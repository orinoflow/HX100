module dxj_top (
input  D11636_SN   ,
input  D505_B      ,
input  D540_GN     ,
input  D2636_B     ,
input  D2667_B     ,
input  D2668_B     ,
input  D2670_B     ,
input  D2671_B     ,
input  D8695_A     ,
input  D8696_A     ,
input  D9934_A     ,
input  D9942_A     ,
input  D9947_A     ,
input  D11631_A    ,
input  D11632_A    ,
input  D12177_RN   ,
input  D13846_A    ,
input  D13859_A    ,
input  D15251_B    ,
input  D15252_B    ,
input  D16018_B    ,
input  D16019_B    ,
input  D16020_B    ,
input  D16021_B    ,
input  D16022_B    ,
input  D16023_B    ,
input  D16024_B    ,
input  D16025_B    ,
input  D16026_B    ,
input  D16027_B    ,
input  D16028_B    ,
input  D16029_B    ,
input  D16030_B    ,
input  D16031_B    ,
input  D16032_B    ,
input  D16033_B    ,
input  D16034_B    ,
input  D16035_B    ,
input  D16036_B    ,
input  D16037_B    ,
input  D16038_B    ,
input  D16039_B    ,
input  D16046_B    ,
input  D16073_B    ,
input  D16074_B    ,
input  D16075_B    ,
input  D16076_B    ,
input  D16081_B    ,
input  D16083_B    ,
input  D16084_B    ,
input  D16099_B    ,
input  D16138_AN   ,
output D499_Y      ,
output D547_Y      ,
output D2144_Y     ,
output D2356_Y     ,
output D9348_Y     ,
output D9936_Y     ,
output D9937_Y     ,
output D9938_Y     ,
output D9939_Y     ,
output D9944_Y     ,
output D9945_Y     ,
output D9952_Y     ,
output D9953_Y     ,
output D9954_Y     ,
output D10115_Y    ,
output D10140_Y    ,
output D10148_Y    ,
output D10149_Y    ,
output D10156_Y    ,
output D10163_Y    ,
output D10373_Y    ,
output D10660_Y    ,
output D12654_Y    ,
output D12655_Y    ,
output D12670_Y    ,
output D13153_Y    ,
output D13155_Y    ,
output D13172_Y    ,
output D14584_Y    ,
output D14585_Y    ,
output D14594_Y    ,
output D14599_Y    ,
output D14610_Y    ,
output D7464_Y     ,
output D15245_Y    ,
output D15247_Y    ,
output D15442_Y    ,
output D16311_Y    ,
output D16403_Y    ,
output D9951_Y     ,
output D9323_Q     ,
output D9353_Q     ,
output D9322_Q     ,
output D9318_Q     ,
output D9336_Q     ,
output D9324_Q     ,
output D9267_Y     ,
output D453_Y      ,
output D10164_Y    ,
output D13204_Y    ,
output D2470_Y     ,
output D16288_Q    ,
output D16404_Y    ,
output D15710_Y    ,
output D2686_Y     ,
output D16300_Y    ,
output D16371_Y    ,
output D15956_Y    ,
output D15957_Y    ,
output D959_Y      ,
output D16302_Y    ,
output D16367_Y    ,
output D2687_Y     ,
output D16401_Y    ,
output D16301_Y    ,
output D16338_Y    ,
output D14774_Y    ,
output D14810_Y    ,
output D14759_Y    ,
output D14773_Y    ,
output D14771_Y    ,
output D14772_Y    ,
output D14811_Y    ,
output D3707_Y     
  );

KC_INV_X8 D16310 ( .Y(D16310_Y), .A(D16341_Y));
KC_AOI22_X3 D15696 ( .A1(D16080_Y), .B0(D15616_Y), .B1(D2521_Y),     .Y(D15696_Y), .A0(D14840_Y));
KC_AOI22_X3 D15695 ( .A1(D14829_Y), .B0(D15634_Y), .B1(D2611_Y),     .Y(D15695_Y), .A0(D15709_Y));
KC_AOI22_X3 D15693 ( .A1(D15616_Y), .B0(D9087_Y), .B1(D14840_Y),     .Y(D15693_Y), .A0(D14311_Y));
KC_AOI22_X3 D15692 ( .A1(D15634_Y), .B0(D15653_Y), .B1(D14829_Y),     .Y(D15692_Y), .A0(D15662_Y));
KC_AOI22_X3 D15690 ( .A1(D15634_Y), .B0(D15654_Y), .B1(D14829_Y),     .Y(D15690_Y), .A0(D15653_Y));
KC_AOI22_X3 D15689 ( .A1(D14840_Y), .B0(D15082_Y), .B1(D15616_Y),     .Y(D15689_Y), .A0(D9085_Y));
KC_AOI22_X3 D15687 ( .A1(D14840_Y), .B0(D15149_Y), .B1(D15616_Y),     .Y(D15687_Y), .A0(D8888_Y));
KC_AOI22_X3 D15686 ( .A1(D15616_Y), .B0(D651_Y), .B1(D14840_Y),     .Y(D15686_Y), .A0(D2583_Y));
KC_AOI22_X3 D15685 ( .A1(D14829_Y), .B0(D15659_Y), .B1(D15634_Y),     .Y(D15685_Y), .A0(D15610_Y));
KC_AOI22_X3 D15682 ( .A1(D15634_Y), .B0(D2648_Y), .B1(D14829_Y),     .Y(D15682_Y), .A0(D15654_Y));
KC_AOI22_X3 D15591 ( .A1(D15529_Y), .B0(D15877_Y), .B1(D15506_Y),     .Y(D15591_Y), .A0(D8902_Y));
KC_AOI22_X3 D15590 ( .A1(D15506_Y), .B0(D6524_Y), .B1(D15529_Y),     .Y(D15590_Y), .A0(D15806_Y));
KC_AOI22_X3 D15589 ( .A1(D755_Y), .B0(D15459_Y), .B1(D14750_Y),     .Y(D15589_Y), .A0(D15411_Y));
KC_AOI22_X3 D15588 ( .A1(D755_Y), .B0(D15411_Y), .B1(D14750_Y),     .Y(D15588_Y), .A0(D15552_Y));
KC_AOI22_X3 D15585 ( .A1(D14750_Y), .B0(D755_Y), .B1(D15341_Y),     .Y(D15585_Y), .A0(D15553_Y));
KC_AOI22_X3 D15584 ( .A1(D16200_Y), .B0(D15506_Y), .B1(D14181_Y),     .Y(D15584_Y), .A0(D15529_Y));
KC_NAND2_X6 D15694 ( .Y(D15694_Y), .B(D15696_Y), .A(D15695_Y));
KC_NAND2_X6 D15691 ( .Y(D15691_Y), .B(D15693_Y), .A(D15692_Y));
KC_NAND2_X6 D15688 ( .Y(D15688_Y), .B(D15689_Y), .A(D15690_Y));
KC_NAND2_X6 D15684 ( .Y(D15684_Y), .B(D15687_Y), .A(D15685_Y));
KC_NAND2_X6 D15683 ( .Y(D15683_Y), .B(D15686_Y), .A(D15682_Y));
KC_NAND2_X6 D15587 ( .Y(D15587_Y), .B(D15590_Y), .A(D15589_Y));
KC_NAND2_X6 D15586 ( .Y(D15586_Y), .B(D15591_Y), .A(D15588_Y));
KC_NAND2_X6 D15583 ( .Y(D15583_Y), .B(D15584_Y), .A(D15585_Y));
KC_MXI2_X8 D16078 ( .Y(D16078_Y), .A(D15239_Y), .BN(D15228_Y),     .S0(D16007_Y));
KC_MXI2_X8 D16077 ( .Y(D16077_Y), .A(D15258_Y), .BN(D14586_Y),     .S0(D15242_Y));
KC_BUF_X15 D14527 ( .Y(D14527_Y), .A(D2574_Q));
KC_OAI211_X3 D14115 ( .B(D14133_Y), .C0(D13309_Y), .A(D14029_Y),     .C1(D13313_Y), .Y(D14115_Y));
KC_XOR2_X5 D16203 ( .Y(D16203_Y), .A(D13320_Y), .B(D13376_Y));
KC_OAI21_X4 D10131 ( .A1(D10099_Y), .B(D10130_Y), .A0(D10085_Y),     .Y(D10131_Y));
KC_NOR2B_X4 D10126 ( .B(D10057_Y), .Y(D10126_Y), .AN(D10048_Q));
KC_AND2BB_X1 D10116 ( .BN(D10106_Y), .Y(D10116_Y), .AN(D10069_Y));
KC_AND2BB_X1 D10115 ( .BN(D10101_Y), .Y(D10115_Y), .AN(D10086_Y));
KC_AND2B_X1 D1665 ( .Y(D1665_Y), .A(D9599_Y), .B(D2110_Y));
KC_OR2_X3 D11634 ( .Y(D11634_Y), .B(D704_Q), .A(D7404_Y));
KC_OR2_X3 D9362 ( .Y(D9362_Y), .B(D9357_Y), .A(D9349_Y));
KC_INV_X4 D9321 ( .Y(D9321_Y), .A(D9947_Y));
KC_MXI2_X9 D16096 ( .Y(D16096_Y), .A(D8294_Y), .BN(D8356_Y),     .S0(D9616_Y));
KC_OAI211B_X2 D6490 ( .B(D8002_Y), .C1(D9371_Y), .A(D1845_Y),     .C0N(D2042_Y), .Y(D6490_Y));
KC_MXI2_X6 D10103 ( .Y(D10103_Y), .B(D10094_Y), .AN(D9456_Y),     .S0(D10091_Y));
KC_MXI2_X6 D16755 ( .Y(D16755_Y), .B(D7669_Y), .AN(D7967_Q),     .S0(D8073_Q));
KC_AO22_X2 D8063 ( .Y(D8063_Y), .B1(D8398_Y), .B0(D8019_Y),     .A1(D3829_Y), .A0(D620_Y));
KC_AO22_X2 D8062 ( .Y(D8062_Y), .B1(D8417_Y), .B0(D8019_Y),     .A1(D5366_Y), .A0(D620_Y));
KC_NAND3_X3 D9298 ( .Y(D9298_Y), .C(D9292_Y), .B(D9290_Y),     .A(D9101_Y));
KC_NAND3_X3 D7991 ( .Y(D7991_Y), .C(D7992_Y), .B(D7940_Y),     .A(D7930_Y));
KC_OAI211_X2 D7990 ( .B(D7939_Y), .C0(D7922_Y), .A(D7989_Y),     .C1(D7946_Y), .Y(D7990_Y));
KC_AOI32_X2 D15608 ( .B1(D15511_Y), .A2(D15494_Y), .Y(D15608_Y),     .A1(D15511_Y), .B0(D15607_Y), .A0(D15387_Y));
KC_AOI32_X2 D13640 ( .B1(D13590_Y), .A2(D13545_Y), .Y(D13640_Y),     .A1(D13590_Y), .B0(D13409_Y), .A0(D13588_Y));
KC_AOI32_X2 D7820 ( .B1(D12301_Y), .A2(D7758_Y), .Y(D7820_Y),     .A1(D12301_Y), .B0(D7779_Y), .A0(D9237_Y));
KC_TINV_X4 D7522 ( .Y(D7522_Y), .A(D7557_Y), .OE(D6110_Y));
KC_BUF_X5 D16659 ( .Y(D16659_Y), .A(D11630_Y));
KC_BUF_X5 D15867 ( .Y(D15867_Y), .A(D15004_Y));
KC_BUF_X5 D12743 ( .Y(D12743_Y), .A(D11638_Q));
KC_BUF_X5 D11627 ( .Y(D11627_Y), .A(D11641_Q));
KC_BUF_X5 D11172 ( .Y(D11172_Y), .A(D11163_Y));
KC_BUF_X5 D7520 ( .Y(D7520_Y), .A(D9315_Y));
KC_TINV_X6 D15450 ( .Y(D15450_Y), .OE(D9136_Y), .A(D7630_Y));
KC_TINV_X6 D15448 ( .Y(D15448_Y), .OE(D1939_Y), .A(D22_Y));
KC_NAND4_X4 D7488 ( .Y(D7488_Y), .D(D7455_Y), .C(D7439_Y), .B(D6019_Y),     .A(D6022_Y));
KC_OR4_X1 D7404 ( .Y(D7404_Y), .C(D5692_Q), .B(D7470_Y), .D(D7274_Y),     .A(D7148_Q));
KC_OR4_X1 D7402 ( .Y(D7402_Y), .C(D7391_Q), .B(D7148_Q), .D(D8903_Y),     .A(D7412_Q));
KC_AND4_X2 D7401 ( .D(D7274_Y), .C(D7328_Y), .B(D7327_Y), .A(D6022_Y),     .Y(D7401_Y));
KC_NOR3B_X1 D16667 ( .Y(D16667_Y), .B(D16672_Y), .CN(D1373_Q),     .A(D16684_Q));
KC_NOR3B_X1 D16641 ( .Y(D16641_Y), .B(D16623_Y), .CN(D16609_Y),     .A(D1400_Q));
KC_NOR3B_X1 D16464 ( .Y(D16464_Y), .B(D16437_Y), .CN(D16440_Y),     .A(D1281_Y));
KC_NOR3B_X1 D14708 ( .Y(D14708_Y), .B(D14639_Y), .CN(D13947_Y),     .A(D13940_Y));
KC_NOR3B_X1 D14005 ( .Y(D14005_Y), .B(D13953_Y), .CN(D13936_Y),     .A(D16559_Y));
KC_NOR3B_X1 D14003 ( .Y(D14003_Y), .B(D13971_Y), .CN(D16117_Y),     .A(D16226_Q));
KC_NOR3B_X1 D12296 ( .Y(D12296_Y), .B(D12261_Y), .CN(D12207_Y),     .A(D2358_Y));
KC_NOR3B_X1 D9492 ( .Y(D9492_Y), .B(D7402_Y), .CN(D9471_Q),     .A(D9582_Q));
KC_NOR3B_X1 D6496 ( .Y(D6496_Y), .B(D468_Y), .CN(D471_Y), .A(D6437_Y));
KC_NOR3B_X1 D6495 ( .Y(D6495_Y), .B(D7929_Y), .CN(D6420_Y),     .A(D7920_Y));
KC_OAI21BB_X2 D14270 ( .BN(D13391_Y), .A1N(D14264_Q), .A0(D14207_Y),     .Y(D14270_Y));
KC_OAI21BB_X2 D13 ( .BN(D294_Y), .A1N(D7426_Y), .A0(D7486_Y),     .Y(D13_Y));
KC_OAI21BB_X2 D6487 ( .BN(D6381_Q), .A1N(D1793_Q), .A0(D6483_Y),     .Y(D6487_Y));
KC_MXI2_X7 D16079 ( .Y(D16079_Y), .A(D16175_Y), .BN(D16104_Y),     .S0(D16106_Y));
KC_MXI2_X7 D15451 ( .Y(D15451_Y), .A(D7701_Y), .BN(D7649_Y),     .S0(D7640_Y));
KC_MXI2_X7 D9144 ( .Y(D9144_Y), .A(D6173_Y), .BN(D13173_Y),     .S0(D6268_Y));
KC_MXI2_X4 D16754 ( .Y(D16754_Y), .A(D7761_Y), .B(D6305_Y),     .S0(D7761_Y));
KC_MXI2_X4 D7617 ( .Y(D7617_Y), .A(D7558_Y), .B(D7573_Y),     .S0(D7558_Y));
KC_MXI2_X4 D6360 ( .Y(D6360_Y), .A(D6336_Y), .B(D6296_Y),     .S0(D6336_Y));
KC_MXI2_X4 D6209 ( .Y(D6209_Y), .A(D6139_Y), .B(D365_Q), .S0(D6139_Y));
KC_AND2B_X2 D1957 ( .Y(D1957_Y), .A(D6087_Y), .B(D6100_Y));
KC_NOR3B_X2 D10097 ( .Y(D10097_Y), .B(D10081_Y), .CN(D9942_Y),     .A(D10080_Y));
KC_NOR3B_X2 D18 ( .Y(D18_Y), .B(D5997_Y), .CN(D5954_Y), .A(D6096_Y));
KC_NOR2_X2 D7164 ( .Y(D7164_Y), .B(D7252_Y), .A(D5756_Y));
KC_NOR2_X2 D5966 ( .Y(D5966_Y), .B(D6075_Y), .A(D7469_Y));
KC_XOR2_X1 D5707 ( .Y(D5707_Y), .A(D5699_Y), .B(D6275_Y));
KC_OAI22B_X1 D15337 ( .A1(D16068_Y), .B0(D16067_Y), .A0(D15281_Y),     .B1N(D15288_Y), .Y(D15337_Y));
KC_OAI22B_X1 D14909 ( .A1(D14809_Y), .B0(D14091_Q), .A0(D14877_Q),     .B1N(D14169_Q), .Y(D14909_Y));
KC_OAI22B_X1 D13413 ( .A1(D13401_Y), .B0(D13300_Y), .A0(D13321_Y),     .B1N(D855_Q), .Y(D13413_Y));
KC_OAI22B_X1 D13412 ( .A1(D13319_Y), .B0(D13299_Y), .A0(D13322_Y),     .B1N(D852_Q), .Y(D13412_Y));
KC_OAI22B_X1 D13407 ( .A1(D13401_Y), .B0(D13406_Y), .A0(D13309_Y),     .B1N(D814_Q), .Y(D13407_Y));
KC_OAI22B_X1 D12370 ( .A1(D12869_Y), .B0(D12313_Y), .A0(D12315_Y),     .B1N(D12346_Q), .Y(D12370_Y));
KC_OAI22B_X1 D9987 ( .A1(D216_Y), .B0(D9955_Y), .A0(D9971_Y),     .B1N(D9981_Q), .Y(D9987_Y));
KC_OAI22B_X1 D9986 ( .A1(D216_Y), .B0(D9966_Y), .A0(D9972_Y),     .B1N(D8823_Q), .Y(D9986_Y));
KC_OAI22B_X1 D9590 ( .A1(D9574_Q), .B0(D9547_Y), .A0(D9577_Q),     .B1N(D9534_Y), .Y(D9590_Y));
KC_OAI22B_X1 D6492 ( .A1(D4863_Y), .B0(D469_Y), .A0(D1700_Y),     .B1N(D480_Q), .Y(D6492_Y));
KC_OAI22B_X1 D4980 ( .A1(D4866_Y), .B0(D4896_Y), .A0(D4868_Y),     .B1N(D4887_Y), .Y(D4980_Y));
KC_OAI22B_X1 D4978 ( .A1(D4895_Y), .B0(D4894_Y), .A0(D1567_Y),     .B1N(D445_Q), .Y(D4978_Y));
KC_OAI22B_X1 D4975 ( .A1(D1566_Y), .B0(D4909_Y), .A0(D3498_Y),     .B1N(D3378_Y), .Y(D4975_Y));
KC_AND2_X6 D10204 ( .Y(D10204_Y), .A(D6328_Y), .B(D7703_Y));
KC_AND2_X6 D10026 ( .Y(D10026_Y), .A(D4702_Y), .B(D4664_Y));
KC_AND4B_X1 D16586 ( .B(D16382_Y), .C(D16654_Y), .D(D16612_Y),     .Y(D16586_Y), .AN(D16608_Y));
KC_AND4B_X1 D8476 ( .B(D8369_Y), .C(D8368_Y), .D(D8403_Y), .Y(D8476_Y),     .AN(D8382_Y));
KC_AND4B_X1 D4650 ( .B(D4687_Y), .C(D4659_Y), .D(D1427_Y), .Y(D4650_Y),     .AN(D3098_Y));
KC_AND3_X1 D14114 ( .C(D14008_Y), .B(D13318_Y), .A(D14133_Y),     .Y(D14114_Y));
KC_AND3_X1 D8264 ( .C(D8243_Q), .B(D8245_Q), .A(D8244_Q), .Y(D8264_Y));
KC_AND3_X1 D6494 ( .C(D7916_Y), .B(D6480_Q), .A(D524_Q), .Y(D6494_Y));
KC_AND3_X1 D4402 ( .C(D5890_Y), .B(D4320_Y), .A(D4457_Y), .Y(D4402_Y));
KC_TINV_X3 D16771 ( .Y(D16771_Y), .A(D16475_Q), .OE(D13326_Y));
KC_TINV_X3 D14610 ( .Y(D14610_Y), .A(D2571_Y), .OE(D14601_Q));
KC_TINV_X3 D16767 ( .Y(D16767_Y), .A(D14282_Y), .OE(D14276_Y));
KC_TINV_X3 D6273 ( .Y(D6273_Y), .A(D5380_Y), .OE(D5417_Y));
KC_TINV_X3 D3499 ( .Y(D3499_Y), .A(D3482_Q), .OE(D16006_Y));
KC_TINV_X3 D3498 ( .Y(D3498_Y), .A(D3588_Y), .OE(D3483_Q));
KC_TINV_X3 D3400 ( .Y(D3400_Y), .A(D3366_Y), .OE(D1517_Q));
KC_AND4_X1 D16281 ( .D(D16261_Y), .C(D16256_Y), .B(D16265_Y),     .A(D16290_Q), .Y(D16281_Y));
KC_AND4_X1 D16279 ( .D(D15630_Y), .C(D16256_Y), .B(D16273_Y),     .A(D16289_Q), .Y(D16279_Y));
KC_AND4_X1 D15943 ( .D(D15884_Y), .C(D15888_Y), .B(D15882_Y),     .A(D15897_Y), .Y(D15943_Y));
KC_AND4_X1 D15865 ( .D(D15820_Y), .C(D15829_Y), .B(D15818_Y),     .A(D15823_Y), .Y(D15865_Y));
KC_AND4_X1 D14994 ( .D(D16359_Q), .C(D16361_Q), .B(D14304_Q),     .A(D2516_Q), .Y(D14994_Y));
KC_AND4_X1 D14471 ( .D(D14413_Y), .C(D14424_Y), .B(D14414_Y),     .A(D13719_Y), .Y(D14471_Y));
KC_AND4_X1 D14470 ( .D(D15172_Y), .C(D1269_Y), .B(D14418_Y),     .A(D15106_Y), .Y(D14470_Y));
KC_AND4_X1 D13753 ( .D(D1185_Y), .C(D13779_Y), .B(D13774_Y),     .A(D13716_Y), .Y(D13753_Y));
KC_AND4_X1 D13700 ( .D(D13670_Y), .C(D13671_Y), .B(D13646_Y),     .A(D13645_Y), .Y(D13700_Y));
KC_AND4_X1 D12221 ( .D(D12228_Y), .C(D16129_Y), .B(D12231_Y),     .A(D12229_Y), .Y(D12221_Y));
KC_AND4_X1 D9320 ( .D(D10142_Y), .C(D9269_Y), .B(D9268_Y), .A(D9266_Y),     .Y(D9320_Y));
KC_AND4_X1 D9002 ( .D(D8963_Y), .C(D342_Y), .B(D7492_Y), .A(D8959_Y),     .Y(D9002_Y));
KC_AND4_X1 D8804 ( .D(D8756_Y), .C(D9481_Y), .B(D9476_Y), .A(D9480_Y),     .Y(D8804_Y));
KC_AND4_X1 D4465 ( .D(D4416_Y), .C(D5953_Y), .B(D165_Y), .A(D5969_Y),     .Y(D4465_Y));
KC_AND4_X1 D4226 ( .D(D4097_Y), .C(D4092_Y), .B(D5754_Y), .A(D4204_Y),     .Y(D4226_Y));
KC_AND4_X1 D3863 ( .D(D3848_Y), .C(D1478_Y), .B(D3849_Y), .A(D1504_Y),     .Y(D3863_Y));
KC_AND4_X1 D3362 ( .D(D3275_Y), .C(D3329_Y), .B(D3369_Y), .A(D3384_Q),     .Y(D3362_Y));
KC_AND4_X1 D3061 ( .D(D44_Y), .C(D3084_Q), .B(D1516_Q), .A(D3078_Q),     .Y(D3061_Y));
KC_TINV_X5 D582 ( .A(D2938_Y), .Y(D582_Y), .OE(D2982_Y));
KC_OAI21B_X2 D14269 ( .A1(D1092_Y), .A0(D870_Y), .BN(D14084_Y),     .Y(D14269_Y));
KC_OAI21B_X2 D12295 ( .A1(D648_Y), .A0(D12249_Y), .BN(D12246_Y),     .Y(D12295_Y));
KC_OAI21B_X2 D10367 ( .A1(D10318_Y), .A0(D10361_Q), .BN(D10362_Q),     .Y(D10367_Y));
KC_OAI21B_X2 D9296 ( .A1(D7784_Y), .A0(D417_Y), .BN(D9111_Y),     .Y(D9296_Y));
KC_OAI21B_X2 D9295 ( .A1(D7785_Y), .A0(D417_Y), .BN(D9106_Y),     .Y(D9295_Y));
KC_OAI21B_X2 D9294 ( .A1(D10162_Y), .A0(D417_Y), .BN(D9111_Y),     .Y(D9294_Y));
KC_OAI21B_X2 D9293 ( .A1(D7730_Y), .A0(D417_Y), .BN(D9106_Y),     .Y(D9293_Y));
KC_OAI21B_X2 D8257 ( .A1(D8296_Y), .A0(D1943_Q), .BN(D1956_Y),     .Y(D8257_Y));
KC_OAI21B_X2 D7403 ( .A1(D4285_Y), .A0(D7361_Y), .BN(D149_Q),     .Y(D7403_Y));
KC_OAI21B_X2 D7400 ( .A1(D7398_Y), .A0(D4434_Y), .BN(D7389_Y),     .Y(D7400_Y));
KC_OAI21B_X2 D7302 ( .A1(D222_Y), .A0(D204_Y), .BN(D7173_Y),     .Y(D7302_Y));
KC_OAI21B_X2 D2808 ( .A1(D2775_Y), .A0(D2845_Y), .BN(D2761_Y),     .Y(D2808_Y));
KC_INV_X3 D16752 ( .Y(D16752_Y), .A(D3054_Y));
KC_INV_X3 D16751 ( .Y(D16751_Y), .A(D4531_Y));
KC_INV_X3 D16750 ( .Y(D16750_Y), .A(D4534_Y));
KC_INV_X3 D16749 ( .Y(D16749_Y), .A(D4533_Y));
KC_INV_X3 D16748 ( .Y(D16748_Y), .A(D315_Y));
KC_INV_X3 D16747 ( .Y(D16747_Y), .A(D10005_Y));
KC_INV_X3 D16746 ( .Y(D16746_Y), .A(D4532_Y));
KC_INV_X3 D16742 ( .Y(D16742_Y), .A(D3056_Y));
KC_INV_X3 D16741 ( .Y(D16741_Y), .A(D4538_Y));
KC_INV_X3 D16740 ( .Y(D16740_Y), .A(D3057_Y));
KC_INV_X3 D16739 ( .Y(D16739_Y), .A(D4544_Y));
KC_INV_X3 D16738 ( .Y(D16738_Y), .A(D3055_Y));
KC_INV_X3 D16737 ( .Y(D16737_Y), .A(D4537_Y));
KC_INV_X3 D10157 ( .Y(D10157_Y), .A(D12300_Y));
KC_INV_X3 D7713 ( .Y(D7713_Y), .A(D12762_Y));
KC_INV_X3 D3597 ( .Y(D3597_Y), .A(D16742_Y));
KC_INV_X3 D3596 ( .Y(D3596_Y), .A(D16752_Y));
KC_INV_X3 D3595 ( .Y(D3595_Y), .A(D16749_Y));
KC_INV_X3 D3593 ( .Y(D3593_Y), .A(D16739_Y));
KC_INV_X3 D3592 ( .Y(D3592_Y), .A(D2698_Y));
KC_INV_X3 D3591 ( .Y(D3591_Y), .A(D16747_Y));
KC_INV_X3 D3590 ( .Y(D3590_Y), .A(D16740_Y));
KC_INV_X3 D3589 ( .Y(D3589_Y), .A(D2699_Y));
KC_INV_X3 D3570 ( .Y(D3570_Y), .A(D16741_Y));
KC_INV_X3 D3569 ( .Y(D3569_Y), .A(D16737_Y));
KC_INV_X3 D3568 ( .Y(D3568_Y), .A(D2697_Y));
KC_INV_X3 D3567 ( .Y(D3567_Y), .A(D16746_Y));
KC_INV_X3 D3566 ( .Y(D3566_Y), .A(D16748_Y));
KC_INV_X3 D3565 ( .Y(D3565_Y), .A(D16750_Y));
KC_INV_X3 D3563 ( .Y(D3563_Y), .A(D16738_Y));
KC_INV_X3 D3562 ( .Y(D3562_Y), .A(D16751_Y));
KC_INV_X3 D2726 ( .Y(D2726_Y), .A(D3569_Y));
KC_INV_X3 D2725 ( .Y(D2725_Y), .A(D3570_Y));
KC_INV_X3 D2735 ( .Y(D2735_Y), .A(D3563_Y));
KC_INV_X3 D2734 ( .Y(D2734_Y), .A(D3596_Y));
KC_INV_X3 D2733 ( .Y(D2733_Y), .A(D3590_Y));
KC_INV_X3 D2732 ( .Y(D2732_Y), .A(D3589_Y));
KC_INV_X3 D2731 ( .Y(D2731_Y), .A(D3592_Y));
KC_INV_X3 D2730 ( .Y(D2730_Y), .A(D3595_Y));
KC_INV_X3 D2729 ( .Y(D2729_Y), .A(D3597_Y));
KC_INV_X3 D2724 ( .Y(D2724_Y), .A(D3567_Y));
KC_INV_X3 D2723 ( .Y(D2723_Y), .A(D3565_Y));
KC_INV_X3 D2722 ( .Y(D2722_Y), .A(D3593_Y));
KC_INV_X3 D2721 ( .Y(D2721_Y), .A(D3591_Y));
KC_INV_X3 D2720 ( .Y(D2720_Y), .A(D3568_Y));
KC_INV_X3 D2719 ( .Y(D2719_Y), .A(D3562_Y));
KC_INV_X3 D2718 ( .Y(D2718_Y), .A(D3566_Y));
KC_INV_X3 D2699 ( .Y(D2699_Y), .A(D4539_Y));
KC_INV_X3 D2698 ( .Y(D2698_Y), .A(D4545_Y));
KC_INV_X3 D2697 ( .Y(D2697_Y), .A(D4530_Y));
KC_MX2_X1 D12174 ( .Y(D12174_Y), .A(D12175_Y), .B(D540_Q),     .S0(D12183_Y));
KC_MX2_X1 D8324 ( .Y(D8324_Y), .A(D8354_Y), .B(D8353_Y), .S0(D8312_Y));
KC_MX2_X1 D7579 ( .Y(D7579_Y), .A(D314_Y), .B(D1706_Y), .S0(D6239_Y));
KC_MX2_X1 D7526 ( .Y(D7526_Y), .A(D281_Y), .B(D1706_Y), .S0(D6239_Y));
KC_MX2_X1 D3764 ( .Y(D3764_Y), .A(D3750_Y), .B(D5253_Y), .S0(D4406_Y));
KC_MX2_X1 D3366 ( .Y(D3366_Y), .A(D6369_Y), .B(D3310_Y), .S0(D3392_Y));
KC_MX2_X1 D3272 ( .Y(D3272_Y), .A(D3222_Y), .B(D3276_Y), .S0(D3249_Y));
KC_MX2_X1 D2262 ( .Y(D2262_Y), .A(D11346_Y), .B(D11418_Y),     .S0(D11417_Y));
KC_AND2_X5 D13841 ( .B(D13844_Y), .A(D14315_Y), .Y(D13841_Y));
KC_AND2_X5 D13840 ( .B(D13844_Y), .A(D14315_Y), .Y(D13840_Y));
KC_AND2_X5 D2176 ( .B(D10298_Q), .A(D2158_Y), .Y(D2176_Y));
KC_MXI2_X5 D7464 ( .Y(D7464_Y), .A(D14549_Y), .B(D14553_Y),     .S0(D14567_Y));
KC_MXI2_X5 D16765 ( .Y(D16765_Y), .A(D13197_Q), .B(D13208_Q),     .S0(D14711_Y));
KC_MXI2_X5 D16762 ( .Y(D16762_Y), .A(D10159_Y), .B(D13288_Y),     .S0(D13157_Y));
KC_MXI2_X5 D7824 ( .Y(D7824_Y), .A(D7481_Q), .B(D409_Y), .S0(D6342_Y));
KC_MXI2_X5 D7757 ( .Y(D7757_Y), .A(D9021_Q), .B(D410_Y), .S0(D6239_Y));
KC_MXI2_X5 D7756 ( .Y(D7756_Y), .A(D8953_Q), .B(D4786_Y),     .S0(D6239_Y));
KC_MXI2_X5 D7755 ( .Y(D7755_Y), .A(D723_Q), .B(D7730_Y), .S0(D6351_Q));
KC_MXI2_X5 D6288 ( .Y(D6288_Y), .A(D239_Q), .B(D4713_Y), .S0(D6239_Y));
KC_MXI2_X5 D6287 ( .Y(D6287_Y), .A(D4235_Q), .B(D4549_Y),     .S0(D6239_Y));
KC_MXI2_X5 D6285 ( .Y(D6285_Y), .A(D8313_Q), .B(D4715_Y),     .S0(D6239_Y));
KC_MXI2_X5 D4747 ( .Y(D4747_Y), .A(D4149_Q), .B(D371_Y), .S0(D6239_Y));
KC_MXI2_X5 D1976 ( .Y(D1976_Y), .A(D8951_Q), .B(D4842_Y),     .S0(D6342_Y));
KC_NAND2_X5 D16632 ( .Y(D16632_Y), .B(D16639_Y), .A(D16614_Y));
KC_NAND2_X5 D13622 ( .Y(D13622_Y), .B(D13419_Y), .A(D2430_Y));
KC_NAND2_X5 D13619 ( .Y(D13619_Y), .B(D13419_Y), .A(D2429_Y));
KC_NAND2_X5 D8551 ( .Y(D8551_Y), .B(D8534_Y), .A(D8466_Y));
KC_NAND2_X5 D8470 ( .Y(D8470_Y), .B(D8415_Y), .A(D8401_Y));
KC_NAND2_X5 D8060 ( .Y(D8060_Y), .B(D7974_Y), .A(D8210_Y));
KC_NAND2_X5 D5082 ( .Y(D5082_Y), .B(D1563_Y), .A(D3413_Y));
KC_NAND2_X5 D2471 ( .Y(D2471_Y), .B(D13419_Y), .A(D2433_Y));
KC_NAND2_X5 D2099 ( .Y(D2099_Y), .B(D382_Y), .A(D7469_Y));
KC_NAND2_X5 D1954 ( .Y(D1954_Y), .B(D7579_Y), .A(D7526_Y));
KC_AOI222_X1 D9228 ( .A1(D9267_Y), .B0(D9114_Y), .B1(D9219_Q),     .C0(D9102_Y), .C1(D8730_Q), .Y(D9228_Y), .A0(D7631_Y));
KC_AOI222_X1 D7306 ( .A1(D199_Y), .B0(D7193_Y), .B1(D9479_Y),     .C0(D5783_Y), .C1(D273_Y), .Y(D7306_Y), .A0(D7293_Y));
KC_AOI222_X1 D16777 ( .A1(D6929_Y), .B0(D1743_Y), .B1(D8542_Y),     .C0(D6930_Y), .C1(D5587_Y), .Y(D16777_Y), .A0(D1743_Y));
KC_AOI222_X1 D16776 ( .A1(D6924_Y), .B0(D6938_Y), .B1(D8542_Y),     .C0(D6919_Y), .C1(D7021_Y), .Y(D16776_Y), .A0(D6938_Y));
KC_AOI222_X1 D16775 ( .A1(D6927_Y), .B0(D1743_Y), .B1(D8542_Y),     .C0(D6930_Y), .C1(D7074_Y), .Y(D16775_Y), .A0(D1743_Y));
KC_AOI222_X1 D5944 ( .A1(D7242_Y), .B0(D4326_Y), .B1(D5871_Y),     .C0(D5848_Y), .C1(D5872_Y), .Y(D5944_Y), .A0(D4341_Y));
KC_AOI222_X1 D4263 ( .A1(D228_Q), .B0(D4167_Y), .B1(D4242_Y),     .C0(D7291_Y), .C1(D4158_Y), .Y(D4263_Y), .A0(D5753_Y));
KC_AOI222_X1 D4262 ( .A1(D8313_Q), .B0(D7288_Y), .B1(D4158_Y),     .C0(D4250_Y), .C1(D3572_Y), .Y(D4262_Y), .A0(D5753_Y));
KC_AOI222_X1 D4257 ( .A1(D165_Y), .B0(D5713_Y), .B1(D5768_Y),     .C0(D4167_Y), .C1(D4243_Y), .Y(D4257_Y), .A0(D5753_Y));
KC_AOI222_X1 D3494 ( .A1(D3477_Y), .B0(D3463_Y), .B1(D3388_Q),     .C0(D3428_Y), .C1(D3409_Y), .Y(D3494_Y), .A0(D3461_Y));
KC_AOI222_X1 D3493 ( .A1(D1570_Y), .B0(D3372_Q), .B1(D4897_Y),     .C0(D69_Y), .C1(D4900_Y), .Y(D3493_Y), .A0(D4923_Y));
KC_AOI222_X1 D16774 ( .A1(D8095_Y), .B0(D8130_Y), .B1(D1840_Y),     .C0(D8095_Y), .C1(D741_Y), .Y(D16774_Y), .A0(D8130_Y));
KC_AOI222_X1 D1969 ( .A1(D5698_Y), .B0(D7194_Y), .B1(D1886_Y),     .C0(D7295_Y), .C1(D7184_Y), .Y(D1969_Y), .A0(D5929_Y));
KC_AOI222_X1 D16773 ( .A1(D1585_Y), .B0(D4449_Y), .B1(D4447_Y),     .C0(D4279_Y), .C1(D4396_Y), .Y(D16773_Y), .A0(D4449_Y));
KC_TINV_X2 D1677 ( .Y(D1677_Y), .A(D2909_Y), .OE(D7636_Y));
KC_NAND3B_X1 D16582 ( .Y(D16582_Y), .A(D16382_Y), .CN(D16285_Y),     .B(D16299_Y));
KC_NAND3B_X1 D16460 ( .Y(D16460_Y), .A(D16470_Q), .CN(D16432_Y),     .B(D16439_Y));
KC_NAND3B_X1 D16398 ( .Y(D16398_Y), .A(D16436_Y), .CN(D16431_Y),     .B(D16470_Q));
KC_NAND3B_X1 D16169 ( .Y(D16169_Y), .A(D16118_Y), .CN(D16174_Y),     .B(D2655_Y));
KC_NAND3B_X1 D16168 ( .Y(D16168_Y), .A(D16105_Y), .CN(D16112_Y),     .B(D16095_Y));
KC_NAND3B_X1 D15582 ( .Y(D15582_Y), .A(D15534_Y), .CN(D15530_Y),     .B(D15362_Y));
KC_NAND3B_X1 D14097 ( .Y(D14097_Y), .A(D14665_Y), .CN(D14044_Y),     .B(D13977_Y));
KC_NAND3B_X1 D13403 ( .Y(D13403_Y), .A(D13330_Y), .CN(D13402_Y),     .B(D13340_Y));
KC_NAND3B_X1 D13402 ( .Y(D13402_Y), .A(D13361_Y), .CN(D13325_Y),     .B(D13372_Y));
KC_NAND3B_X1 D13401 ( .Y(D13401_Y), .A(D13256_Y), .CN(D12241_Y),     .B(D7668_Y));
KC_NAND3B_X1 D11112 ( .Y(D11112_Y), .A(D11101_Y), .CN(D10605_Y),     .B(D11101_Y));
KC_NAND3B_X1 D10819 ( .Y(D10819_Y), .A(D10831_Y), .CN(D10870_Y),     .B(D10870_Y));
KC_NAND3B_X1 D9946 ( .Y(D9946_Y), .A(D9925_Y), .CN(D9966_Y),     .B(D9933_Y));
KC_NAND3B_X1 D9281 ( .Y(D9281_Y), .A(D9258_Y), .CN(D8893_Y),     .B(D9200_Y));
KC_NAND3B_X1 D9152 ( .Y(D9152_Y), .A(D6095_Y), .CN(D7700_Y),     .B(D9179_Y));
KC_NAND3B_X1 D8827 ( .Y(D8827_Y), .A(D8750_Y), .CN(D2028_Y),     .B(D8792_Y));
KC_NAND3B_X1 D8718 ( .Y(D8718_Y), .A(D8685_Y), .CN(D8685_Y),     .B(D61_Y));
KC_NAND3B_X1 D8717 ( .Y(D8717_Y), .A(D8671_Y), .CN(D8685_Y),     .B(D8685_Y));
KC_NAND3B_X1 D8351 ( .Y(D8351_Y), .A(D16755_Y), .CN(D8047_Y),     .B(D8292_Y));
KC_NAND3B_X1 D8350 ( .Y(D8350_Y), .A(D8047_Y), .CN(D16755_Y),     .B(D8292_Y));
KC_NAND3B_X1 D8254 ( .Y(D8254_Y), .A(D8250_Q), .CN(D8204_Y),     .B(D1840_Y));
KC_NAND3B_X1 D8157 ( .Y(D8157_Y), .A(D5174_Y), .CN(D8060_Y),     .B(D8102_Y));
KC_NAND3B_X1 D8156 ( .Y(D8156_Y), .A(D8108_Y), .CN(D9437_Y),     .B(D8120_Y));
KC_NAND3B_X1 D7975 ( .Y(D7975_Y), .A(D6787_Y), .CN(D7921_Y),     .B(D7931_Y));
KC_NAND3B_X1 D7797 ( .Y(D7797_Y), .A(D7762_Y), .CN(D7792_Y),     .B(D447_Y));
KC_NAND3B_X1 D7739 ( .Y(D7739_Y), .A(D7709_Y), .CN(D7673_Y),     .B(D7710_Y));
KC_NAND3B_X1 D7396 ( .Y(D7396_Y), .A(D7225_Y), .CN(D8841_Y),     .B(D5840_Y));
KC_NAND3B_X1 D7395 ( .Y(D7395_Y), .A(D7438_Y), .CN(D6071_Y),     .B(D7340_Y));
KC_NAND3B_X1 D7297 ( .Y(D7297_Y), .A(D8734_Y), .CN(D7224_Y),     .B(D7214_Y));
KC_NAND3B_X1 D6489 ( .Y(D6489_Y), .A(D485_Q), .CN(D6433_Y),     .B(D6481_Q));
KC_NAND3B_X1 D6272 ( .Y(D6272_Y), .A(D6282_Y), .CN(D6227_Y),     .B(D6244_Y));
KC_NAND3B_X1 D6269 ( .Y(D6269_Y), .A(D6265_Y), .CN(D13173_Y),     .B(D6235_Y));
KC_NAND3B_X1 D6079 ( .Y(D6079_Y), .A(D6035_Y), .CN(D6014_Y),     .B(D6009_Y));
KC_NAND3B_X1 D6078 ( .Y(D6078_Y), .A(D7353_Y), .CN(D5963_Y),     .B(D5952_Y));
KC_NAND3B_X1 D5935 ( .Y(D5935_Y), .A(D6019_Y), .CN(D5835_Y),     .B(D5864_Y));
KC_NAND3B_X1 D4740 ( .Y(D4740_Y), .A(D1571_Y), .CN(D4734_Y),     .B(D4741_Y));
KC_NAND3B_X1 D4730 ( .Y(D4730_Y), .A(D4735_Y), .CN(D4654_Y),     .B(D10026_Y));
KC_NAND3B_X1 D4124 ( .Y(D4124_Y), .A(D4547_Y), .CN(D1653_Y),     .B(D2716_Y));
KC_NAND3B_X1 D3389 ( .Y(D3389_Y), .A(D3342_Y), .CN(D3357_Y),     .B(D1454_Y));
KC_NAND3B_X1 D3192 ( .Y(D3192_Y), .A(D1430_Y), .CN(D3188_Q),     .B(D3144_Y));
KC_NAND3B_X1 D2892 ( .Y(D2892_Y), .A(D268_Q), .CN(D2902_Q),     .B(D2792_Y));
KC_NAND3B_X1 D2802 ( .Y(D2802_Y), .A(D2784_Y), .CN(D2783_Y),     .B(D2767_Y));
KC_NAND3B_X1 D1805 ( .Y(D1805_Y), .A(D6172_Y), .CN(D6196_Y),     .B(D56_Y));
KC_NAND3B_X1 D1661 ( .Y(D1661_Y), .A(D4389_Y), .CN(D4546_Y),     .B(D4389_Y));
KC_NAND2_X2 D16722 ( .Y(D16722_Y), .B(D16715_Y), .A(D16720_Y));
KC_NAND2_X2 D16701 ( .Y(D16701_Y), .B(D16772_Y), .A(D16704_Y));
KC_NAND2_X2 D16700 ( .Y(D16700_Y), .B(D16772_Y), .A(D16697_Y));
KC_NAND2_X2 D16615 ( .Y(D16615_Y), .B(D16639_Y), .A(D16649_Y));
KC_NAND2_X2 D16578 ( .Y(D16578_Y), .B(D16588_Y), .A(D16594_Y));
KC_NAND2_X2 D16576 ( .Y(D16576_Y), .B(D16588_Y), .A(D16575_Y));
KC_NAND2_X2 D16313 ( .Y(D16313_Y), .B(D16341_Y), .A(GND));
KC_NAND2_X2 D15132 ( .Y(D15132_Y), .B(D15159_Y), .A(D15124_Y));
KC_NAND2_X2 D15131 ( .Y(D15131_Y), .B(D15159_Y), .A(D15123_Y));
KC_NAND2_X2 D14682 ( .Y(D14682_Y), .B(D14712_Y), .A(D14675_Y));
KC_NAND2_X2 D14681 ( .Y(D14681_Y), .B(D14712_Y), .A(D14674_Y));
KC_NAND2_X2 D13988 ( .Y(D13988_Y), .B(D13996_Q), .A(D13275_Q));
KC_NAND2_X2 D13824 ( .Y(D13824_Y), .B(D13843_Y), .A(D13817_Y));
KC_NAND2_X2 D13823 ( .Y(D13823_Y), .B(D13843_Y), .A(D13818_Y));
KC_NAND2_X2 D13610 ( .Y(D13610_Y), .B(D13419_Y), .A(D13549_Y));
KC_NAND2_X2 D13609 ( .Y(D13609_Y), .B(D1076_Y), .A(D13605_Y));
KC_NAND2_X2 D13607 ( .Y(D13607_Y), .B(D1076_Y), .A(D13604_Y));
KC_NAND2_X2 D13089 ( .Y(D13089_Y), .B(D13094_Y), .A(D13079_Y));
KC_NAND2_X2 D13085 ( .Y(D13085_Y), .B(D13094_Y), .A(D104_Y));
KC_NAND2_X2 D12272 ( .Y(D12272_Y), .B(D12304_Y), .A(D12263_Y));
KC_NAND2_X2 D12269 ( .Y(D12269_Y), .B(D12304_Y), .A(D12262_Y));
KC_NAND2_X2 D12123 ( .Y(D12123_Y), .B(D11612_Y), .A(D12112_Y));
KC_NAND2_X2 D11597 ( .Y(D11597_Y), .B(D11612_Y), .A(D11593_Y));
KC_NAND2_X2 D11334 ( .Y(D11334_Y), .B(D11417_Y), .A(D11315_Y));
KC_NAND2_X2 D11333 ( .Y(D11333_Y), .B(D11417_Y), .A(D11316_Y));
KC_NAND2_X2 D11036 ( .Y(D11036_Y), .B(D11055_Y), .A(D11023_Y));
KC_NAND2_X2 D11029 ( .Y(D11029_Y), .B(D11055_Y), .A(D11022_Y));
KC_NAND2_X2 D10799 ( .Y(D10799_Y), .B(D16082_Y), .A(D10786_Y));
KC_NAND2_X2 D10796 ( .Y(D10796_Y), .B(D16082_Y), .A(D10784_Y));
KC_NAND2_X2 D9904 ( .Y(D9904_Y), .B(D8663_Y), .A(D9900_Y));
KC_NAND2_X2 D9902 ( .Y(D9902_Y), .B(D8663_Y), .A(D9899_Y));
KC_NAND2_X2 D9713 ( .Y(D9713_Y), .B(D8478_Y), .A(D9700_Y));
KC_NAND2_X2 D8590 ( .Y(D8590_Y), .B(D8607_Y), .A(D8579_Y));
KC_NAND2_X2 D8587 ( .Y(D8587_Y), .B(D8607_Y), .A(D8569_Y));
KC_NAND2_X2 D8464 ( .Y(D8464_Y), .B(D8415_Y), .A(D8418_Y));
KC_NAND2_X2 D8462 ( .Y(D8462_Y), .B(D8478_Y), .A(D8453_Y));
KC_NAND2_X2 D8461 ( .Y(D8461_Y), .B(D8286_Y), .A(D8279_Y));
KC_NAND2_X2 D6665 ( .Y(D6665_Y), .B(D16753_Y), .A(GND));
KC_NAND2_X2 D6653 ( .Y(D6653_Y), .B(D16753_Y), .A(D6646_Y));
KC_NAND2_X2 D6543 ( .Y(D6543_Y), .B(D16696_Y), .A(D6522_Y));
KC_NAND2_X2 D6542 ( .Y(D6542_Y), .B(D16696_Y), .A(D6520_Y));
KC_NAND2_X2 D6380 ( .Y(D6380_Y), .B(D14591_Y), .A(D6372_Y));
KC_NAND2_X2 D6379 ( .Y(D6379_Y), .B(D14591_Y), .A(D6373_Y));
KC_NAND2_X2 D5803 ( .Y(D5803_Y), .B(D6275_Y), .A(D224_Y));
KC_NAND2_X2 D5802 ( .Y(D5802_Y), .B(D6275_Y), .A(D185_Y));
KC_NAND2_X2 D5478 ( .Y(D5478_Y), .B(D5489_Y), .A(D5460_Y));
KC_NAND2_X2 D5475 ( .Y(D5475_Y), .B(D5489_Y), .A(D5459_Y));
KC_NAND2_X2 D5079 ( .Y(D5079_Y), .B(D3501_Y), .A(D4985_Y));
KC_NAND2_X2 D4845 ( .Y(D4845_Y), .B(D4819_Q), .A(D3383_Q));
KC_NAND2_X2 D4725 ( .Y(D4725_Y), .B(D6197_Y), .A(D4716_Y));
KC_NAND2_X2 D4632 ( .Y(D4632_Y), .B(D6197_Y), .A(D4618_Y));
KC_NAND2_X2 D4480 ( .Y(D4480_Y), .B(D6128_Y), .A(D4459_Y));
KC_NAND2_X2 D4044 ( .Y(D4044_Y), .B(D4072_Y), .A(D4039_Y));
KC_NAND2_X2 D4043 ( .Y(D4043_Y), .B(D4072_Y), .A(D4034_Y));
KC_NAND2_X2 D4017 ( .Y(D4017_Y), .B(D4571_Y), .A(D1460_Y));
KC_NAND2_X2 D3971 ( .Y(D3971_Y), .B(D4571_Y), .A(D3958_Y));
KC_NAND2_X2 D3732 ( .Y(D3732_Y), .B(D4406_Y), .A(D3719_Y));
KC_NAND2_X2 D3731 ( .Y(D3731_Y), .B(D4406_Y), .A(D3718_Y));
KC_NAND2_X2 D3295 ( .Y(D3295_Y), .B(D3266_Y), .A(D3265_Y));
KC_NAND2_X2 D2695 ( .Y(D2695_Y), .B(D16715_Y), .A(D2694_Y));
KC_NAND2_X2 D1647 ( .Y(D1647_Y), .B(D6128_Y), .A(D1625_Y));
KC_TINV_X1 D8267 ( .Y(D8267_Y), .A(D616_Y), .OE(D101_Y));
KC_TINV_X1 D6286 ( .Y(D6286_Y), .A(D16147_Y), .OE(D7547_Y));
KC_TINV_X1 D5949 ( .Y(D5949_Y), .A(D5937_Y), .OE(D6186_Y));
KC_TINV_X1 D5640 ( .Y(D5640_Y), .A(D4037_Y), .OE(D5556_Y));
KC_TINV_X1 D3599 ( .Y(D3599_Y), .A(D3586_Y), .OE(D3481_Q));
KC_TINV_X1 D1825 ( .Y(D1825_Y), .A(D6268_Y), .OE(D1815_Y));
KC_TINV_X1 D1537 ( .Y(D1537_Y), .A(D4966_Y), .OE(D1527_Q));
KC_INV_X6 D16726 ( .Y(D16726_Y), .A(D2695_Y));
KC_INV_X6 D16721 ( .Y(D16721_Y), .A(D16722_Y));
KC_INV_X6 D16699 ( .Y(D16699_Y), .A(D16700_Y));
KC_INV_X6 D16698 ( .Y(D16698_Y), .A(D16701_Y));
KC_INV_X6 D16637 ( .Y(D16637_Y), .A(D16632_Y));
KC_INV_X6 D16621 ( .Y(D16621_Y), .A(D16615_Y));
KC_INV_X6 D16584 ( .Y(D16584_Y), .A(D16578_Y));
KC_INV_X6 D16577 ( .Y(D16577_Y), .A(D16576_Y));
KC_INV_X6 D16312 ( .Y(D16312_Y), .A(D16313_Y));
KC_INV_X6 D16311 ( .Y(D16311_Y), .A(D16308_Y));
KC_INV_X6 D15130 ( .Y(D15130_Y), .A(D15131_Y));
KC_INV_X6 D15129 ( .Y(D15129_Y), .A(D15132_Y));
KC_INV_X6 D14784 ( .Y(D14784_Y), .A(D14681_Y));
KC_INV_X6 D14680 ( .Y(D14680_Y), .A(D14682_Y));
KC_INV_X6 D13822 ( .Y(D13822_Y), .A(D13824_Y));
KC_INV_X6 D13821 ( .Y(D13821_Y), .A(D13823_Y));
KC_INV_X6 D13608 ( .Y(D13608_Y), .A(D13609_Y));
KC_INV_X6 D13606 ( .Y(D13606_Y), .A(D13607_Y));
KC_INV_X6 D13084 ( .Y(D13084_Y), .A(D13089_Y));
KC_INV_X6 D12338 ( .Y(D12338_Y), .A(D12272_Y));
KC_INV_X6 D12271 ( .Y(D12271_Y), .A(D12269_Y));
KC_INV_X6 D12176 ( .Y(D12176_Y), .A(D13847_Y));
KC_INV_X6 D12175 ( .Y(D12175_Y), .A(D10821_Y));
KC_INV_X6 D12118 ( .Y(D12118_Y), .A(D12123_Y));
KC_INV_X6 D11660 ( .Y(D11660_Y), .A(D4747_Y));
KC_INV_X6 D11657 ( .Y(D11657_Y), .A(D392_Y));
KC_INV_X6 D11655 ( .Y(D11655_Y), .A(D6281_Y));
KC_INV_X6 D11628 ( .Y(D11628_Y), .A(D10187_Y));
KC_INV_X6 D11596 ( .Y(D11596_Y), .A(D11597_Y));
KC_INV_X6 D11332 ( .Y(D11332_Y), .A(D11334_Y));
KC_INV_X6 D11331 ( .Y(D11331_Y), .A(D11333_Y));
KC_INV_X6 D11032 ( .Y(D11032_Y), .A(D11036_Y));
KC_INV_X6 D11028 ( .Y(D11028_Y), .A(D11029_Y));
KC_INV_X6 D10798 ( .Y(D10798_Y), .A(D10799_Y));
KC_INV_X6 D10797 ( .Y(D10797_Y), .A(D7757_Y));
KC_INV_X6 D10795 ( .Y(D10795_Y), .A(D10796_Y));
KC_INV_X6 D10794 ( .Y(D10794_Y), .A(D7756_Y));
KC_INV_X6 D10514 ( .Y(D10514_Y), .A(D6793_Y));
KC_INV_X6 D10291 ( .Y(D10291_Y), .A(D1976_Y));
KC_INV_X6 D10216 ( .Y(D10216_Y), .A(D6405_Y));
KC_INV_X6 D10133 ( .Y(D10133_Y), .A(D10069_Y));
KC_INV_X6 D10044 ( .Y(D10044_Y), .A(D8898_Q));
KC_INV_X6 D10043 ( .Y(D10043_Y), .A(D8895_Q));
KC_INV_X6 D10028 ( .Y(D10028_Y), .A(D10006_Q));
KC_INV_X6 D10027 ( .Y(D10027_Y), .A(D10008_Q));
KC_INV_X6 D9907 ( .Y(D9907_Y), .A(D9904_Y));
KC_INV_X6 D9901 ( .Y(D9901_Y), .A(D9902_Y));
KC_INV_X6 D9716 ( .Y(D9716_Y), .A(D8462_Y));
KC_INV_X6 D9715 ( .Y(D9715_Y), .A(D9713_Y));
KC_INV_X6 D9266 ( .Y(D9266_Y), .A(D13287_Y));
KC_INV_X6 D9017 ( .Y(D9017_Y), .A(D8896_Q));
KC_INV_X6 D9016 ( .Y(D9016_Y), .A(D326_Q));
KC_INV_X6 D9015 ( .Y(D9015_Y), .A(D8897_Q));
KC_INV_X6 D9014 ( .Y(D9014_Y), .A(D9023_Q));
KC_INV_X6 D9013 ( .Y(D9013_Y), .A(D305_Q));
KC_INV_X6 D9012 ( .Y(D9012_Y), .A(D2090_Q));
KC_INV_X6 D8949 ( .Y(D8949_Y), .A(D303_Q));
KC_INV_X6 D8948 ( .Y(D8948_Y), .A(D8955_Q));
KC_INV_X6 D8815 ( .Y(D8815_Y), .A(D147_Q));
KC_INV_X6 D8592 ( .Y(D8592_Y), .A(D8590_Y));
KC_INV_X6 D8586 ( .Y(D8586_Y), .A(D8587_Y));
KC_INV_X6 D8542 ( .Y(D8542_Y), .A(D8466_Y));
KC_INV_X6 D8540 ( .Y(D8540_Y), .A(D5461_Y));
KC_INV_X6 D8146 ( .Y(D8146_Y), .A(D6759_Y));
KC_INV_X6 D7992 ( .Y(D7992_Y), .A(D7936_Y));
KC_INV_X6 D7989 ( .Y(D7989_Y), .A(D8466_Y));
KC_INV_X6 D7784 ( .Y(D7784_Y), .A(D13285_Y));
KC_INV_X6 D7783 ( .Y(D7783_Y), .A(D7819_Y));
KC_INV_X6 D7782 ( .Y(D7782_Y), .A(D1772_Y));
KC_INV_X6 D7470 ( .Y(D7470_Y), .A(D7319_Y));
KC_INV_X6 D7469 ( .Y(D7469_Y), .A(D5704_Y));
KC_INV_X6 D6664 ( .Y(D6664_Y), .A(D6665_Y));
KC_INV_X6 D6654 ( .Y(D6654_Y), .A(D6653_Y));
KC_INV_X6 D6545 ( .Y(D6545_Y), .A(D6543_Y));
KC_INV_X6 D6541 ( .Y(D6541_Y), .A(D6542_Y));
KC_INV_X6 D6378 ( .Y(D6378_Y), .A(D6379_Y));
KC_INV_X6 D6377 ( .Y(D6377_Y), .A(D6380_Y));
KC_INV_X6 D6262 ( .Y(D6262_Y), .A(D4725_Y));
KC_INV_X6 D6177 ( .Y(D6177_Y), .A(D346_Y));
KC_INV_X6 D5801 ( .Y(D5801_Y), .A(D5803_Y));
KC_INV_X6 D5681 ( .Y(D5681_Y), .A(D5802_Y));
KC_INV_X6 D5477 ( .Y(D5477_Y), .A(D5478_Y));
KC_INV_X6 D5473 ( .Y(D5473_Y), .A(D5475_Y));
KC_INV_X6 D5403 ( .Y(D5403_Y), .A(D5392_Y));
KC_INV_X6 D4960 ( .Y(D4960_Y), .A(D3400_Y));
KC_INV_X6 D4811 ( .Y(D4811_Y), .A(D3163_Y));
KC_INV_X6 D4479 ( .Y(D4479_Y), .A(D4480_Y));
KC_INV_X6 D4478 ( .Y(D4478_Y), .A(D1647_Y));
KC_INV_X6 D4084 ( .Y(D4084_Y), .A(D4043_Y));
KC_INV_X6 D4046 ( .Y(D4046_Y), .A(D4044_Y));
KC_INV_X6 D3970 ( .Y(D3970_Y), .A(D3971_Y));
KC_INV_X6 D3730 ( .Y(D3730_Y), .A(D3731_Y));
KC_INV_X6 D3729 ( .Y(D3729_Y), .A(D3732_Y));
KC_INV_X6 D3371 ( .Y(D3371_Y), .A(D3479_Y));
KC_INV_X6 D2386 ( .Y(D2386_Y), .A(D13085_Y));
KC_INV_X6 D2343 ( .Y(D2343_Y), .A(D7668_Y));
KC_INV_X6 D2222 ( .Y(D2222_Y), .A(D545_Y));
KC_INV_X6 D2160 ( .Y(D2160_Y), .A(D230_Q));
KC_INV_X6 D2158 ( .Y(D2158_Y), .A(D2175_Q));
KC_INV_X6 D2086 ( .Y(D2086_Y), .A(D272_Y));
KC_INV_X6 D1932 ( .Y(D1932_Y), .A(D545_Y));
KC_INV_X6 D20 ( .Y(D20_Y), .A(D235_Y));
KC_INV_X6 D1787 ( .Y(D1787_Y), .A(D4150_Y));
KC_INV_X6 D1646 ( .Y(D1646_Y), .A(D4632_Y));
KC_INV_X6 D1492 ( .Y(D1492_Y), .A(D4017_Y));
KC_INV_X7 D16732 ( .Y(D16732_Y), .A(D16731_Y));
KC_INV_X7 D16724 ( .Y(D16724_Y), .A(D1328_Y));
KC_INV_X7 D16707 ( .Y(D16707_Y), .A(D16711_Y));
KC_INV_X7 D16683 ( .Y(D16683_Y), .A(D1329_Y));
KC_INV_X7 D16628 ( .Y(D16628_Y), .A(D16636_Y));
KC_INV_X7 D16619 ( .Y(D16619_Y), .A(D16618_Y));
KC_INV_X7 D16585 ( .Y(D16585_Y), .A(D1389_Y));
KC_INV_X7 D16553 ( .Y(D16553_Y), .A(D16554_Y));
KC_INV_X7 D16326 ( .Y(D16326_Y), .A(D16404_Y));
KC_INV_X7 D16325 ( .Y(D16325_Y), .A(D16405_Y));
KC_INV_X7 D15142 ( .Y(D15142_Y), .A(D15154_Y));
KC_INV_X7 D15135 ( .Y(D15135_Y), .A(D15155_Y));
KC_INV_X7 D14791 ( .Y(D14791_Y), .A(D14800_Y));
KC_INV_X7 D14697 ( .Y(D14697_Y), .A(D14801_Y));
KC_INV_X7 D13832 ( .Y(D13832_Y), .A(D1397_Y));
KC_INV_X7 D13830 ( .Y(D13830_Y), .A(D13838_Y));
KC_INV_X7 D13615 ( .Y(D13615_Y), .A(D13623_Y));
KC_INV_X7 D13612 ( .Y(D13612_Y), .A(D13618_Y));
KC_INV_X7 D12548 ( .Y(D12548_Y), .A(D1244_Y));
KC_INV_X7 D12511 ( .Y(D12511_Y), .A(D12513_Y));
KC_INV_X7 D12293 ( .Y(D12293_Y), .A(D12288_Y));
KC_INV_X7 D12284 ( .Y(D12284_Y), .A(D12292_Y));
KC_INV_X7 D11603 ( .Y(D11603_Y), .A(D11607_Y));
KC_INV_X7 D11598 ( .Y(D11598_Y), .A(D12126_Y));
KC_INV_X7 D11407 ( .Y(D11407_Y), .A(D2257_Y));
KC_INV_X7 D11347 ( .Y(D11347_Y), .A(D941_Y));
KC_INV_X7 D11041 ( .Y(D11041_Y), .A(D11047_Y));
KC_INV_X7 D11037 ( .Y(D11037_Y), .A(D2228_Y));
KC_INV_X7 D10814 ( .Y(D10814_Y), .A(D10827_Y));
KC_INV_X7 D10810 ( .Y(D10810_Y), .A(D10820_Y));
KC_INV_X7 D9914 ( .Y(D9914_Y), .A(D9920_Y));
KC_INV_X7 D9720 ( .Y(D9720_Y), .A(D160_Y));
KC_INV_X7 D8660 ( .Y(D8660_Y), .A(D9919_Y));
KC_INV_X7 D8468 ( .Y(D8468_Y), .A(D1058_Y));
KC_INV_X7 D7015 ( .Y(D7015_Y), .A(D7019_Y));
KC_INV_X7 D6682 ( .Y(D6682_Y), .A(D713_Y));
KC_INV_X7 D6680 ( .Y(D6680_Y), .A(D712_Y));
KC_INV_X7 D6565 ( .Y(D6565_Y), .A(D6561_Y));
KC_INV_X7 D6558 ( .Y(D6558_Y), .A(D6564_Y));
KC_INV_X7 D6395 ( .Y(D6395_Y), .A(D6398_Y));
KC_INV_X7 D6388 ( .Y(D6388_Y), .A(D6412_Y));
KC_INV_X7 D6121 ( .Y(D6121_Y), .A(D6126_Y));
KC_INV_X7 D6074 ( .Y(D6074_Y), .A(D1807_Y));
KC_INV_X7 D5696 ( .Y(D5696_Y), .A(D5700_Y));
KC_INV_X7 D5695 ( .Y(D5695_Y), .A(D5811_Y));
KC_INV_X7 D5486 ( .Y(D5486_Y), .A(D1662_Y));
KC_INV_X7 D5483 ( .Y(D5483_Y), .A(D5487_Y));
KC_INV_X7 D4646 ( .Y(D4646_Y), .A(D4648_Y));
KC_INV_X7 D4055 ( .Y(D4055_Y), .A(D4087_Y));
KC_INV_X7 D4052 ( .Y(D4052_Y), .A(D4067_Y));
KC_INV_X7 D4021 ( .Y(D4021_Y), .A(D4025_Y));
KC_INV_X7 D3982 ( .Y(D3982_Y), .A(D3984_Y));
KC_INV_X7 D3760 ( .Y(D3760_Y), .A(D3759_Y));
KC_INV_X7 D3751 ( .Y(D3751_Y), .A(D711_Y));
KC_INV_X7 D1656 ( .Y(D1656_Y), .A(D362_Y));
KC_INV_X7 D1238 ( .Y(D1238_Y), .A(D1240_Y));
KC_TIEHI_X1 D16715 ( .Y(D16715_Y));
KC_TIEHI_X1 D16772 ( .Y(D16772_Y));
KC_TIEHI_X1 D16639 ( .Y(D16639_Y));
KC_TIEHI_X1 D16588 ( .Y(D16588_Y));
KC_TIEHI_X1 D16341 ( .Y(D16341_Y));
KC_TIEHI_X1 D15159 ( .Y(D15159_Y));
KC_TIEHI_X1 D14712 ( .Y(D14712_Y));
KC_TIEHI_X1 D13843 ( .Y(D13843_Y));
KC_TIEHI_X1 D13094 ( .Y(D13094_Y));
KC_TIEHI_X1 D12304 ( .Y(D12304_Y));
KC_TIEHI_X1 D16761 ( .Y(D16761_Y));
KC_TIEHI_X1 D11612 ( .Y(D11612_Y));
KC_TIEHI_X1 D11417 ( .Y(D11417_Y));
KC_TIEHI_X1 D11055 ( .Y(D11055_Y));
KC_TIEHI_X1 D16082 ( .Y(D16082_Y));
KC_TIEHI_X1 D10313 ( .Y(D10313_Y));
KC_TIEHI_X1 D8663 ( .Y(D8663_Y));
KC_TIEHI_X1 D8607 ( .Y(D8607_Y));
KC_TIEHI_X1 D8478 ( .Y(D8478_Y));
KC_TIEHI_X1 D8359 ( .Y(D8359_Y));
KC_TIEHI_X1 D16753 ( .Y(D16753_Y));
KC_TIEHI_X1 D16696 ( .Y(D16696_Y));
KC_TIEHI_X1 D14591 ( .Y(D14591_Y));
KC_TIEHI_X1 D6275 ( .Y(D6275_Y));
KC_TIEHI_X1 D5489 ( .Y(D5489_Y));
KC_TIEHI_X1 D6197 ( .Y(D6197_Y));
KC_TIEHI_X1 D6128 ( .Y(D6128_Y));
KC_TIEHI_X1 D4072 ( .Y(D4072_Y));
KC_TIEHI_X1 D4571 ( .Y(D4571_Y));
KC_TIEHI_X1 D4406 ( .Y(D4406_Y));
KC_TIEHI_X1 D1076 ( .Y(D1076_Y));
KC_NOR4_X1 D16000 ( .Y(D16000_Y), .D(D16013_Q), .C(D15999_Q),     .B(D16012_Q), .A(D15997_Q));
KC_NOR4_X1 D14476 ( .Y(D14476_Y), .D(D1383_Q), .C(D14496_Q),     .B(D15235_Q), .A(D1379_Q));
KC_NOR4_X1 D14193 ( .Y(D14193_Y), .D(D14196_Q), .C(D926_Q),     .B(D14164_Q), .A(D14167_Q));
KC_NOR4_X1 D9387 ( .Y(D9387_Y), .D(D266_Y), .C(D16_Y), .B(D11660_Y),     .A(D10177_Y));
KC_NOR4_X1 D4836 ( .Y(D4836_Y), .D(D4825_Q), .C(D4817_Q), .B(D4824_Q),     .A(D1654_Q));
KC_NOR4_X1 D2584 ( .Y(D2584_Y), .D(D145_Q), .C(D925_Q), .B(D14874_Q),     .A(D15670_Q));
KC_NOR4_X1 D1525 ( .Y(D1525_Y), .D(D2672_Y), .C(D2851_Y), .B(D2814_Q),     .A(D1524_Q));
KC_NOR4_X1 D1075 ( .Y(D1075_Y), .D(D16319_Q), .C(D15797_Q),     .B(D15711_Q), .A(D1074_Q));
KC_OAI31_X3 D7984 ( .A2(D7973_Q), .A1(D6381_Q), .Y(D7984_Y),     .A0(D7653_Y), .B(D1849_Y));
KC_OAI31_X3 D1073 ( .A2(D13575_Y), .A1(D13569_Y), .Y(D1073_Y),     .A0(D13409_Y), .B(D2426_Y));
KC_OAI31_X2 D16295 ( .B2(D16271_Y), .B1(D16285_Y), .B0(D16279_Y),     .Y(D16295_Y), .A(D16249_Y));
KC_OAI31_X2 D13710 ( .B2(D85_Y), .B1(D13649_Y), .B0(D13409_Y),     .Y(D13710_Y), .A(D13547_Y));
KC_OAI31_X2 D8258 ( .B2(D8185_Y), .B1(D9369_Y), .B0(D9365_Y),     .Y(D8258_Y), .A(D8029_Y));
KC_OAI31_X2 D2477 ( .B2(D13565_Y), .B1(D13579_Y), .B0(D13409_Y),     .Y(D2477_Y), .A(D13546_Y));
KC_OAI31_X2 D2476 ( .B2(D13624_Y), .B1(D13559_Y), .B0(D13409_Y),     .Y(D2476_Y), .A(D13555_Y));
KC_OAI31_X2 D2475 ( .B2(D13416_Y), .B1(D13420_Y), .B0(D13409_Y),     .Y(D2475_Y), .A(D13429_Y));
KC_OAI31_X2 D2260 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11552_Y),     .Y(D2260_Y), .A(D11536_Y));
KC_OAI31_X2 D1330 ( .B2(D2243_Y), .B1(D11565_Y), .B0(D11505_Y),     .Y(D1330_Y), .A(D11536_Y));
KC_OAI31_X2 D1071 ( .B2(D13551_Y), .B1(D13544_Y), .B0(D13409_Y),     .Y(D1071_Y), .A(D13554_Y));
KC_ADDF_X1 D16350 ( .S(D16350_S), .Ci(D1000_S), .B(D16363_Q),     .A(D16347_Y));
KC_ADDF_X1 D16306 ( .S(D16306_S), .Ci(D15778_S), .B(D16346_Q),     .A(D16305_Y));
KC_ADDF_X1 D15942 ( .S(D15942_S), .Ci(D15933_Y), .B(D16390_Q),     .A(D15913_Y));
KC_ADDF_X1 D15939 ( .S(D15939_S), .Ci(D15938_Y), .B(D16391_Q),     .A(D15909_Y));
KC_ADDF_X1 D15937 ( .S(D15937_S), .Ci(D15940_Y), .B(D16364_Q),     .A(D2596_Y));
KC_ADDF_X1 D15936 ( .S(D15936_S), .Ci(D15922_Y), .B(D15910_Y),     .A(D1234_Q));
KC_ADDF_X1 D15935 ( .S(D15935_S), .Ci(D15932_Y), .B(D16389_Q),     .A(D15895_Y));
KC_ADDF_X1 D15862 ( .S(D15862_S), .Ci(D15826_Y), .B(D16359_Q),     .A(D15781_S));
KC_ADDF_X1 D15861 ( .S(D15861_S), .Ci(D15780_S), .B(D15823_Y),     .A(D15868_Q));
KC_ADDF_X1 D15860 ( .S(D15860_S), .Ci(D15821_Y), .B(D16353_Q),     .A(D16306_S));
KC_ADDF_X1 D15859 ( .S(D15859_S), .Ci(D2567_S), .B(D15818_Y),     .A(D15870_Q));
KC_ADDF_X1 D15858 ( .S(D15858_S), .Ci(D15862_S), .B(D15829_Y),     .A(D1148_Q));
KC_ADDF_X1 D15857 ( .S(D15857_S), .Ci(D15810_Y), .B(D16350_S),     .A(D16355_Q));
KC_ADDF_X1 D15856 ( .S(D15856_S), .Ci(D15860_S), .B(D15831_Y),     .A(D16357_Q));
KC_ADDF_X1 D15785 ( .S(D15785_S), .Ci(D2632_Y), .B(D2603_Y),     .A(D1074_Q));
KC_ADDF_X1 D15783 ( .S(D15783_S), .Ci(D15784_Y), .B(D15735_Y),     .A(D15797_Q));
KC_ADDF_X1 D15782 ( .S(D15782_S), .Ci(D15740_Y), .B(D1053_Q),     .A(D15739_Y));
KC_ADDF_X1 D15781 ( .S(D15781_S), .Ci(D15783_S), .B(D15792_Q),     .A(D15720_Y));
KC_ADDF_X1 D15780 ( .S(D15780_S), .Ci(D15715_Y), .B(D16361_Q),     .A(D15779_S));
KC_ADDF_X1 D15779 ( .S(D15779_S), .Ci(D15785_S), .B(D15791_Q),     .A(D15729_Y));
KC_ADDF_X1 D15778 ( .S(D15778_S), .Ci(D15731_Y), .B(D15734_Y),     .A(D1077_Q));
KC_ADDF_X1 D15248 ( .S(D15248_S), .Ci(D15306_Y), .B(D15243_Y),     .A(D15242_Y));
KC_ADDF_X1 D15127 ( .S(D15127_S), .Ci(D15125_Y), .B(D16393_Q),     .A(D15102_Y));
KC_ADDF_X1 D15126 ( .S(D15126_S), .Ci(D2566_Y), .B(D16365_Q),     .A(D15048_Y));
KC_ADDF_X1 D15072 ( .S(D15072_S), .Ci(D14984_S), .B(D15032_Y),     .A(D1157_Q));
KC_ADDF_X1 D15071 ( .S(D15071_S), .Ci(D15069_Y), .B(D2678_Q),     .A(D15018_Y));
KC_ADDF_X1 D15070 ( .S(D15070_S), .Ci(D14982_S), .B(D15019_Y),     .A(D15084_Q));
KC_ADDF_X1 D15068 ( .S(D15068_S), .Ci(D14981_S), .B(D15025_Y),     .A(D1163_Q));
KC_ADDF_X1 D14993 ( .S(D14993_S), .Ci(D2536_Y), .B(D2539_Y),     .A(D14870_Q));
KC_ADDF_X1 D14990 ( .S(D14990_S), .Ci(D14991_Y), .B(D14941_Y),     .A(D15711_Q));
KC_ADDF_X1 D14989 ( .S(D14989_S), .Ci(D15006_Y), .B(D14947_Y),     .A(D14997_Q));
KC_ADDF_X1 D14988 ( .S(D14988_S), .Ci(D14993_S), .B(D14873_Q),     .A(D14933_Y));
KC_ADDF_X1 D14986 ( .S(D14986_S), .Ci(D14979_S), .B(D14996_Q),     .A(D14935_Y));
KC_ADDF_X1 D14984 ( .S(D14984_S), .Ci(D14922_Y), .B(D2516_Q),     .A(D14988_S));
KC_ADDF_X1 D14982 ( .S(D14982_S), .Ci(D14916_Y), .B(D2679_Q),     .A(D14986_S));
KC_ADDF_X1 D14981 ( .S(D14981_S), .Ci(D14915_Y), .B(D14304_Q),     .A(D14978_S));
KC_ADDF_X1 D14980 ( .S(D14980_S), .Ci(D14990_S), .B(D15793_Q),     .A(D14924_Y));
KC_ADDF_X1 D14979 ( .S(D14979_S), .Ci(D14945_Y), .B(D14928_Y),     .A(D15669_Q));
KC_ADDF_X1 D14978 ( .S(D14978_S), .Ci(D14989_S), .B(D1051_Q),     .A(D14934_Y));
KC_ADDF_X1 D13749 ( .S(D13749_S), .Ci(D14322_Y), .B(D13727_Y),     .A(D2468_Q));
KC_ADDF_X1 D13748 ( .S(D13748_S), .Ci(D14353_Y), .B(D2414_Y),     .A(D13765_Q));
KC_ADDF_X1 D13695 ( .S(D13695_S), .Ci(D13778_Y), .B(D13671_Y),     .A(D13705_Q));
KC_ADDF_X1 D13694 ( .S(D13694_S), .Ci(D14412_Y), .B(D13646_Y),     .A(D1150_Q));
KC_ADDF_X1 D13693 ( .S(D13693_S), .Ci(D13722_Y), .B(D13645_Y),     .A(D1159_Q));
KC_ADDF_X1 D9377 ( .S(D9377_S), .Ci(D9373_Y), .B(D9386_Y),     .A(D8946_Y));
KC_ADDF_X1 D8798 ( .S(D8798_S), .Ci(D8805_Y), .B(D8774_Y),     .A(D8816_Y));
KC_ADDF_X1 D8689 ( .S(D8689_S), .Ci(D8671_Y), .B(D8671_Y),     .A(D8685_Y));
KC_ADDF_X1 D7577 ( .S(D7577_S), .Ci(D7537_Y), .B(D7571_Y),     .A(D7578_Y));
KC_ADDF_X1 D6887 ( .S(D6887_S), .Ci(D6888_Y), .B(D6836_Y),     .A(D6879_Y));
KC_ADDF_X1 D5384 ( .S(D5384_S), .Ci(D5383_Y), .B(D5481_Y),     .A(D5404_Y));
KC_ADDF_X1 D5068 ( .S(D5068_S), .Ci(D466_Y), .B(D5096_Y), .A(D3633_Y));
KC_ADDF_X1 D4801 ( .S(D4801_S), .Ci(D4787_Y), .B(D4840_Y),     .A(D4769_Y));
KC_ADDF_X1 D4718 ( .S(D4718_S), .Ci(D3267_Y), .B(D2995_Y),     .A(D3274_Y));
KC_ADDF_X1 D3260 ( .S(D3260_S), .Ci(D3291_Y), .B(D3290_Y),     .A(D3223_Y));
KC_ADDF_X1 D3171 ( .S(D3171_S), .Ci(D3170_Y), .B(D3182_Y),     .A(D3122_Y));
KC_ADDF_X1 D2567 ( .S(D2567_S), .Ci(D15039_Y), .B(D1155_Q),     .A(D14980_S));
KC_ADDF_X1 D2457 ( .S(D2457_S), .Ci(D14403_Y), .B(D13673_Y),     .A(D13704_Q));
KC_ADDF_X1 D2456 ( .S(D2456_S), .Ci(D14483_Y), .B(D2413_Y),     .A(D1235_Q));
KC_ADDF_X1 D2145 ( .S(D2145_S), .Ci(D2135_Y), .B(D10860_Y),     .A(D10856_Y));
KC_ADDF_X1 D2060 ( .S(D2060_S), .Ci(D9554_Y), .B(D9496_Y),     .A(D9496_Y));
KC_ADDF_X1 D2057 ( .S(D2057_S), .Ci(D8817_Y), .B(D8807_Y),     .A(D8807_Y));
KC_ADDF_X1 D1914 ( .S(D1914_S), .Ci(D8368_Y), .B(D8414_Y),     .A(D1837_Y));
KC_ADDF_X1 D1000 ( .S(D1000_S), .Ci(D15745_Y), .B(D16315_Q),     .A(D15782_S));
KC_NAND4_X3 D16559 ( .Y(D16559_Y), .D(D16558_Q), .C(D16557_Q),     .B(D1381_Q), .A(D16539_Y));
KC_NAND4_X3 D16299 ( .Y(D16299_Y), .D(D15630_Y), .C(D16266_Y),     .B(D16273_Y), .A(D16292_Q));
KC_NAND4_X3 D14806 ( .Y(D14806_Y), .D(D14743_Y), .C(D15611_Y),     .B(D13325_Y), .A(D16271_Y));
KC_NAND4_X3 D7818 ( .Y(D7818_Y), .D(D7770_Y), .C(D7776_Y), .B(D723_Q),     .A(D13285_Y));
KC_NAND4_X3 D7750 ( .Y(D7750_Y), .D(D10161_Y), .C(D7784_Y),     .B(D13289_Y), .A(D723_Q));
KC_NAND4_X3 D5705 ( .Y(D5705_Y), .D(D5670_Y), .C(D5652_Y), .B(D5686_Q),     .A(D5691_Q));
KC_NAND4_X3 D5703 ( .Y(D5703_Y), .D(D5664_Y), .C(D5667_Y), .B(D5666_Y),     .A(D5691_Q));
KC_NAND4_X3 D14 ( .Y(D14_Y), .D(D4421_Y), .C(D1787_Y), .B(D4424_Y),     .A(D4418_Y));
KC_NAND4_X3 D3829 ( .Y(D3829_Y), .D(D3827_Y), .C(D3795_Y), .B(D3782_Y),     .A(D3793_Y));
KC_NAND4_X3 D955 ( .Y(D955_Y), .D(D15630_Y), .C(D16276_Y), .B(D1378_Q),     .A(D14686_Q));
KC_BUF_X9 D16554 ( .Y(D16554_Y), .A(D16580_Y));
KC_BUF_X9 D14801 ( .Y(D14801_Y), .A(D14792_Y));
KC_BUF_X9 D14800 ( .Y(D14800_Y), .A(D14793_Y));
KC_BUF_X9 D13618 ( .Y(D13618_Y), .A(D13613_Y));
KC_BUF_X9 D12288 ( .Y(D12288_Y), .A(D12365_Y));
KC_BUF_X9 D12126 ( .Y(D12126_Y), .A(D12125_Y));
KC_BUF_X9 D11047 ( .Y(D11047_Y), .A(D11040_Y));
KC_BUF_X9 D10820 ( .Y(D10820_Y), .A(D10812_Y));
KC_BUF_X9 D7019 ( .Y(D7019_Y), .A(D8600_Y));
KC_BUF_X9 D6561 ( .Y(D6561_Y), .A(D6559_Y));
KC_BUF_X9 D6412 ( .Y(D6412_Y), .A(D6393_Y));
KC_BUF_X9 D6398 ( .Y(D6398_Y), .A(D6396_Y));
KC_BUF_X9 D5811 ( .Y(D5811_Y), .A(D5809_Y));
KC_BUF_X9 D5487 ( .Y(D5487_Y), .A(D5484_Y));
KC_BUF_X9 D4123 ( .Y(D4123_Y), .A(D4312_Y));
KC_BUF_X9 D3087 ( .Y(D3087_Y), .A(D377_Y));
KC_BUF_X9 D2228 ( .Y(D2228_Y), .A(D11038_Y));
KC_BUF_X9 D1662 ( .Y(D1662_Y), .A(D1660_Y));
KC_BUF_X9 D1389 ( .Y(D1389_Y), .A(D16593_Y));
KC_BUF_X9 D1240 ( .Y(D1240_Y), .A(D8599_Y));
KC_BUF_X9 D1058 ( .Y(D1058_Y), .A(D9718_Y));
KC_BUF_X9 D942 ( .Y(D942_Y), .A(D9637_Q));
KC_BUF_X9 D941 ( .Y(D941_Y), .A(D935_Y));
KC_NOR3_X2 D16597 ( .B(D16598_Q), .Y(D16597_Y), .C(D16571_Y),     .A(D16590_Q));
KC_NOR3_X2 D16285 ( .B(D16256_Y), .Y(D16285_Y), .C(D16250_Y),     .A(D16265_Y));
KC_NOR3_X2 D13393 ( .B(D12756_Q), .Y(D13393_Y), .C(D13268_Q),     .A(D12814_Y));
KC_NOR3_X2 D12048 ( .B(D6793_Y), .Y(D12048_Y), .C(D12027_Y),     .A(D6791_Y));
KC_NOR3_X2 D12047 ( .B(D8222_Y), .Y(D12047_Y), .C(D12018_Y),     .A(D11990_Y));
KC_NOR3_X2 D11989 ( .B(D8222_Y), .Y(D11989_Y), .C(D11942_Y),     .A(D11969_Y));
KC_NOR3_X2 D11982 ( .B(D6793_Y), .Y(D11982_Y), .C(D11945_Y),     .A(D6791_Y));
KC_NOR3_X2 D11981 ( .B(D760_Y), .Y(D11981_Y), .C(D11940_Y),     .A(D2277_Y));
KC_NOR3_X2 D11007 ( .B(D6793_Y), .Y(D11007_Y), .C(D10967_Y),     .A(D6791_Y));
KC_NOR3_X2 D11006 ( .B(D8222_Y), .Y(D11006_Y), .C(D10966_Y),     .A(D10990_Y));
KC_NOR3_X2 D11005 ( .B(D760_Y), .Y(D11005_Y), .C(D10971_Y),     .A(D10985_Y));
KC_NOR3_X2 D11004 ( .B(D5376_Y), .Y(D11004_Y), .C(D10963_Y),     .A(D5377_Y));
KC_NOR3_X2 D11003 ( .B(D760_Y), .Y(D11003_Y), .C(D10975_Y),     .A(D10985_Y));
KC_NOR3_X2 D10806 ( .B(D6793_Y), .Y(D10806_Y), .C(D10734_Y),     .A(D6791_Y));
KC_NOR3_X2 D10805 ( .B(D760_Y), .Y(D10805_Y), .C(D10728_Y),     .A(D10765_Y));
KC_NOR3_X2 D10804 ( .B(D8222_Y), .Y(D10804_Y), .C(D10730_Y),     .A(D10766_Y));
KC_NOR3_X2 D10516 ( .B(D6793_Y), .Y(D10516_Y), .C(D10965_Y),     .A(D6791_Y));
KC_NOR3_X2 D8340 ( .B(D8048_Y), .Y(D8340_Y), .C(D8288_Y), .A(D1920_Y));
KC_NOR3_X2 D8339 ( .B(D16755_Y), .Y(D8339_Y), .C(D8291_Y),     .A(D8047_Y));
KC_NOR3_X2 D8337 ( .B(D16755_Y), .Y(D8337_Y), .C(D8289_Y),     .A(D8047_Y));
KC_NOR3_X2 D7473 ( .B(D7418_Y), .Y(D7473_Y), .C(D7419_Y), .A(D6022_Y));
KC_NOR3_X2 D7295 ( .B(D5756_Y), .Y(D7295_Y), .C(D7279_Y), .A(D7097_Y));
KC_NOR3_X2 D6972 ( .B(D8222_Y), .Y(D6972_Y), .C(D6934_Y), .A(D5522_Y));
KC_NOR3_X2 D6971 ( .B(D6793_Y), .Y(D6971_Y), .C(D6935_Y), .A(D6791_Y));
KC_NOR3_X2 D5684 ( .B(D5662_Y), .Y(D5684_Y), .C(D5661_Y), .A(D5686_Q));
KC_NOR3_X2 D5540 ( .B(D760_Y), .Y(D5540_Y), .C(D5518_Y), .A(D1596_Y));
KC_NOR3_X2 D5409 ( .B(D6808_Y), .Y(D5409_Y), .C(D5358_Y), .A(D6809_Y));
KC_NOR3_X2 D5408 ( .B(D8222_Y), .Y(D5408_Y), .C(D5359_Y), .A(D5392_Y));
KC_NOR3_X2 D5407 ( .B(D760_Y), .Y(D5407_Y), .C(D5368_Y), .A(D8267_Y));
KC_NOR3_X2 D5406 ( .B(D5389_Y), .Y(D5406_Y), .C(D5357_Y), .A(D5388_Y));
KC_NOR3_X2 D5405 ( .B(D8222_Y), .Y(D5405_Y), .C(D5350_Y), .A(D5449_Y));
KC_NOR3_X2 D5323 ( .B(D5389_Y), .Y(D5323_Y), .C(D5267_Y), .A(D5388_Y));
KC_NOR3_X2 D5322 ( .B(D760_Y), .Y(D5322_Y), .C(D1556_Y), .A(D5301_Y));
KC_NOR3_X2 D3379 ( .B(D3318_Y), .Y(D3379_Y), .C(D3351_Y), .A(D3317_Y));
KC_NOR3_X2 D2301 ( .B(D760_Y), .Y(D2301_Y), .C(D11956_Y),     .A(D11438_Y));
KC_NOR3_X2 D2300 ( .B(D5376_Y), .Y(D2300_Y), .C(D11957_Y),     .A(D5377_Y));
KC_NOR3_X2 D2227 ( .B(D5376_Y), .Y(D2227_Y), .C(D10972_Y),     .A(D5377_Y));
KC_NOR3_X2 D1651 ( .B(D5389_Y), .Y(D1651_Y), .C(D5520_Y), .A(D5388_Y));
KC_NOR3_X2 D1144 ( .B(D8222_Y), .Y(D1144_Y), .C(D10467_Y),     .A(D10990_Y));
KC_NOR3_X2 D921 ( .B(D6808_Y), .Y(D921_Y), .C(D6782_Y), .A(D6809_Y));
KC_CELL_X1 D9301 ( .Y(D9301_Y), .A(D9316_Y), .B(D9212_QN),     .C(D9271_Y));
KC_CELL_X1 D3707 ( .Y(D3707_Y), .A(D15596_Y), .B(D15663_Y),     .C(D16383_Y));
KC_DFFRNHQ_X3 D10239 ( .Q(D10239_Q), .S0(D10209_Y), .D(D10221_Q),     .RN(D9381_Y), .CK(D10707_Y));
KC_DFFRNHQ_X3 D9493 ( .Q(D9493_Q), .S0(D9409_Y), .D(D9445_Y),     .RN(D9446_Y), .CK(D9321_Y));
KC_DFFRNHQ_X3 D9302 ( .Q(D9302_Q), .S0(D5966_Y), .D(D13859_Y),     .RN(D9271_Y), .CK(D9211_QN));
KC_DFFRNHQ_X3 D9231 ( .Q(D9231_Q), .S0(D5966_Y), .D(D9302_Q),     .RN(D9271_Y), .CK(D9211_QN));
KC_DFFRNHQ_X3 D7412 ( .Q(D7412_Q), .S0(D7363_Y), .D(D5698_Y),     .RN(D8894_Y), .CK(D4462_Y));
KC_DFFRNHQ_X3 D4568 ( .Q(D4568_Q), .S0(D4542_Y), .D(D4395_Y),     .RN(D1652_Y), .CK(D4462_Y));
KC_DFFRNHQ_X3 D4567 ( .Q(D4567_Q), .S0(D1624_Y), .D(D4395_Y),     .RN(D1652_Y), .CK(D4462_Y));
KC_DFFRNHQ_X3 D4566 ( .Q(D4566_Q), .S0(D4548_Y), .D(D4274_Y),     .RN(D1652_Y), .CK(D4462_Y));
KC_DFFRNHQ_X3 D4495 ( .Q(D4495_Q), .S0(D4451_Y), .D(D5936_Y),     .RN(D1652_Y), .CK(D5931_QN));
KC_DFFRNHQ_X3 D3302 ( .Q(D3302_Q), .S0(D3262_Y), .D(D3248_Y),     .RN(D4827_Y), .CK(D4799_Y));
KC_DFFRNHQ_X3 D2816 ( .Q(D2816_Q), .S0(D2763_Y), .D(D2752_Y),     .RN(D2882_Y), .CK(D2864_Y));
KC_DFFRNHQ_X3 D1536 ( .Q(D1536_Q), .S0(D1477_Y), .D(D1442_Y),     .RN(D2882_Y), .CK(D7712_Y));
KC_DFFRNHQ_X3 D857 ( .Q(D857_Q), .S0(D8175_Y), .D(D8359_Y),     .RN(D9562_Y), .CK(D7962_Y));
KC_OA22_X1 D12371 ( .A1(D12311_Y), .B0(D12345_Y), .B1(D12347_Y),     .A0(D12310_Y), .Y(D12371_Y));
KC_OA22_X1 D12307 ( .A1(D648_Y), .B0(D12251_Y), .B1(D12704_Y),     .A0(D12323_Y), .Y(D12307_Y));
KC_OA22_X1 D5093 ( .A1(D4866_Y), .B0(D5031_Y), .B1(D1564_Y),     .A0(D5023_Y), .Y(D5093_Y));
KC_OA22_X1 D5092 ( .A1(D3420_Y), .B0(D4865_Y), .B1(D5021_Y),     .A0(D5023_Y), .Y(D5092_Y));
KC_OA22_X1 D850 ( .A1(D11767_Y), .B0(D12361_Y), .B1(D12354_Y),     .A0(D12324_Y), .Y(D850_Y));
KC_AOI21B_X2 D16520 ( .A0N(D16519_Y), .A1(D16506_Y), .Y(D16520_Y),     .B(D16496_Y));
KC_AOI21B_X2 D16516 ( .A0N(D16518_Y), .A1(D16498_Y), .Y(D16516_Y),     .B(D16496_Y));
KC_AOI21B_X2 D16297 ( .A0N(D16269_Y), .A1(D2628_Y), .Y(D16297_Y),     .B(D16260_Y));
KC_AOI21B_X2 D16296 ( .A0N(D16288_Q), .A1(D16299_Y), .Y(D16296_Y),     .B(D16251_Y));
KC_AOI21B_X2 D16227 ( .A0N(D2615_Y), .A1(D13374_Y), .Y(D16227_Y),     .B(D2658_Y));
KC_AOI21B_X2 D13637 ( .A0N(D13555_Y), .A1(D14236_Q), .Y(D13637_Y),     .B(D14074_Y));
KC_AOI21B_X2 D13527 ( .A0N(D14133_Y), .A1(D14025_Y), .Y(D13527_Y),     .B(D13472_Y));
KC_AOI21B_X2 D12297 ( .A0N(D12801_Y), .A1(D12362_Y), .Y(D12297_Y),     .B(D12657_Y));
KC_AOI21B_X2 D11675 ( .A0N(D11654_Y), .A1(D11649_Y), .Y(D11675_Y),     .B(D11654_Y));
KC_AOI21B_X2 D11674 ( .A0N(D11671_Y), .A1(D11646_Y), .Y(D11674_Y),     .B(D11654_Y));
KC_AOI21B_X2 D10831 ( .A0N(D10870_Y), .A1(D2223_Y), .Y(D10831_Y),     .B(D10807_Y));
KC_AOI21B_X2 D9593 ( .A0N(D2100_Y), .A1(D1665_Y), .Y(D9593_Y),     .B(D2102_Y));
KC_AOI21B_X2 D9489 ( .A0N(D9397_Y), .A1(D9443_Y), .Y(D9489_Y),     .B(D9403_Y));
KC_AOI21B_X2 D8731 ( .A0N(D8688_Y), .A1(D8691_Y), .Y(D8731_Y),     .B(D8675_Y));
KC_AOI21B_X2 D8729 ( .A0N(D8707_Y), .A1(D188_Y), .Y(D8729_Y),     .B(D8679_Y));
KC_AOI21B_X2 D8265 ( .A0N(D8243_Q), .A1(D8293_Y), .Y(D8265_Y),     .B(D8264_Y));
KC_AOI21B_X2 D7821 ( .A0N(D7762_Y), .A1(D447_Y), .Y(D7821_Y),     .B(D7792_Y));
KC_AOI21B_X2 D7616 ( .A0N(D7572_Y), .A1(D7639_Y), .Y(D7616_Y),     .B(D7569_Y));
KC_AOI21B_X2 D37 ( .A0N(D7514_Y), .A1(D1677_Y), .Y(D37_Y),     .B(D7567_Y));
KC_AOI21B_X2 D17 ( .A0N(D5959_Y), .A1(D7415_Y), .Y(D17_Y),     .B(D6014_Y));
KC_AOI21B_X2 D7406 ( .A0N(D7347_Y), .A1(D202_Y), .Y(D7406_Y),     .B(D7199_Y));
KC_AOI21B_X2 D7310 ( .A0N(D7200_Y), .A1(D7304_Y), .Y(D7310_Y),     .B(D7307_Y));
KC_AOI21B_X2 D6355 ( .A0N(D6295_Y), .A1(D10161_Y), .Y(D6355_Y),     .B(D6312_Y));
KC_AOI21B_X2 D6204 ( .A0N(D6145_Y), .A1(D6117_Y), .Y(D6204_Y),     .B(D6146_Y));
KC_AOI21B_X2 D5948 ( .A0N(D5905_Y), .A1(D5857_Y), .Y(D5948_Y),     .B(D7103_Y));
KC_AOI21B_X2 D4746 ( .A0N(D4673_Y), .A1(D4591_Y), .Y(D4746_Y),     .B(D3097_Y));
KC_AOI21B_X2 D4651 ( .A0N(D4817_Q), .A1(D47_Y), .Y(D4651_Y),     .B(D4613_Y));
KC_AOI21B_X2 D29 ( .A0N(D4466_Y), .A1(D4513_Y), .Y(D29_Y),     .B(D4518_Y));
KC_AOI21B_X2 D4399 ( .A0N(D4366_Y), .A1(D2956_Y), .Y(D4399_Y),     .B(D2829_Y));
KC_AOI21B_X2 D3202 ( .A0N(D3155_Y), .A1(D3180_Y), .Y(D3202_Y),     .B(D3195_Y));
KC_AOI21B_X2 D49 ( .A0N(D4615_Y), .A1(D310_Y), .Y(D49_Y), .B(D7641_Y));
KC_AOI21B_X2 D32 ( .A0N(D2948_Y), .A1(D2948_Y), .Y(D32_Y),     .B(D4525_Y));
KC_AOI21B_X2 D31 ( .A0N(D3045_Y), .A1(D316_Y), .Y(D31_Y), .B(D3034_Y));
KC_AOI21B_X2 D15 ( .A0N(D2911_Y), .A1(D2953_Y), .Y(D15_Y),     .B(D2953_Y));
KC_AOI21B_X2 D23 ( .A0N(D1905_Y), .A1(D5703_Y), .Y(D23_Y),     .B(D7507_Y));
KC_AOI21B_X2 D22 ( .A0N(D7505_Y), .A1(D5703_Y), .Y(D22_Y),     .B(D7507_Y));
KC_AOI21B_X2 D21 ( .A0N(D5960_Y), .A1(D1710_Y), .Y(D21_Y),     .B(D6083_Y));
KC_AOI21B_X2 D1672 ( .A0N(D4696_Y), .A1(D4572_Y), .Y(D1672_Y),     .B(D3097_Y));
KC_AOI21B_X2 D958 ( .A0N(D865_Y), .A1(D10859_Y), .Y(D958_Y),     .B(D2145_S));
KC_AOI21B_X2 D845 ( .A0N(D15534_Y), .A1(D15534_Y), .Y(D845_Y),     .B(D15582_Y));
KC_AOI21B_X2 D844 ( .A0N(D13363_Y), .A1(D819_Q), .Y(D844_Y),     .B(D13221_Y));
KC_AOI22B_X1 D15698 ( .A1(D15466_Y), .B0(D15485_Y), .B1(D15647_Y),     .Y(D15698_Y), .A0N(D15658_Y));
KC_AOI22B_X1 D15697 ( .A1(D15470_Y), .B0(D15484_Y), .B1(D14847_Y),     .Y(D15697_Y), .A0N(D15627_Y));
KC_AOI22B_X1 D15455 ( .A1(D15361_Y), .B0(D15378_Y), .B1(D15355_Y),     .Y(D15455_Y), .A0N(D15559_Y));
KC_AOI22B_X1 D15454 ( .A1(D15362_Y), .B0(D15367_Y), .B1(D15404_Y),     .Y(D15454_Y), .A0N(D15525_Y));
KC_AOI22B_X1 D15156 ( .A1(D16008_Q), .B0(D15996_Q), .B1(D15094_Y),     .Y(D15156_Y), .A0N(D16011_Q));
KC_AOI22B_X1 D15005 ( .A1(D14304_Q), .B0(D1054_Q), .B1(D14946_Y),     .Y(D15005_Y), .A0N(D2679_Q));
KC_AOI22B_X1 D14703 ( .A1(D14745_Y), .B0(D14655_Y), .B1(D14589_Y),     .Y(D14703_Y), .A0N(D14639_Y));
KC_AOI22B_X1 D14477 ( .A1(D1383_Q), .B0(D14419_Y), .B1(D14461_Y),     .Y(D14477_Y), .A0N(D15214_Q));
KC_AOI22B_X1 D14397 ( .A1(D1380_Q), .B0(D15871_Q), .B1(D15019_Y),     .Y(D14397_Y), .A0N(D16014_Q));
KC_AOI22B_X1 D14268 ( .A1(D14241_Q), .B0(D14302_Q), .B1(D14200_Y),     .Y(D14268_Y), .A0N(D14239_Q));
KC_AOI22B_X1 D14267 ( .A1(D14244_Q), .B0(D16314_Q), .B1(D14935_Y),     .Y(D14267_Y), .A0N(D1066_Q));
KC_AOI22B_X1 D14194 ( .A1(D14168_Q), .B0(D14091_Q), .B1(D14725_Y),     .Y(D14194_Y), .A0N(D14118_Q));
KC_AOI22B_X1 D14099 ( .A1(D14034_Y), .B0(D14038_Y), .B1(D14030_Y),     .Y(D14099_Y), .A0N(D14001_Y));
KC_AOI22B_X1 D14098 ( .A1(D14034_Y), .B0(D14038_Y), .B1(D14021_Y),     .Y(D14098_Y), .A0N(D14004_Y));
KC_AOI22B_X1 D13628 ( .A1(D11276_Y), .B0(D14247_Y), .B1(D15774_Y),     .Y(D13628_Y), .A0N(D2421_Y));
KC_AOI22B_X1 D13627 ( .A1(D11276_Y), .B0(D14247_Y), .B1(D15765_Y),     .Y(D13627_Y), .A0N(D2420_Y));
KC_AOI22B_X1 D13626 ( .A1(D11276_Y), .B0(D13540_Y), .B1(D15765_Y),     .Y(D13626_Y), .A0N(D2471_Y));
KC_AOI22B_X1 D13625 ( .A1(D11276_Y), .B0(D14220_Y), .B1(D15765_Y),     .Y(D13625_Y), .A0N(D13622_Y));
KC_AOI22B_X1 D13624 ( .A1(D12879_Y), .B0(D13393_Y), .B1(D12955_Y),     .Y(D13624_Y), .A0N(D13709_Y));
KC_AOI22B_X1 D13277 ( .A1(D14811_Y), .B0(D2454_Y), .B1(D12683_Q),     .Y(D13277_Y), .A0N(D13186_Y));
KC_AOI22B_X1 D9483 ( .A1(D8148_Q), .B0(D826_Q), .B1(D1986_Y),     .Y(D9483_Y), .A0N(D9405_Y));
KC_AOI22B_X1 D7978 ( .A1(D7921_Y), .B0(D7916_Y), .B1(D7907_Y),     .Y(D7978_Y), .A0N(D727_Y));
KC_AOI22B_X1 D5817 ( .A1(D5737_Y), .B0(D7193_Y), .B1(D9475_Y),     .Y(D5817_Y), .A0N(D1617_Y));
KC_AOI22B_X1 D5084 ( .A1(D1563_Y), .B0(D4877_Y), .B1(D3501_Y),     .Y(D5084_Y), .A0N(D3420_Y));
KC_AOI22B_X1 D2804 ( .A1(D2845_Y), .B0(D2746_Y), .B1(D2838_Y),     .Y(D2804_Y), .A0N(D2755_Y));
KC_AOI22B_X1 D1069 ( .A1(D11276_Y), .B0(D984_Y), .B1(D15774_Y),     .Y(D1069_Y), .A0N(D13641_Y));
KC_AOI22B_X1 D1068 ( .A1(D11276_Y), .B0(D13540_Y), .B1(D15774_Y),     .Y(D1068_Y), .A0N(D16767_Y));
KC_AOI22B_X1 D1067 ( .A1(D11276_Y), .B0(D984_Y), .B1(D15765_Y),     .Y(D1067_Y), .A0N(D13619_Y));
KC_AOI22B_X1 D948 ( .A1(D820_Q), .B0(D14118_Q), .B1(D14011_Y),     .Y(D948_Y), .A0N(D2517_Q));
KC_AOI22B_X1 D840 ( .A1(D13323_Y), .B0(D12748_Q), .B1(D13349_Y),     .Y(D840_Y), .A0N(D13380_Y));
KC_AOI22B_X1 D839 ( .A1(D14034_Y), .B0(D14038_Y), .B1(D14718_Y),     .Y(D839_Y), .A0N(D14087_Y));
KC_AOI22B_X1 D838 ( .A1(D14034_Y), .B0(D14038_Y), .B1(D14828_Y),     .Y(D838_Y), .A0N(D14088_Y));
KC_AND2_X3 D12057 ( .B(D12035_Y), .A(D11465_Y), .Y(D12057_Y));
KC_AND2_X3 D12056 ( .B(D2278_Y), .A(D11465_Y), .Y(D12056_Y));
KC_AND2_X3 D12055 ( .B(D12036_Y), .A(D11465_Y), .Y(D12055_Y));
KC_AND2_X3 D12054 ( .B(D12038_Y), .A(D11465_Y), .Y(D12054_Y));
KC_AND2_X3 D12053 ( .B(D12039_Y), .A(D11465_Y), .Y(D12053_Y));
KC_AND2_X3 D11995 ( .B(D11449_Y), .A(D2244_Y), .Y(D11995_Y));
KC_AND2_X3 D11994 ( .B(D11447_Y), .A(D11465_Y), .Y(D11994_Y));
KC_AND2_X3 D11993 ( .B(D1114_Y), .A(D11465_Y), .Y(D11993_Y));
KC_AND2_X3 D11992 ( .B(D11445_Y), .A(D11465_Y), .Y(D11992_Y));
KC_AND2_X3 D11586 ( .B(D11531_Y), .A(D11535_Y), .Y(D11586_Y));
KC_AND2_X3 D11477 ( .B(D11446_Y), .A(D11465_Y), .Y(D11477_Y));
KC_AND2_X3 D10824 ( .B(D10785_Y), .A(D11257_Y), .Y(D10824_Y));
KC_AND2_X3 D10823 ( .B(D10869_Y), .A(D11257_Y), .Y(D10823_Y));
KC_AND2_X3 D10563 ( .B(D9831_Y), .A(D8532_Y), .Y(D10563_Y));
KC_AND2_X3 D10562 ( .B(D1110_Y), .A(D8532_Y), .Y(D10562_Y));
KC_AND2_X3 D9360 ( .B(D12302_Y), .A(D9342_Y), .Y(D9360_Y));
KC_AND2_X3 D7018 ( .B(D6947_Y), .A(D6958_Y), .Y(D7018_Y));
KC_AND2_X3 D6909 ( .B(D6885_Y), .A(D8049_Y), .Y(D6909_Y));
KC_AND2_X3 D2303 ( .B(D2279_Y), .A(D11465_Y), .Y(D2303_Y));
KC_AND2_X3 D2302 ( .B(D2236_Y), .A(D11465_Y), .Y(D2302_Y));
KC_AND2_X3 D1956 ( .B(D8296_Y), .A(D8343_Q), .Y(D1956_Y));
KC_AND2_X3 D1955 ( .B(D1911_Y), .A(D8532_Y), .Y(D1955_Y));
KC_AND2_X3 D1161 ( .B(D11455_Y), .A(D2244_Y), .Y(D1161_Y));
KC_AND2_X3 D834 ( .B(D10781_Y), .A(D11257_Y), .Y(D834_Y));
KC_BUF_X8 D16581 ( .Y(D16581_Y), .A(D16587_QN));
KC_BUF_X8 D14177 ( .Y(D14177_Y), .A(D13249_Y));
KC_BUF_X8 D14095 ( .Y(D14095_Y), .A(D13249_Y));
KC_BUF_X8 D13276 ( .Y(D13276_Y), .A(D13249_Y));
KC_BUF_X8 D13205 ( .Y(D13205_Y), .A(D13249_Y));
KC_BUF_X8 D11633 ( .Y(D11633_Y), .A(D11641_Q));
KC_BUF_X8 D11632 ( .Y(D11632_Y), .A(D11632_A));
KC_BUF_X8 D11631 ( .Y(D11631_Y), .A(D11631_A));
KC_BUF_X8 D11630 ( .Y(D11630_Y), .A(D11637_Q));
KC_BUF_X8 D11133 ( .Y(D11133_Y), .A(D11124_Y));
KC_BUF_X8 D10187 ( .Y(D10187_Y), .A(D11625_Y));
KC_BUF_X8 D9985 ( .Y(D9985_Y), .A(D9947_Y));
KC_BUF_X8 D9474 ( .Y(D9474_Y), .A(D9359_Y));
KC_BUF_X8 D6076 ( .Y(D6076_Y), .A(D11630_Y));
KC_BUF_X8 D4965 ( .Y(D4965_Y), .A(D4958_QN));
KC_BUF_X8 D1947 ( .Y(D1947_Y), .A(D5812_Y));
KC_BUF_X8 D830 ( .Y(D830_Y), .A(D13249_Y));
KC_XOR2_X2 D15432 ( .Y(D15432_Y), .A(D16212_Y), .B(D16207_Y));
KC_XOR2_X2 D15431 ( .Y(D15431_Y), .A(D16210_Y), .B(D16213_Y));
KC_XOR2_X2 D15430 ( .Y(D15430_Y), .A(D16206_Y), .B(D16208_Y));
KC_XOR2_X2 D15325 ( .Y(D15325_Y), .A(D16218_Y), .B(D16220_Y));
KC_XOR2_X2 D15324 ( .Y(D15324_Y), .A(D16150_Y), .B(D16237_Y));
KC_XOR2_X2 D15318 ( .Y(D15318_Y), .A(D16162_Y), .B(D15447_Y));
KC_XOR2_X2 D15317 ( .Y(D15317_Y), .A(D16159_Y), .B(D16157_Y));
KC_XOR2_X2 D15315 ( .Y(D15315_Y), .A(D16149_Y), .B(D16221_Y));
KC_XOR2_X2 D14575 ( .Y(D14575_Y), .A(D16153_Y), .B(D16146_Y));
KC_XOR2_X2 D14574 ( .Y(D14574_Y), .A(D16152_Y), .B(D16183_Y));
KC_XOR2_X2 D14573 ( .Y(D14573_Y), .A(D16145_Y), .B(D16151_Y));
KC_XOR2_X2 D13381 ( .Y(D13381_Y), .A(D16073_Y), .B(D2669_Y));
KC_XOR2_X2 D13156 ( .Y(D13156_Y), .A(D16019_Y), .B(D15391_Y));
KC_XOR2_X2 D12139 ( .Y(D12139_Y), .A(D16038_Y), .B(D15392_Y));
KC_XOR2_X2 D10205 ( .Y(D10205_Y), .A(D16046_Y), .B(D15422_Y));
KC_XOR2_X2 D9087 ( .Y(D9087_Y), .A(D16039_Y), .B(D15419_Y));
KC_XOR2_X2 D9085 ( .Y(D9085_Y), .A(D16036_Y), .B(D15383_Y));
KC_XOR2_X2 D8998 ( .Y(D8998_Y), .A(D16021_Y), .B(D15382_Y));
KC_XOR2_X2 D8997 ( .Y(D8997_Y), .A(D16035_Y), .B(D15428_Y));
KC_XOR2_X2 D8902 ( .Y(D8902_Y), .A(D16018_Y), .B(D15312_Y));
KC_XOR2_X2 D8889 ( .Y(D8889_Y), .A(D16022_Y), .B(D15423_Y));
KC_XOR2_X2 D8888 ( .Y(D8888_Y), .A(D16034_Y), .B(D15396_Y));
KC_XOR2_X2 D8887 ( .Y(D8887_Y), .A(D505_Y), .B(D16048_Y));
KC_XOR2_X2 D8886 ( .Y(D8886_Y), .A(D16099_Y), .B(D15313_Y));
KC_XOR2_X2 D8885 ( .Y(D8885_Y), .A(D16076_Y), .B(D15268_Y));
KC_XOR2_X2 D6524 ( .Y(D6524_Y), .A(D16028_Y), .B(D15314_Y));
KC_XOR2_X2 D2871 ( .Y(D2871_Y), .A(D16020_Y), .B(D15299_Y));
KC_XOR2_X2 D2870 ( .Y(D2870_Y), .A(D16029_Y), .B(D15298_Y));
KC_XOR2_X2 D2866 ( .Y(D2866_Y), .A(D10206_Y), .B(D13189_Y));
KC_XOR2_X2 D2863 ( .Y(D2863_Y), .A(D12143_Q), .B(D12184_Y));
KC_XOR2_X2 D2862 ( .Y(D2862_Y), .A(D11276_Y), .B(D10216_Y));
KC_XOR2_X2 D2861 ( .Y(D2861_Y), .A(D8953_Q), .B(D7959_Y));
KC_XOR2_X2 D2665 ( .Y(D2665_Y), .A(D9021_Q), .B(D7957_Y));
KC_XOR2_X2 D2066 ( .Y(D2066_Y), .A(D7481_Q), .B(D7958_Y));
KC_XOR2_X2 D1476 ( .Y(D1476_Y), .A(D51_Y), .B(D8069_Y));
KC_XOR2_X2 D1475 ( .Y(D1475_Y), .A(D8895_Q), .B(D8869_Y));
KC_XOR2_X2 D1474 ( .Y(D1474_Y), .A(D3647_Q), .B(D727_Y));
KC_XOR2_X2 D1473 ( .Y(D1473_Y), .A(D2671_Y), .B(D2152_Y));
KC_XOR2_X2 D1472 ( .Y(D1472_Y), .A(D273_Y), .B(D7320_Y));
KC_XOR2_X2 D774 ( .Y(D774_Y), .A(D10681_Y), .B(D11228_Y));
KC_XOR2_X2 D651 ( .Y(D651_Y), .A(D16024_Y), .B(D15420_Y));
KC_BUF_X12 D15004 ( .Y(D15004_Y), .A(D833_Y));
KC_BUF_X12 D12860 ( .Y(D12860_Y), .A(D13249_Y));
KC_BUF_X12 D9359 ( .Y(D9359_Y), .A(D9347_Y));
KC_BUF_X12 D1059 ( .Y(D1059_Y), .A(D2522_Y));
KC_BUF_X12 D965 ( .Y(D965_Y), .A(D9360_Y));
KC_BUF_X12 D709 ( .Y(D709_Y), .A(D10706_Y));
KC_AND2_X2 D16716 ( .B(D16725_Y), .A(D16659_Y), .Y(D16716_Y));
KC_AND2_X2 D16705 ( .B(D16714_Y), .A(D16659_Y), .Y(D16705_Y));
KC_AND2_X2 D16629 ( .B(D16644_Y), .A(D16659_Y), .Y(D16629_Y));
KC_AND2_X2 D16567 ( .B(D16589_Y), .A(D16659_Y), .Y(D16567_Y));
KC_AND2_X2 D16321 ( .B(D16324_Y), .A(D12177_RN), .Y(D16321_Y));
KC_AND2_X2 D16294 ( .B(D16325_Y), .A(D16326_Y), .Y(D16294_Y));
KC_AND2_X2 D16167 ( .B(D16102_Y), .A(D16126_Y), .Y(D16167_Y));
KC_AND2_X2 D15259 ( .B(D15244_Y), .A(D15242_Y), .Y(D15259_Y));
KC_AND2_X2 D15144 ( .B(D15157_Y), .A(D14315_Y), .Y(D15144_Y));
KC_AND2_X2 D15143 ( .B(D15157_Y), .A(D14315_Y), .Y(D15143_Y));
KC_AND2_X2 D14693 ( .B(D14804_Y), .A(D14315_Y), .Y(D14693_Y));
KC_AND2_X2 D14691 ( .B(D14804_Y), .A(D14315_Y), .Y(D14691_Y));
KC_AND2_X2 D13399 ( .B(D13236_Y), .A(D10797_Y), .Y(D13399_Y));
KC_AND2_X2 D13091 ( .B(D13093_Y), .A(D14315_Y), .Y(D13091_Y));
KC_AND2_X2 D13052 ( .B(D13093_Y), .A(D14315_Y), .Y(D13052_Y));
KC_AND2_X2 D12998 ( .B(D13009_Y), .A(D14315_Y), .Y(D12998_Y));
KC_AND2_X2 D12364 ( .B(D12308_Y), .A(D11183_Y), .Y(D12364_Y));
KC_AND2_X2 D12287 ( .B(D850_Y), .A(D9345_Y), .Y(D12287_Y));
KC_AND2_X2 D12281 ( .B(D12308_Y), .A(D11183_Y), .Y(D12281_Y));
KC_AND2_X2 D11642 ( .B(D12748_Q), .A(D9345_Y), .Y(D11642_Y));
KC_AND2_X2 D11602 ( .B(D11611_Y), .A(D9850_Y), .Y(D11602_Y));
KC_AND2_X2 D11601 ( .B(D11611_Y), .A(D9850_Y), .Y(D11601_Y));
KC_AND2_X2 D11411 ( .B(D11418_Y), .A(D11183_Y), .Y(D11411_Y));
KC_AND2_X2 D11116 ( .B(D12371_Y), .A(D9345_Y), .Y(D11116_Y));
KC_AND2_X2 D11044 ( .B(D11054_Y), .A(D9850_Y), .Y(D11044_Y));
KC_AND2_X2 D11043 ( .B(D11054_Y), .A(D9850_Y), .Y(D11043_Y));
KC_AND2_X2 D10815 ( .B(D10829_Y), .A(D11183_Y), .Y(D10815_Y));
KC_AND2_X2 D10811 ( .B(D10829_Y), .A(D11183_Y), .Y(D10811_Y));
KC_AND2_X2 D10807 ( .B(D779_Y), .A(D779_Y), .Y(D10807_Y));
KC_AND2_X2 D9795 ( .B(D9774_Y), .A(D9781_Y), .Y(D9795_Y));
KC_AND2_X2 D9626 ( .B(D9721_Y), .A(D9850_Y), .Y(D9626_Y));
KC_AND2_X2 D9151 ( .B(D7630_Y), .A(D383_Y), .Y(D9151_Y));
KC_AND2_X2 D9024 ( .B(D8989_Y), .A(D8701_Y), .Y(D9024_Y));
KC_AND2_X2 D8826 ( .B(D8755_Y), .A(D7260_Y), .Y(D8826_Y));
KC_AND2_X2 D8661 ( .B(D8662_Y), .A(D9850_Y), .Y(D8661_Y));
KC_AND2_X2 D8601 ( .B(D8608_Y), .A(D9850_Y), .Y(D8601_Y));
KC_AND2_X2 D8597 ( .B(D8608_Y), .A(D9850_Y), .Y(D8597_Y));
KC_AND2_X2 D8155 ( .B(D8165_Y), .A(D11183_Y), .Y(D8155_Y));
KC_AND2_X2 D8154 ( .B(D8165_Y), .A(D11183_Y), .Y(D8154_Y));
KC_AND2_X2 D8059 ( .B(D8046_Y), .A(D8049_Y), .Y(D8059_Y));
KC_AND2_X2 D7796 ( .B(D7775_Y), .A(D7797_Y), .Y(D7796_Y));
KC_AND2_X2 D7738 ( .B(D6328_Y), .A(D7706_Y), .Y(D7738_Y));
KC_AND2_X2 D7392 ( .B(D5932_Y), .A(D7381_Y), .Y(D7392_Y));
KC_AND2_X2 D6614 ( .B(D8032_Y), .A(D8049_Y), .Y(D6614_Y));
KC_AND2_X2 D6613 ( .B(D6650_Y), .A(D8049_Y), .Y(D6613_Y));
KC_AND2_X2 D6390 ( .B(D6413_Y), .A(D11633_Y), .Y(D6390_Y));
KC_AND2_X2 D6389 ( .B(D6413_Y), .A(D11633_Y), .Y(D6389_Y));
KC_AND2_X2 D6206 ( .B(D1818_Y), .A(D6076_Y), .Y(D6206_Y));
KC_AND2_X2 D6122 ( .B(D30_Y), .A(D6076_Y), .Y(D6122_Y));
KC_AND2_X2 D6120 ( .B(D30_Y), .A(D6076_Y), .Y(D6120_Y));
KC_AND2_X2 D5808 ( .B(D5822_Y), .A(D6076_Y), .Y(D5808_Y));
KC_AND2_X2 D5807 ( .B(D5822_Y), .A(D6076_Y), .Y(D5807_Y));
KC_AND2_X2 D5411 ( .B(D5490_Y), .A(D11633_Y), .Y(D5411_Y));
KC_AND2_X2 D5410 ( .B(D5490_Y), .A(D11633_Y), .Y(D5410_Y));
KC_AND2_X2 D5248 ( .B(D5253_Y), .A(D11633_Y), .Y(D5248_Y));
KC_AND2_X2 D4642 ( .B(D1818_Y), .A(D6076_Y), .Y(D4642_Y));
KC_AND2_X2 D4395 ( .B(D4319_Y), .A(D5833_Y), .Y(D4395_Y));
KC_AND2_X2 D4061 ( .B(D4073_Y), .A(D9850_Y), .Y(D4061_Y));
KC_AND2_X2 D4059 ( .B(D4073_Y), .A(D9850_Y), .Y(D4059_Y));
KC_AND2_X2 D3983 ( .B(D1535_Y), .A(D11633_Y), .Y(D3983_Y));
KC_AND2_X2 D3191 ( .B(D3202_Y), .A(D4607_Y), .Y(D3191_Y));
KC_AND2_X2 D3085 ( .B(D3072_Y), .A(D3072_Y), .Y(D3085_Y));
KC_AND2_X2 D2693 ( .B(D16725_Y), .A(D16659_Y), .Y(D2693_Y));
KC_AND2_X2 D2692 ( .B(D16714_Y), .A(D16659_Y), .Y(D2692_Y));
KC_AND2_X2 D2689 ( .B(D16644_Y), .A(D16659_Y), .Y(D2689_Y));
KC_AND2_X2 D2688 ( .B(D16589_Y), .A(D16659_Y), .Y(D2688_Y));
KC_AND2_X2 D2263 ( .B(D11418_Y), .A(D11183_Y), .Y(D2263_Y));
KC_AND2_X2 D1946 ( .B(D9721_Y), .A(D9850_Y), .Y(D1946_Y));
KC_AND2_X2 D1800 ( .B(D6567_Y), .A(D11633_Y), .Y(D1800_Y));
KC_AND2_X2 D1799 ( .B(D6567_Y), .A(D11633_Y), .Y(D1799_Y));
KC_AND2_X2 D1795 ( .B(D56_Y), .A(D6149_Y), .Y(D1795_Y));
KC_AND2_X2 D1520 ( .B(D1535_Y), .A(D11633_Y), .Y(D1520_Y));
KC_AND2_X2 D1388 ( .B(D8662_Y), .A(D9850_Y), .Y(D1388_Y));
KC_AND2_X2 D1055 ( .B(D13009_Y), .A(D14315_Y), .Y(D1055_Y));
KC_AND2_X2 D708 ( .B(D5253_Y), .A(D11633_Y), .Y(D708_Y));
KC_XNOR2_X2 D16202 ( .Y(D16202_Y), .A(D16215_Y), .B(D16229_Y));
KC_XNOR2_X2 D16201 ( .Y(D16201_Y), .A(D16219_Y), .B(D16236_Y));
KC_XNOR2_X2 D16200 ( .Y(D16200_Y), .A(D16031_Y), .B(D2588_Y));
KC_XNOR2_X2 D16198 ( .Y(D16198_Y), .A(D16023_Y), .B(D15307_Y));
KC_XNOR2_X2 D16166 ( .Y(D16166_Y), .A(D16027_Y), .B(D15275_Y));
KC_XNOR2_X2 D16139 ( .Y(D16139_Y), .A(D16025_Y), .B(D15287_Y));
KC_XNOR2_X2 D16132 ( .Y(D16132_Y), .A(D16075_Y), .B(D15297_Y));
KC_XNOR2_X2 D16800 ( .Y(D16800_Y), .A(D15252_Y), .B(D15308_Y));
KC_XNOR2_X2 D9553 ( .Y(D9553_Y), .A(D2670_Y), .B(D15296_Y));
KC_XNOR2_X2 D6977 ( .Y(D6977_Y), .A(D16032_Y), .B(D566_Y));
KC_XNOR2_X2 D6976 ( .Y(D6976_Y), .A(D2512_Y), .B(D14640_Y));
KC_XNOR2_X2 D6975 ( .Y(D6975_Y), .A(D15251_Y), .B(D572_Y));
KC_XNOR2_X2 D6111 ( .Y(D6111_Y), .A(D16030_Y), .B(D15285_Y));
KC_XNOR2_X2 D16130 ( .Y(D16130_Y), .A(D9371_Y), .B(D605_Q));
KC_XNOR2_X2 D16129 ( .Y(D16129_Y), .A(D10179_Y), .B(D12236_Q));
KC_XNOR2_X2 D16128 ( .Y(D16128_Y), .A(D2329_Y), .B(D12185_Q));
KC_XNOR2_X2 D16070 ( .Y(D16070_Y), .A(D10797_Y), .B(D10794_Y));
KC_XNOR2_X2 D15460 ( .Y(D15460_Y), .A(D10311_Q), .B(D9406_Y));
KC_XNOR2_X2 D15457 ( .Y(D15457_Y), .A(D10303_Q), .B(D10196_Y));
KC_XNOR2_X2 D15440 ( .Y(D15440_Y), .A(D10701_Y), .B(D11212_Y));
KC_XNOR2_X2 D15439 ( .Y(D15439_Y), .A(D2127_Y), .B(D326_Q));
KC_XNOR2_X2 D16794 ( .Y(D16794_Y), .A(D8864_Y), .B(D8899_Q));
KC_XNOR2_X2 D16793 ( .Y(D16793_Y), .A(D8860_Y), .B(D8898_Q));
KC_XNOR2_X2 D16792 ( .Y(D16792_Y), .A(D8866_Y), .B(D8896_Q));
KC_XNOR2_X2 D16791 ( .Y(D16791_Y), .A(D8919_Y), .B(D8824_Q));
KC_XNOR2_X2 D16790 ( .Y(D16790_Y), .A(D8918_Y), .B(D305_Q));
KC_XNOR2_X2 D2874 ( .Y(D2874_Y), .A(D300_Q), .B(D2710_Y));
KC_XNOR2_X2 D16788 ( .Y(D16788_Y), .A(D2999_Q), .B(D2715_Y));
KC_XNOR2_X2 D16787 ( .Y(D16787_Y), .A(D2883_Q), .B(D2713_Y));
KC_XNOR2_X2 D16786 ( .Y(D16786_Y), .A(D4485_Q), .B(D2714_Y));
KC_XNOR2_X2 D16785 ( .Y(D16785_Y), .A(D3003_Q), .B(D2707_Y));
KC_XNOR2_X2 D16784 ( .Y(D16784_Y), .A(D297_Q), .B(D2709_Y));
KC_XNOR2_X2 D16783 ( .Y(D16783_Y), .A(D3001_Q), .B(D2701_Y));
KC_XNOR2_X2 D16782 ( .Y(D16782_Y), .A(D265_Q), .B(D2706_Y));
KC_XNOR2_X2 D16779 ( .Y(D16779_Y), .A(D298_Q), .B(D2702_Y));
KC_XNOR2_X2 D15246 ( .Y(D15246_Y), .A(D3002_Q), .B(D2703_Y));
KC_XNOR2_X2 D14583 ( .Y(D14583_Y), .A(D3000_Q), .B(D2705_Y));
KC_XNOR2_X2 D14580 ( .Y(D14580_Y), .A(D4486_Q), .B(D2704_Y));
KC_XNOR2_X2 D14578 ( .Y(D14578_Y), .A(D299_Q), .B(D2700_Y));
KC_XNOR2_X2 D15438 ( .Y(D15438_Y), .A(D16081_Y), .B(D15292_Y));
KC_XNOR2_X2 D15437 ( .Y(D15437_Y), .A(D16074_Y), .B(D15286_Y));
KC_XNOR2_X2 D15433 ( .Y(D15433_Y), .A(D15274_Y), .B(D16026_Y));
KC_BUF_X16 D610 ( .Y(D610_Y), .A(D1848_Y));
KC_AOI31_X2 D621 ( .B0(D2312_Y), .B1(D8001_Y), .B2(D7668_Y),     .Y(D621_Y), .A(D8003_Y));
KC_NOR3_X3 D10372 ( .B(D2176_Y), .Y(D10372_Y), .C(D8295_Y),     .A(D10362_Q));
KC_NOR3_X3 D10369 ( .B(D2155_Y), .Y(D10369_Y), .C(D8295_Y),     .A(D10362_Q));
KC_NOR3_X3 D620 ( .B(D10186_Y), .Y(D620_Y), .C(D9364_Y), .A(D8044_Y));
KC_OAI22_X2 D547 ( .A1(D14506_Y), .B0(D14505_Y), .B1(D14567_Y),     .A0(D14643_Y), .Y(D547_Y));
KC_TLATHQ_X3 D12179 ( .D(D14806_Y), .Q(D12179_Q), .GN(D534_Y));
KC_TLATHQ_X3 D11673 ( .D(D12138_Y), .Q(D11673_Q), .GN(D540_Q));
KC_TLATHQ_X3 D11641 ( .D(D7488_Y), .Q(D11641_Q), .GN(D11629_Y));
KC_TLATHQ_X3 D11640 ( .D(D7164_Y), .Q(D11640_Q), .GN(D11621_Y));
KC_TLATHQ_X3 D11639 ( .D(D12136_Y), .Q(D11639_Q), .GN(D11637_Q));
KC_TLATHQ_X3 D11638 ( .D(D11616_Y), .Q(D11638_Q), .GN(D11637_Q));
KC_TLATHQ_X3 D2174 ( .D(D11634_Y), .Q(D2174_Q), .GN(D11636_Q));
KC_TLATHQ_X3 D2104 ( .D(D11634_Y), .Q(D2104_Q), .GN(D11620_Y));
KC_TLATHQ_X3 D540 ( .D(D11614_Y), .Q(D540_Q), .GN(D540_GN));
KC_TLATHQ_X3 D539 ( .D(D11616_Y), .Q(D539_Q), .GN(D11624_Y));
KC_BUF_X10 D15807 ( .Y(D15807_Y), .A(D14228_Y));
KC_BUF_X10 D15219 ( .Y(D15219_Y), .A(D14228_Y));
KC_BUF_X10 D15083 ( .Y(D15083_Y), .A(D14228_Y));
KC_BUF_X10 D10821 ( .Y(D10821_Y), .A(D10705_Y));
KC_BUF_X10 D10633 ( .Y(D10633_Y), .A(D11640_Q));
KC_BUF_X10 D10176 ( .Y(D10176_Y), .A(D10187_Y));
KC_BUF_X10 D6615 ( .Y(D6615_Y), .A(D9359_Y));
KC_BUF_X10 D5812 ( .Y(D5812_Y), .A(D9315_Y));
KC_BUF_X10 D1663 ( .Y(D1663_Y), .A(D6615_Y));
KC_BUF_X10 D833 ( .Y(D833_Y), .A(D1059_Y));
KC_BUF_X10 D536 ( .Y(D536_Y), .A(D6615_Y));
KC_NOR2_X4 D10132 ( .Y(D10132_Y), .B(D10106_Y), .A(D10133_Y));
KC_NOR2_X4 D7609 ( .Y(D7609_Y), .B(D7430_Y), .A(D7470_Y));
KC_NOR2_X4 D7305 ( .Y(D7305_Y), .B(D7273_Y), .A(D7250_Y));
KC_NOR2_X4 D5936 ( .Y(D5936_Y), .B(D5685_Y), .A(D7460_Y));
KC_NOR2_X4 D1953 ( .Y(D1953_Y), .B(D8017_Y), .A(D2343_Y));
KC_NOR2_X4 D535 ( .Y(D535_Y), .B(D9343_Y), .A(D9349_Y));
KC_BUF_X11 D16476 ( .Y(D16476_Y), .A(D15988_QN));
KC_BUF_X11 D14315 ( .Y(D14315_Y), .A(D11630_Y));
KC_BUF_X11 D13910 ( .Y(D13910_Y), .A(D13249_Y));
KC_BUF_X11 D13404 ( .Y(D13404_Y), .A(D13249_Y));
KC_BUF_X11 D13283 ( .Y(D13283_Y), .A(D13214_QN));
KC_BUF_X11 D13206 ( .Y(D13206_Y), .A(D13214_QN));
KC_BUF_X11 D12859 ( .Y(D12859_Y), .A(D13249_Y));
KC_BUF_X11 D12750 ( .Y(D12750_Y), .A(D833_Y));
KC_BUF_X11 D12104 ( .Y(D12104_Y), .A(D11567_Y));
KC_BUF_X11 D11183 ( .Y(D11183_Y), .A(D11630_Y));
KC_BUF_X11 D9947 ( .Y(D9947_Y), .A(D9947_A));
KC_BUF_X11 D9850 ( .Y(D9850_Y), .A(D11630_Y));
KC_BUF_X11 D9224 ( .Y(D9224_Y), .A(D9208_Y));
KC_BUF_X11 D6484 ( .Y(D6484_Y), .A(D6461_Y));
KC_BUF_X11 D4827 ( .Y(D4827_Y), .A(D965_Y));
KC_BUF_X11 D2522 ( .Y(D2522_Y), .A(D12743_Y));
KC_BUF_X11 D2356 ( .Y(D2356_Y), .A(D12179_Q));
KC_BUF_X11 D534 ( .Y(D534_Y), .A(D10187_Y));
KC_AO222_X1 D8828 ( .A1(D8753_Y), .B0(D8757_Y), .B1(D8757_Y),     .C0(D8793_Y), .C1(D8773_Y), .Y(D8828_Y), .A0(D8782_Y));
KC_AO222_X1 D7977 ( .A1(D6547_Q), .B0(D7932_Y), .B1(D8272_Y),     .C0(D8399_Y), .C1(D7919_Y), .Y(D7977_Y), .A0(D7920_Y));
KC_AO222_X1 D7976 ( .A1(D517_Q), .B0(D7932_Y), .B1(D8270_Y),     .C0(D8409_Y), .C1(D7919_Y), .Y(D7976_Y), .A0(D7920_Y));
KC_AO222_X1 D7814 ( .A1(D4811_Y), .B0(D725_Y), .B1(D7767_Y),     .C0(D7771_Y), .C1(D8065_Y), .Y(D7814_Y), .A0(D6383_Q));
KC_AO222_X1 D7813 ( .A1(D4811_Y), .B0(D13171_Y), .B1(D7767_Y),     .C0(D7771_Y), .C1(D7958_Y), .Y(D7813_Y), .A0(D1792_Q));
KC_AO222_X1 D7812 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D6385_Q),     .C0(D8072_Y), .C1(D7771_Y), .Y(D7812_Y), .A0(D12764_Y));
KC_AO222_X1 D7811 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D7793_Q),     .C0(D8061_Y), .C1(D7771_Y), .Y(D7811_Y), .A0(D13287_Y));
KC_AO222_X1 D7810 ( .A1(D4811_Y), .B0(D12863_Y), .B1(D7767_Y),     .C0(D7771_Y), .C1(D7957_Y), .Y(D7810_Y), .A0(D452_Q));
KC_AO222_X1 D7809 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D6382_Q),     .C0(D8070_Y), .C1(D7771_Y), .Y(D7809_Y), .A0(D13288_Y));
KC_AO222_X1 D7807 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D450_Q),     .C0(D8068_Y), .C1(D7771_Y), .Y(D7807_Y), .A0(D12300_Y));
KC_AO222_X1 D7806 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D7789_Q),     .C0(D8071_Y), .C1(D7771_Y), .Y(D7806_Y), .A0(D724_Y));
KC_AO222_X1 D7805 ( .A1(D4811_Y), .B0(D12762_Y), .B1(D7767_Y),     .C0(D7771_Y), .C1(D8063_Y), .Y(D7805_Y), .A0(D7794_Q));
KC_AO222_X1 D7804 ( .A1(D7763_Y), .B0(D9254_Y), .B1(D7763_Y),     .C0(D7821_Y), .C1(D447_Y), .Y(D7804_Y), .A0(D7762_Y));
KC_AO222_X1 D7802 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D7790_Q),     .C0(D8067_Y), .C1(D7771_Y), .Y(D7802_Y), .A0(D12763_Y));
KC_AO222_X1 D7801 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D7791_Q),     .C0(D8066_Y), .C1(D7771_Y), .Y(D7801_Y), .A0(D12761_Y));
KC_AO222_X1 D7798 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D6387_Q),     .C0(D8069_Y), .C1(D7771_Y), .Y(D7798_Y), .A0(D723_Q));
KC_AO222_X1 D7298 ( .A1(D7249_Y), .B0(D5804_Y), .B1(D7213_Y),     .C0(D7140_Y), .C1(D7098_Y), .Y(D7298_Y), .A0(D7302_Y));
KC_AO222_X1 D6485 ( .A1(D1695_Y), .B0(D6465_Y), .B1(D4961_Y),     .C0(D1746_Y), .C1(D1745_Y), .Y(D6485_Y), .A0(D1817_Y));
KC_AO222_X1 D6196 ( .A1(D6205_Y), .B0(D6166_Y), .B1(D6172_Y),     .C0(D6166_Y), .C1(D6209_Y), .Y(D6196_Y), .A0(D6160_Y));
KC_AO222_X1 D6127 ( .A1(D4307_Y), .B0(D4392_Y), .B1(D2893_Y),     .C0(D4388_Y), .C1(D4385_Y), .Y(D6127_Y), .A0(D4308_Y));
KC_AO222_X1 D5937 ( .A1(D4721_Y), .B0(D259_Y), .B1(D5934_Y),     .C0(D7392_Y), .C1(D7367_Y), .Y(D5937_Y), .A0(D5932_Y));
KC_AO222_X1 D4828 ( .A1(D4772_Y), .B0(D4776_Y), .B1(D4662_Y),     .C0(D4771_Y), .C1(D4834_Y), .Y(D4828_Y), .A0(D1456_Y));
KC_AO222_X1 D4559 ( .A1(D4513_Y), .B0(D29_Y), .B1(D4411_Y),     .C0(D1593_Y), .C1(D4466_Y), .Y(D4559_Y), .A0(D4466_Y));
KC_AO222_X1 D4492 ( .A1(D4407_Y), .B0(D4389_Y), .B1(D4404_Y),     .C0(D4546_Y), .C1(D10045_Y), .Y(D4492_Y), .A0(D4450_Y));
KC_AO222_X1 D4236 ( .A1(D5863_Y), .B0(D4233_Y), .B1(D4264_Y),     .C0(D228_Q), .C1(D4196_Y), .Y(D4236_Y), .A0(D4220_Y));
KC_AO222_X1 D4128 ( .A1(D4106_Y), .B0(D1595_Y), .B1(D1538_Y),     .C0(D4124_Y), .C1(D2716_Y), .Y(D4128_Y), .A0(D1595_Y));
KC_AO222_X1 D3090 ( .A1(D3050_Y), .B0(D3035_Y), .B1(D3010_Y),     .C0(D3035_Y), .C1(D6255_Y), .Y(D3090_Y), .A0(D3010_Y));
KC_AO222_X1 D1959 ( .A1(D7767_Y), .B0(D4811_Y), .B1(D1791_Q),     .C0(D8064_Y), .C1(D7771_Y), .Y(D1959_Y), .A0(D13280_Q));
KC_AO222_X1 D1958 ( .A1(D4811_Y), .B0(D13289_Y), .B1(D7767_Y),     .C0(D7771_Y), .C1(D7959_Y), .Y(D1958_Y), .A0(D6386_Q));
KC_AO222_X1 D537 ( .A1(D521_Q), .B0(D7932_Y), .B1(D8277_Y),     .C0(D8417_Y), .C1(D7919_Y), .Y(D537_Y), .A0(D7920_Y));
KC_AO222_X1 D457 ( .A1(D4811_Y), .B0(D13285_Y), .B1(D7767_Y),     .C0(D7771_Y), .C1(D615_Y), .Y(D457_Y), .A0(D6384_Q));
KC_NAND4B_X1 D16551 ( .B(D1381_Q), .C(D16538_Y), .Y(D16551_Y),     .DN(D16535_Y), .A(D16556_Q));
KC_NAND4B_X1 D16550 ( .B(D16534_Y), .C(D16536_Y), .Y(D16550_Y),     .DN(D16542_Y), .A(D1381_Q));
KC_NAND4B_X1 D16458 ( .B(D16473_Q), .C(D16434_Y), .Y(D16458_Y),     .DN(D16448_Y), .A(D1322_Q));
KC_NAND4B_X1 D16457 ( .B(D1322_Q), .C(D16439_Y), .Y(D16457_Y),     .DN(D16417_Y), .A(D16471_Q));
KC_NAND4B_X1 D16286 ( .B(D16289_Q), .C(D16256_Y), .Y(D16286_Y),     .DN(D16290_Q), .A(D16293_Q));
KC_NAND4B_X1 D16224 ( .B(D15508_Y), .C(D16191_Y), .Y(D16224_Y),     .DN(D16379_Y), .A(D16382_Y));
KC_NAND4B_X1 D15567 ( .B(D15533_Y), .C(D15515_Y), .Y(D15567_Y),     .DN(D15582_Y), .A(D15530_Y));
KC_NAND4B_X1 D15258 ( .B(D14586_Y), .C(D15243_Y), .Y(D15258_Y),     .DN(D15306_Y), .A(D327_Y));
KC_NAND4B_X1 D14683 ( .B(D14634_Y), .C(D14630_Y), .Y(D14683_Y),     .DN(D14621_Y), .A(D14685_Q));
KC_NAND4B_X1 D12988 ( .B(D12933_Y), .C(D13001_Y), .Y(D12988_Y),     .DN(D12949_Y), .A(D12942_Y));
KC_NAND4B_X1 D12847 ( .B(D12813_Y), .C(D12703_Y), .Y(D12847_Y),     .DN(D13268_Q), .A(D12756_Q));
KC_NAND4B_X1 D12273 ( .B(D11660_Y), .C(D12268_Y), .Y(D12273_Y),     .DN(D12190_Y), .A(D11655_Y));
KC_NAND4B_X1 D10186 ( .B(D392_Y), .C(D6285_Y), .Y(D10186_Y),     .DN(D16_Y), .A(D11655_Y));
KC_NAND4B_X1 D9382 ( .B(D10179_Y), .C(D9387_Y), .Y(D9382_Y),     .DN(D4619_Y), .A(D12187_Y));
KC_NAND4B_X1 D9270 ( .B(D9247_Y), .C(D9300_Y), .Y(D9270_Y),     .DN(D9282_Y), .A(D9300_Y));
KC_NAND4B_X1 D8819 ( .B(D8775_Y), .C(D8755_Y), .Y(D8819_Y),     .DN(D8774_Y), .A(D8774_Y));
KC_NAND4B_X1 D8338 ( .B(D8281_Y), .C(D957_Y), .Y(D8338_Y),     .DN(D8281_Y), .A(D8282_Y));
KC_NAND4B_X1 D8242 ( .B(D8246_Q), .C(D8201_Y), .Y(D8242_Y),     .DN(D8247_Q), .A(D8249_Q));
KC_NAND4B_X1 D7972 ( .B(D7985_Y), .C(D7961_Y), .Y(D7972_Y),     .DN(D7928_Y), .A(D7934_Y));
KC_NAND4B_X1 D7891 ( .B(D7838_Y), .C(D6429_Y), .Y(D7891_Y),     .DN(D1857_Y), .A(D7832_Y));
KC_NAND4B_X1 D7787 ( .B(D9320_Y), .C(D7776_Y), .Y(D7787_Y),     .DN(D10154_Y), .A(D10155_Y));
KC_NAND4B_X1 D7474 ( .B(D8991_Y), .C(D7465_Y), .Y(D7474_Y),     .DN(D6048_Y), .A(D8938_Y));
KC_NAND4B_X1 D7389 ( .B(D5825_Y), .C(D7396_Y), .Y(D7389_Y),     .DN(D5837_Y), .A(D7336_Y));
KC_NAND4B_X1 D7296 ( .B(D186_Y), .C(D7260_Y), .Y(D7296_Y),     .DN(D7097_Y), .A(D7140_Y));
KC_NAND4B_X1 D7143 ( .B(D7109_Y), .C(D7124_Y), .Y(D7143_Y),     .DN(D5880_Y), .A(D192_Q));
KC_NAND4B_X1 D6479 ( .B(D5030_Y), .C(D6443_Y), .Y(D6479_Y),     .DN(D6445_Y), .A(D5039_Y));
KC_NAND4B_X1 D6265 ( .B(D6268_Y), .C(D6274_Y), .Y(D6265_Y),     .DN(D6240_Y), .A(D6236_Y));
KC_NAND4B_X1 D5933 ( .B(D7335_Y), .C(D7330_Y), .Y(D5933_Y),     .DN(D5932_Y), .A(D7335_Y));
KC_NAND4B_X1 D5685 ( .B(D5669_Y), .C(D5665_Y), .Y(D5685_Y),     .DN(D5675_Y), .A(D5689_Q));
KC_NAND4B_X1 D5080 ( .B(D4983_Y), .C(D5054_Y), .Y(D5080_Y),     .DN(D5055_Y), .A(D5084_Y));
KC_NAND4B_X1 D4964 ( .B(D445_Q), .C(D446_Q), .Y(D4964_Y), .DN(D6363_Y),     .A(D444_Q));
KC_NAND4B_X1 D4963 ( .B(D5085_Y), .C(D4879_Y), .Y(D4963_Y),     .DN(D3410_Y), .A(D3534_Y));
KC_NAND4B_X1 D4816 ( .B(D4779_Y), .C(D6329_Y), .Y(D4816_Y),     .DN(D4835_Y), .A(D4785_Y));
KC_NAND4B_X1 D4815 ( .B(D4836_Y), .C(D4781_Y), .Y(D4815_Y),     .DN(D1655_Q), .A(D4756_Y));
KC_NAND4B_X1 D4726 ( .B(D3274_Y), .C(D4718_S), .Y(D4726_Y),     .DN(D3274_Y), .A(D3274_Y));
KC_NAND4B_X1 D4635 ( .B(D344_Y), .C(D4612_Y), .Y(D4635_Y),     .DN(D4596_Y), .A(D72_Y));
KC_NAND4B_X1 D4552 ( .B(D4500_Y), .C(D4504_Y), .Y(D4552_Y),     .DN(D3040_Y), .A(D1431_Y));
KC_NAND4B_X1 D4392 ( .B(D2956_Y), .C(D4115_Y), .Y(D4392_Y),     .DN(D4310_Y), .A(D2881_Y));
KC_NAND4B_X1 D4234 ( .B(D5726_Y), .C(D4120_Q), .Y(D4234_Y),     .DN(D4197_Y), .A(D4204_Y));
KC_NAND4B_X1 D3480 ( .B(D3305_Y), .C(D3306_Y), .Y(D3480_Y),     .DN(D3427_Y), .A(D3371_Y));
KC_NAND4B_X1 D3381 ( .B(D3380_Y), .C(D3331_Y), .Y(D3381_Y),     .DN(D3284_Y), .A(D3321_Y));
KC_NAND4B_X1 D3380 ( .B(D3323_Y), .C(D3208_Y), .Y(D3380_Y),     .DN(D3206_Y), .A(D3369_Y));
KC_NAND4B_X1 D3378 ( .B(D3372_Q), .C(D3303_Y), .Y(D3378_Y),     .DN(D3304_Y), .A(D3376_Q));
KC_NAND4B_X1 D3278 ( .B(D3222_Y), .C(D1428_Y), .Y(D3278_Y),     .DN(D1574_Y), .A(D3264_Y));
KC_NAND4B_X1 D3277 ( .B(D1427_Y), .C(D3225_Y), .Y(D3277_Y),     .DN(D396_Y), .A(D3348_Y));
KC_NAND4B_X1 D3183 ( .B(D3185_Q), .C(D1430_Y), .Y(D3183_Y),     .DN(D3132_Y), .A(D3188_Q));
KC_NAND4B_X1 D3074 ( .B(D3029_Y), .C(D4506_Y), .Y(D3074_Y),     .DN(D3029_Y), .A(D3029_Y));
KC_NAND4B_X1 D2881 ( .B(D2831_Y), .C(D4310_Y), .Y(D2881_Y),     .DN(D4115_Y), .A(D2831_Y));
KC_NAND4B_X1 D2793 ( .B(D2766_Y), .C(D2737_Y), .Y(D2793_Y),     .DN(D2746_Y), .A(D2755_Y));
KC_NAND4B_X1 D812 ( .B(D12814_Y), .C(D12813_Y), .Y(D812_Y),     .DN(D13268_Q), .A(D12756_Q));
KC_NAND4B_X1 D528 ( .B(D15259_Y), .C(D705_Y), .Y(D528_Y),     .DN(D16077_Y), .A(D15248_S));
KC_NAND4B_X1 D448 ( .B(D454_Y), .C(D6370_Y), .Y(D448_Y), .DN(D4917_Y),     .A(D4940_Y));
KC_OR3_X1 D16549 ( .Y(D16549_Y), .C(D16544_Y), .B(D16487_Y),     .A(D16556_Q));
KC_OR3_X1 D14233 ( .Y(D14233_Y), .C(D14236_Q), .B(D14265_Q),     .A(D14245_Q));
KC_OR3_X1 D10106 ( .Y(D10106_Y), .C(D10067_Y), .B(D10085_Y),     .A(D10086_Y));
KC_OR3_X1 D9350 ( .Y(D9350_Y), .C(D9343_Y), .B(D9357_Y), .A(D9344_Y));
KC_OR3_X1 D9003 ( .Y(D9003_Y), .C(D9216_Q), .B(D7739_Y), .A(D9159_Q));
KC_OR3_X1 D8807 ( .Y(D8807_Y), .C(D8705_Y), .B(D8817_Y), .A(D8786_Y));
KC_OR3_X1 D6464 ( .Y(D6464_Y), .C(D468_Y), .B(D5017_Y), .A(D4989_Y));
KC_OR3_X1 D4956 ( .Y(D4956_Y), .C(D4960_Y), .B(D3371_Y), .A(D7968_Q));
KC_OR3_X1 D2633 ( .Y(D2633_Y), .C(D16392_Q), .B(D16389_Q),     .A(D16391_Q));
KC_OR3_X1 D441 ( .Y(D441_Y), .C(D6375_Q), .B(D6376_Q), .A(D444_Q));
KC_OAI22_X3 D431 ( .A1(D9113_Y), .B0(D1904_Y), .B1(D5963_Y),     .A0(D7684_Y), .Y(D431_Y));
KC_OA21_X1 D16687 ( .A0(D16682_Q), .B(D16690_Y), .A1(D16689_Y),     .Y(D16687_Y));
KC_OA21_X1 D16686 ( .A0(D16684_Q), .B(D16688_Y), .A1(D16695_Y),     .Y(D16686_Y));
KC_OA21_X1 D16685 ( .A0(D16681_Q), .B(D16692_Y), .A1(D16691_Y),     .Y(D16685_Y));
KC_OA21_X1 D16664 ( .A0(D16650_Q), .B(D16670_Y), .A1(D16643_Y),     .Y(D16664_Y));
KC_OA21_X1 D16663 ( .A0(D16660_Q), .B(D16666_Y), .A1(D16669_Y),     .Y(D16663_Y));
KC_OA21_X1 D16662 ( .A0(D1373_Q), .B(D16668_Y), .A1(D16646_Y),     .Y(D16662_Y));
KC_OA21_X1 D16638 ( .A0(D1396_Q), .B(D16642_Y), .A1(D16640_Y),     .Y(D16638_Y));
KC_OA21_X1 D16170 ( .A0(D16148_Y), .B(D16187_Y), .A1(D16095_Y),     .Y(D16170_Y));
KC_OA21_X1 D16085 ( .A0(D16051_Y), .B(D16100_Y), .A1(D16120_Y),     .Y(D16085_Y));
KC_OA21_X1 D15239 ( .A0(D15228_Y), .B(D15240_Y), .A1(D15183_Y),     .Y(D15239_Y));
KC_OA21_X1 D14592 ( .A0(D14519_Q), .B(D16770_Y), .A1(D14609_Y),     .Y(D14592_Y));
KC_OA21_X1 D14590 ( .A0(D14601_Q), .B(D14602_Y), .A1(D16769_Y),     .Y(D14590_Y));
KC_OA21_X1 D14589 ( .A0(D14518_Q), .B(D14608_Y), .A1(D14607_Y),     .Y(D14589_Y));
KC_OA21_X1 D14588 ( .A0(D2512_Y), .B(D14606_Y), .A1(D14605_Y),     .Y(D14588_Y));
KC_OA21_X1 D14587 ( .A0(D14688_Q), .B(D14604_Y), .A1(D14687_Q),     .Y(D14587_Y));
KC_OA21_X1 D13912 ( .A0(D14520_Q), .B(D13922_Y), .A1(D13925_Y),     .Y(D13912_Y));
KC_OA21_X1 D13911 ( .A0(D608_Q), .B(D13924_Y), .A1(D14603_Y),     .Y(D13911_Y));
KC_OA21_X1 D13863 ( .A0(D13865_Q), .B(D13873_Y), .A1(D13872_Q),     .Y(D13863_Y));
KC_OA21_X1 D13862 ( .A0(D543_Q), .B(D13868_Y), .A1(D13870_Y),     .Y(D13862_Y));
KC_OA21_X1 D13861 ( .A0(D13864_Q), .B(D13871_Y), .A1(D13874_Y),     .Y(D13861_Y));
KC_OA21_X1 D13174 ( .A0(D13175_Q), .B(D16763_Y), .A1(D13869_Y),     .Y(D13174_Y));
KC_OA21_X1 D9282 ( .A0(D9246_Y), .B(D9299_Y), .A1(D9247_Y),     .Y(D9282_Y));
KC_OA21_X1 D8352 ( .A0(D8294_Y), .B(D8357_Y), .A1(D6773_Y),     .Y(D8352_Y));
KC_OA21_X1 D8256 ( .A0(D8239_Y), .B(D8262_Y), .A1(D8219_Y),     .Y(D8256_Y));
KC_OA21_X1 D7740 ( .A0(D7706_Y), .B(D7753_Y), .A1(D9210_Y),     .Y(D7740_Y));
KC_OA21_X1 D6276 ( .A0(D6254_Y), .B(D14139_Y), .A1(D6238_Y),     .Y(D6276_Y));
KC_OA21_X1 D6274 ( .A0(D6212_Y), .B(D12130_Y), .A1(D6240_Y),     .Y(D6274_Y));
KC_OA21_X1 D6198 ( .A0(D6157_Y), .B(D9105_Y), .A1(D6183_Y),     .Y(D6198_Y));
KC_OA21_X1 D6129 ( .A0(D16143_Y), .B(D6368_Y), .A1(D6105_Y),     .Y(D6129_Y));
KC_OA21_X1 D5083 ( .A0(D5064_Y), .B(D5097_Y), .A1(D3633_Y),     .Y(D5083_Y));
KC_OA21_X1 D4835 ( .A0(D4700_Y), .B(D4843_Y), .A1(D4779_Y),     .Y(D4835_Y));
KC_OA21_X1 D4834 ( .A0(D3385_Q), .B(D3391_Y), .A1(D4846_Y),     .Y(D4834_Y));
KC_OA21_X1 D4833 ( .A0(D4817_Q), .B(D4850_Y), .A1(D4853_Y),     .Y(D4833_Y));
KC_OA21_X1 D4832 ( .A0(D1655_Q), .B(D4851_Y), .A1(D4849_Y),     .Y(D4832_Y));
KC_OA21_X1 D4831 ( .A0(D4825_Q), .B(D4854_Y), .A1(D4848_Y),     .Y(D4831_Y));
KC_OA21_X1 D4830 ( .A0(D4824_Q), .B(D4858_Y), .A1(D4856_Y),     .Y(D4830_Y));
KC_OA21_X1 D4829 ( .A0(D4823_Q), .B(D4855_Y), .A1(D4852_Y),     .Y(D4829_Y));
KC_OA21_X1 D4245 ( .A0(D232_Q), .B(D4251_Y), .A1(D4258_Y),     .Y(D4245_Y));
KC_OA21_X1 D4244 ( .A0(D4136_Q), .B(D4254_Y), .A1(D5693_Q),     .Y(D4244_Y));
KC_OA21_X1 D4243 ( .A0(D165_Y), .B(D4255_Y), .A1(D4261_Y),     .Y(D4243_Y));
KC_OA21_X1 D4242 ( .A0(D228_Q), .B(D4260_Y), .A1(D2810_Y),     .Y(D4242_Y));
KC_OA21_X1 D4241 ( .A0(D229_Q), .B(D4259_Y), .A1(D4253_Y),     .Y(D4241_Y));
KC_OA21_X1 D4240 ( .A0(D4150_Y), .B(D4265_Y), .A1(D235_Y),     .Y(D4240_Y));
KC_OA21_X1 D4239 ( .A0(D8838_Y), .B(D4268_Y), .A1(D4266_Y),     .Y(D4239_Y));
KC_OA21_X1 D4238 ( .A0(D4235_Q), .B(D237_Y), .A1(D2815_Y),     .Y(D4238_Y));
KC_OA21_X1 D4237 ( .A0(D239_Q), .B(D238_Y), .A1(D4267_Y), .Y(D4237_Y));
KC_OA21_X1 D4133 ( .A0(D4121_Q), .B(D4147_Y), .A1(D4252_Y),     .Y(D4133_Y));
KC_OA21_X1 D4132 ( .A0(D4149_Q), .B(D4152_Y), .A1(D4256_Y),     .Y(D4132_Y));
KC_OA21_X1 D4131 ( .A0(D4122_Q), .B(D4142_Y), .A1(D4139_Y),     .Y(D4131_Y));
KC_OA21_X1 D4130 ( .A0(D4120_Q), .B(D4143_Y), .A1(D4141_Y),     .Y(D4130_Y));
KC_OA21_X1 D4129 ( .A0(D4119_Q), .B(D4140_Y), .A1(D4148_Y),     .Y(D4129_Y));
KC_OA21_X1 D3288 ( .A0(D3265_Y), .B(D3295_Y), .A1(D3266_Y),     .Y(D3288_Y));
KC_OA21_X1 D2895 ( .A0(D2885_Q), .B(D2900_Y), .A1(D2788_Y),     .Y(D2895_Y));
KC_OA21_X1 D2690 ( .A0(D16599_Q), .B(D2691_Y), .A1(D16665_Y),     .Y(D2690_Y));
KC_OA21_X1 D2102 ( .A0(D9672_Y), .B(D2109_Y), .A1(D2061_Y),     .Y(D2102_Y));
KC_OA21_X1 D1399 ( .A0(D1395_Q), .B(D16694_Y), .A1(D16671_Y),     .Y(D1399_Y));
KC_OA21_X1 D1398 ( .A0(D1400_Q), .B(D1406_Y), .A1(D1320_Q),     .Y(D1398_Y));
KC_OA21_X1 D426 ( .A0(D3383_Q), .B(D4845_Y), .A1(D4819_Q), .Y(D426_Y));
KC_OA21_X1 D425 ( .A0(D4826_Q), .B(D4847_Y), .A1(D3993_Y), .Y(D425_Y));
KC_DFFSNHQ_X1 D12143 ( .Q(D12143_Q), .D(D12146_Y), .SN(D11636_SN),     .CK(D709_Y));
KC_DFFSNHQ_X1 D9353 ( .Q(D9353_Q), .D(D9317_Y), .SN(D7893_Y),     .CK(D10107_QN));
KC_DFFSNHQ_X1 D9324 ( .Q(D9324_Q), .D(D9311_Y), .SN(D7892_Y),     .CK(D9212_QN));
KC_DFFSNHQ_X1 D9323 ( .Q(D9323_Q), .D(D9311_Y), .SN(D7892_Y),     .CK(D10107_QN));
KC_DFFSNHQ_X1 D9322 ( .Q(D9322_Q), .D(D9316_Y), .SN(D7892_Y),     .CK(D10107_QN));
KC_DFFSNHQ_X1 D9319 ( .Q(D9319_Q), .D(D9310_Y), .SN(D7892_Y),     .CK(D9212_QN));
KC_DFFSNHQ_X1 D9318 ( .Q(D9318_Q), .D(D9310_Y), .SN(D7892_Y),     .CK(D10107_QN));
KC_DFFSNHQ_X1 D9260 ( .Q(D9260_Q), .D(D9294_Y), .SN(D7892_Y),     .CK(D9212_QN));
KC_DFFSNHQ_X1 D9209 ( .Q(D9209_Q), .D(D9199_Y), .SN(D9214_Y),     .CK(D9212_QN));
KC_DFFSNHQ_X1 D442 ( .Q(D442_Q), .D(D9295_Y), .SN(D9271_Y),     .CK(D10107_QN));
KC_DFFSNHQ_X1 D414 ( .Q(D414_Q), .D(D9176_Y), .SN(D9271_Y),     .CK(D10107_QN));
KC_NAND3_X2 D16524 ( .Y(D16524_Y), .C(D16537_Y), .B(D16536_Y),     .A(D16493_Y));
KC_NAND3_X2 D14805 ( .Y(D14805_Y), .C(D14754_Y), .B(D14807_Y),     .A(D14057_Y));
KC_NAND3_X2 D13409 ( .Y(D13409_Y), .C(D812_Y), .B(D13334_Y),     .A(D14017_Y));
KC_NAND3_X2 D7407 ( .Y(D7407_Y), .C(D8841_Y), .B(D7225_Y),     .A(D5804_Y));
KC_NAND3_X2 D5825 ( .Y(D5825_Y), .C(D5712_Y), .B(D7184_Y),     .A(D1956_Y));
KC_NAND3_X2 D5704 ( .Y(D5704_Y), .C(D5678_Y), .B(D5691_Q),     .A(D5687_Q));
KC_NAND3_X2 D396 ( .Y(D396_Y), .C(D3218_Y), .B(D3234_Y), .A(D3243_Y));
KC_BUF_X14 D9954 ( .Y(D9954_Y), .A(D9970_Y));
KC_BUF_X14 D394 ( .Y(D394_Y), .A(D9149_Q));
KC_MXI2_X3 D10192 ( .Y(D10192_Y), .A(D40_Q), .B(D1702_Y),     .S0(D6342_Y));
KC_MXI2_X3 D10191 ( .Y(D10191_Y), .A(D6248_Q), .B(D6309_Y),     .S0(D6342_Y));
KC_MXI2_X3 D7670 ( .Y(D7670_Y), .A(D4150_Y), .B(D4676_Y),     .S0(D6239_Y));
KC_MXI2_X3 D7669 ( .Y(D7669_Y), .A(D8838_Y), .B(D4677_Y),     .S0(D6239_Y));
KC_MXI2_X3 D7668 ( .Y(D7668_Y), .A(D235_Y), .B(D4675_Y), .S0(D6239_Y));
KC_MXI2_X3 D6410 ( .Y(D6410_Y), .A(D41_Y), .B(D6353_Y), .S0(D6342_Y));
KC_MXI2_X3 D6407 ( .Y(D6407_Y), .A(D7509_Y), .B(D456_Y), .S0(D6342_Y));
KC_MXI2_X3 D6406 ( .Y(D6406_Y), .A(D7613_Y), .B(D6310_Y),     .S0(D6342_Y));
KC_MXI2_X3 D6405 ( .Y(D6405_Y), .A(D334_Q), .B(D455_Y), .S0(D6342_Y));
KC_MXI2_X3 D6281 ( .Y(D6281_Y), .A(D228_Q), .B(D381_Y), .S0(D6239_Y));
KC_MXI2_X3 D1964 ( .Y(D1964_Y), .A(D9099_Y), .B(D7800_Y),     .S0(D6342_Y));
KC_MXI2_X3 D1814 ( .Y(D1814_Y), .A(D51_Y), .B(D4784_Y), .S0(D6342_Y));
KC_MXI2_X3 D1813 ( .Y(D1813_Y), .A(D57_Y), .B(D4841_Y), .S0(D6342_Y));
KC_MXI2_X3 D464 ( .Y(D464_Y), .A(D7502_Y), .B(D7808_Y), .S0(D6342_Y));
KC_MXI2_X3 D463 ( .Y(D463_Y), .A(D36_Y), .B(D7799_Y), .S0(D6342_Y));
KC_MXI2_X3 D462 ( .Y(D462_Y), .A(D9023_Q), .B(D7803_Y), .S0(D6342_Y));
KC_MXI2_X3 D392 ( .Y(D392_Y), .A(D165_Y), .B(D371_Y), .S0(D6239_Y));
KC_OAI21B_X1 D16171 ( .A1(D16079_Y), .B(D16185_Y), .A0N(D16123_Y),     .Y(D16171_Y));
KC_OAI21B_X1 D16086 ( .A1(D16067_Y), .B(D16055_Y), .A0N(D567_Y),     .Y(D16086_Y));
KC_OAI21B_X1 D16001 ( .A1(D14785_Y), .B(D13966_Y), .A0N(D16524_Y),     .Y(D16001_Y));
KC_OAI21B_X1 D15456 ( .A1(D646_Y), .B(D15429_Y), .A0N(D15379_Y),     .Y(D15456_Y));
KC_OAI21B_X1 D13768 ( .A1(D13763_Y), .B(D13752_Y), .A0N(D13747_Y),     .Y(D13768_Y));
KC_OAI21B_X1 D13516 ( .A1(D852_Q), .B(D866_Y), .A0N(D13512_Y),     .Y(D13516_Y));
KC_OAI21B_X1 D12999 ( .A1(D13497_Y), .B(D12995_Q), .A0N(D13590_Y),     .Y(D12999_Y));
KC_OAI21B_X1 D12927 ( .A1(D855_Q), .B(D12872_Y), .A0N(D13697_Y),     .Y(D12927_Y));
KC_OAI21B_X1 D10517 ( .A1(D9746_Y), .B(D10488_Y), .A0N(D10926_Y),     .Y(D10517_Y));
KC_OAI21B_X1 D9585 ( .A1(D622_Y), .B(D9389_Y), .A0N(D9519_Y),     .Y(D9585_Y));
KC_OAI21B_X1 D9584 ( .A1(D9554_Y), .B(D9494_Y), .A0N(D9494_Y),     .Y(D9584_Y));
KC_OAI21B_X1 D9285 ( .A1(D9282_Y), .B(D9270_Y), .A0N(D7547_Y),     .Y(D9285_Y));
KC_OAI21B_X1 D8830 ( .A1(D8827_Y), .B(D2029_Y), .A0N(D8827_Y),     .Y(D8830_Y));
KC_OAI21B_X1 D8829 ( .A1(D8826_Y), .B(D8819_Y), .A0N(D8796_Y),     .Y(D8829_Y));
KC_OAI21B_X1 D8724 ( .A1(D9949_Y), .B(D7781_Y), .A0N(D8681_Y),     .Y(D8724_Y));
KC_OAI21B_X1 D8723 ( .A1(D7142_Y), .B(D8690_Y), .A0N(D190_Y),     .Y(D8723_Y));
KC_OAI21B_X1 D8473 ( .A1(D1835_Y), .B(D8029_Y), .A0N(D8418_Y),     .Y(D8473_Y));
KC_OAI21B_X1 D8472 ( .A1(D1835_Y), .B(D8029_Y), .A0N(D8286_Y),     .Y(D8472_Y));
KC_OAI21B_X1 D8471 ( .A1(D1835_Y), .B(D8029_Y), .A0N(D8410_Y),     .Y(D8471_Y));
KC_OAI21B_X1 D7980 ( .A1(D7950_Y), .B(D7979_Y), .A0N(D6518_Y),     .Y(D7980_Y));
KC_OAI21B_X1 D7979 ( .A1(D1937_Y), .B(D8057_Y), .A0N(D3647_Q),     .Y(D7979_Y));
KC_OAI21B_X1 D7898 ( .A1(D7855_Y), .B(D7859_Y), .A0N(D7890_Q),     .Y(D7898_Y));
KC_OAI21B_X1 D7537 ( .A1(D7571_Y), .B(D37_Y), .A0N(D7514_Y),     .Y(D7537_Y));
KC_OAI21B_X1 D7483 ( .A1(D7446_Y), .B(D7428_Y), .A0N(D7471_Y),     .Y(D7483_Y));
KC_OAI21B_X1 D6279 ( .A1(D6227_Y), .B(D6282_Y), .A0N(D6231_Y),     .Y(D6279_Y));
KC_OAI21B_X1 D6278 ( .A1(D6220_Y), .B(D6337_Y), .A0N(D16147_Y),     .Y(D6278_Y));
KC_OAI21B_X1 D6199 ( .A1(D6166_Y), .B(D56_Y), .A0N(D6160_Y),     .Y(D6199_Y));
KC_OAI21B_X1 D6080 ( .A1(D6011_Y), .B(D5993_Y), .A0N(D284_Y),     .Y(D6080_Y));
KC_OAI21B_X1 D5818 ( .A1(D5901_Y), .B(D4188_Y), .A0N(D5782_Y),     .Y(D5818_Y));
KC_OAI21B_X1 D4966 ( .A1(D4954_Y), .B(D4955_Y), .A0N(D4921_Y),     .Y(D4966_Y));
KC_OAI21B_X1 D4564 ( .A1(D6031_Y), .B(D7337_Y), .A0N(D4563_Q),     .Y(D4564_Y));
KC_OAI21B_X1 D4396 ( .A1(D5863_Y), .B(D4327_Y), .A0N(D4280_Y),     .Y(D4396_Y));
KC_OAI21B_X1 D3583 ( .A1(D4895_Y), .B(D3585_Y), .A0N(D3525_Y),     .Y(D3583_Y));
KC_OAI21B_X1 D3291 ( .A1(D3223_Y), .B(D3217_Y), .A0N(D3259_Y),     .Y(D3291_Y));
KC_OAI21B_X1 D3290 ( .A1(D3259_Y), .B(D3207_Y), .A0N(D3052_Y),     .Y(D3290_Y));
KC_OAI21B_X1 D3193 ( .A1(D3155_Y), .B(D3094_Y), .A0N(D4607_Y),     .Y(D3193_Y));
KC_OAI21B_X1 D3091 ( .A1(D4525_Y), .B(D32_Y), .A0N(D316_Y),     .Y(D3091_Y));
KC_OAI21B_X1 D1961 ( .A1(D1835_Y), .B(D8029_Y), .A0N(D8401_Y),     .Y(D1961_Y));
KC_OAI21B_X1 D1960 ( .A1(D1828_Y), .B(D1888_Y), .A0N(D105_Y),     .Y(D1960_Y));
KC_OAI21B_X1 D1667 ( .A1(D1648_Y), .B(D309_Y), .A0N(D4505_Y),     .Y(D1667_Y));
KC_OAI21B_X1 D487 ( .A1(D469_Y), .B(D435_Y), .A0N(D479_Q), .Y(D487_Y));
KC_OAI21B_X1 D391 ( .A1(D4728_Q), .B(D3255_Y), .A0N(D372_Y),     .Y(D391_Y));
KC_OAI21B_X1 D390 ( .A1(D2995_Y), .B(D4717_Y), .A0N(D3268_Y),     .Y(D390_Y));
KC_OAI21BB_X1 D16477 ( .Y(D16477_Y), .B(D16483_Q), .C(D16467_Y),     .A(D16410_Y));
KC_OAI21BB_X1 D14521 ( .Y(D14521_Y), .B(D14548_Y), .C(D14532_Y),     .A(D2512_Y));
KC_OAI21BB_X1 D12751 ( .Y(D12751_Y), .B(D12738_Y), .C(D13234_Y),     .A(D13220_Y));
KC_OAI21BB_X1 D11588 ( .Y(D11588_Y), .B(D8472_Y), .C(D11535_Y),     .A(D6792_Y));
KC_OAI21BB_X1 D11587 ( .Y(D11587_Y), .B(D6792_Y), .C(D11535_Y),     .A(D8472_Y));
KC_OAI21BB_X1 D11415 ( .Y(D11415_Y), .B(D8302_Y), .C(D11386_Y),     .A(D6792_Y));
KC_OAI21BB_X1 D11414 ( .Y(D11414_Y), .B(D6792_Y), .C(D11386_Y),     .A(D8302_Y));
KC_OAI21BB_X1 D11348 ( .Y(D11348_Y), .B(D6792_Y), .C(D11256_Y),     .A(D1961_Y));
KC_OAI21BB_X1 D11052 ( .Y(D11052_Y), .B(D6792_Y), .C(D11536_Y),     .A(D8473_Y));
KC_OAI21BB_X1 D10894 ( .Y(D10894_Y), .B(D1961_Y), .C(D11256_Y),     .A(D6792_Y));
KC_OAI21BB_X1 D8552 ( .Y(D8552_Y), .B(D2032_Y), .C(D1891_Y),     .A(D5508_Y));
KC_OAI21BB_X1 D8255 ( .Y(D8255_Y), .B(D6759_Y), .C(D1899_Y),     .A(D6709_Y));
KC_OAI21BB_X1 D7897 ( .Y(D7897_Y), .B(D7878_Y), .C(D7874_Y),     .A(D7842_Y));
KC_OAI21BB_X1 D7808 ( .Y(D7808_Y), .B(D1453_Y), .C(D4659_Y),     .A(D450_Q));
KC_OAI21BB_X1 D7803 ( .Y(D7803_Y), .B(D1453_Y), .C(D4659_Y),     .A(D7791_Q));
KC_OAI21BB_X1 D7800 ( .Y(D7800_Y), .B(D1453_Y), .C(D4655_Y),     .A(D7790_Q));
KC_OAI21BB_X1 D7799 ( .Y(D7799_Y), .B(D1453_Y), .C(D4655_Y),     .A(D7789_Q));
KC_OAI21BB_X1 D7536 ( .Y(D7536_Y), .B(D7508_Y), .C(D7416_Y),     .A(D7534_Q));
KC_OAI21BB_X1 D7535 ( .Y(D7535_Y), .B(D5966_Y), .C(D7508_Y),     .A(D8730_Q));
KC_OAI21BB_X1 D7397 ( .Y(D7397_Y), .B(D5768_Y), .C(D5916_Y),     .A(D7333_Y));
KC_OAI21BB_X1 D6831 ( .Y(D6831_Y), .B(D8031_Y), .C(D5391_Y),     .A(D6260_Y));
KC_OAI21BB_X1 D5938 ( .Y(D5938_Y), .B(D5651_Y), .C(D5863_Y),     .A(D5997_Y));
KC_OAI21BB_X1 D5816 ( .Y(D5816_Y), .B(D5877_Y), .C(D213_Y),     .A(D5856_Y));
KC_OAI21BB_X1 D5249 ( .Y(D5249_Y), .B(D6792_Y), .C(D5215_Y),     .A(D561_Y));
KC_OAI21BB_X1 D4026 ( .Y(D4026_Y), .B(D8471_Y), .C(D5558_Y),     .A(D6260_Y));
KC_OAI21BB_X1 D3888 ( .Y(D3888_Y), .B(D6260_Y), .C(D3862_Y),     .A(D8309_Y));
KC_OAI21BB_X1 D3887 ( .Y(D3887_Y), .B(D8309_Y), .C(D3862_Y),     .A(D6260_Y));
KC_OAI21BB_X1 D3761 ( .Y(D3761_Y), .B(D561_Y), .C(D5215_Y),     .A(D6792_Y));
KC_OAI21BB_X1 D2894 ( .Y(D2894_Y), .B(D2887_Q), .C(D2854_Y),     .A(D2827_Y));
KC_OAI21BB_X1 D2803 ( .Y(D2803_Y), .B(D2805_Y), .C(D2766_Y),     .A(D2814_Q));
KC_OAI21BB_X1 D2259 ( .Y(D2259_Y), .B(D6792_Y), .C(D11258_Y),     .A(D8258_Y));
KC_OAI21BB_X1 D2258 ( .Y(D2258_Y), .B(D8258_Y), .C(D11258_Y),     .A(D6792_Y));
KC_OAI21BB_X1 D2101 ( .Y(D2101_Y), .B(D9523_Y), .C(D825_Q),     .A(D1985_Y));
KC_OAI21BB_X1 D1666 ( .Y(D1666_Y), .B(D4926_Y), .C(D4968_Y),     .A(D4927_Y));
KC_OAI21BB_X1 D1523 ( .Y(D1523_Y), .B(D6260_Y), .C(D6958_Y),     .A(D8471_Y));
KC_OAI21BB_X1 D456 ( .Y(D456_Y), .B(D1453_Y), .C(D4697_Y),     .A(D7794_Q));
KC_OAI21BB_X1 D455 ( .Y(D455_Y), .B(D1453_Y), .C(D4655_Y),     .A(D7793_Q));
KC_OAI21BB_X1 D424 ( .Y(D424_Y), .B(D10079_Y), .C(D7683_Y),     .A(D9218_Q));
KC_OAI21BB_X1 D423 ( .Y(D423_Y), .B(D10079_Y), .C(D9101_Y),     .A(D419_Q));
KC_OAI21BB_X1 D422 ( .Y(D422_Y), .B(D10079_Y), .C(D9180_Y),     .A(D10108_Q));
KC_OAI21BB_X1 D389 ( .Y(D389_Y), .B(D10079_Y), .C(D9175_Y),     .A(D9148_Q));
KC_OR2_X1 D16672 ( .Y(D16672_Y), .B(D16677_Q), .A(D16682_Q));
KC_OR2_X1 D16546 ( .Y(D16546_Y), .B(D16549_Y), .A(D16654_Y));
KC_OR2_X1 D16511 ( .Y(D16511_Y), .B(D16501_Y), .A(D16484_Y));
KC_OR2_X1 D16506 ( .Y(D16506_Y), .B(D16490_Y), .A(D16484_Y));
KC_OR2_X1 D16451 ( .Y(D16451_Y), .B(D16457_Y), .A(D16375_Y));
KC_OR2_X1 D16193 ( .Y(D16193_Y), .B(D16190_Y), .A(D16379_Y));
KC_OR2_X1 D15122 ( .Y(D15122_Y), .B(D15089_Y), .A(D15170_Y));
KC_OR2_X1 D15111 ( .Y(D15111_Y), .B(D1177_Y), .A(D1275_Y));
KC_OR2_X1 D14775 ( .Y(D14775_Y), .B(D13392_Y), .A(D14807_Y));
KC_OR2_X1 D14667 ( .Y(D14667_Y), .B(D14630_Y), .A(D14629_Y));
KC_OR2_X1 D14566 ( .Y(D14566_Y), .B(D14547_Y), .A(D14560_Y));
KC_OR2_X1 D14365 ( .Y(D14365_Y), .B(D14324_Y), .A(D14328_Y));
KC_OR2_X1 D14363 ( .Y(D14363_Y), .B(D14327_Y), .A(D14437_Y));
KC_OR2_X1 D14287 ( .Y(D14287_Y), .B(D14274_Y), .A(D14285_Y));
KC_OR2_X1 D13971 ( .Y(D13971_Y), .B(D13975_Y), .A(D12690_Y));
KC_OR2_X1 D13736 ( .Y(D13736_Y), .B(D13725_Y), .A(D13747_Y));
KC_OR2_X1 D13245 ( .Y(D13245_Y), .B(D12195_Y), .A(D2407_Y));
KC_OR2_X1 D12663 ( .Y(D12663_Y), .B(D16_Y), .A(D6342_Y));
KC_OR2_X1 D12136 ( .Y(D12136_Y), .B(D12183_Y), .A(D2304_Q));
KC_OR2_X1 D11649 ( .Y(D11649_Y), .B(D12197_Y), .A(D11651_Y));
KC_OR2_X1 D11616 ( .Y(D11616_Y), .B(D7401_Y), .A(D7404_Y));
KC_OR2_X1 D10863 ( .Y(D10863_Y), .B(D10807_Y), .A(D10864_Y));
KC_OR2_X1 D10091 ( .Y(D10091_Y), .B(D10078_Y), .A(D9104_Y));
KC_OR2_X1 D9540 ( .Y(D9540_Y), .B(D9583_Y), .A(D9524_Y));
KC_OR2_X1 D9434 ( .Y(D9434_Y), .B(D9436_Y), .A(D9469_Y));
KC_OR2_X1 D9432 ( .Y(D9432_Y), .B(D9407_Y), .A(D9404_Y));
KC_OR2_X1 D9130 ( .Y(D9130_Y), .B(D9119_Y), .A(D9123_Y));
KC_OR2_X1 D8990 ( .Y(D8990_Y), .B(D8701_Y), .A(D9025_Y));
KC_OR2_X1 D8989 ( .Y(D8989_Y), .B(D7490_Y), .A(D9025_Y));
KC_OR2_X1 D8927 ( .Y(D8927_Y), .B(D9122_Y), .A(D7485_Y));
KC_OR2_X1 D8882 ( .Y(D8882_Y), .B(D8952_Q), .A(D8050_Y));
KC_OR2_X1 D8775 ( .Y(D8775_Y), .B(D8798_S), .A(D7427_Y));
KC_OR2_X1 D8686 ( .Y(D8686_Y), .B(D8729_Y), .A(D8729_Y));
KC_OR2_X1 D8219 ( .Y(D8219_Y), .B(D8239_Y), .A(D1840_Y));
KC_OR2_X1 D7952 ( .Y(D7952_Y), .B(D7921_Y), .A(D7943_Y));
KC_OR2_X1 D7640 ( .Y(D7640_Y), .B(D6215_Y), .A(D7649_Y));
KC_OR2_X1 D7453 ( .Y(D7453_Y), .B(D4490_Q), .A(D268_Q));
KC_OR2_X1 D7370 ( .Y(D7370_Y), .B(D1716_Y), .A(D7389_Y));
KC_OR2_X1 D7123 ( .Y(D7123_Y), .B(D6333_Y), .A(D7120_Y));
KC_OR2_X1 D6880 ( .Y(D6880_Y), .B(D8371_Y), .A(D970_Y));
KC_OR2_X1 D6370 ( .Y(D6370_Y), .B(D4962_Y), .A(D6441_Y));
KC_OR2_X1 D6235 ( .Y(D6235_Y), .B(D13173_Y), .A(D9144_Y));
KC_OR2_X1 D6158 ( .Y(D6158_Y), .B(D6138_Y), .A(D6156_Y));
KC_OR2_X1 D6106 ( .Y(D6106_Y), .B(D6089_Y), .A(D7515_Y));
KC_OR2_X1 D5787 ( .Y(D5787_Y), .B(D1728_Y), .A(D5788_Y));
KC_OR2_X1 D4700 ( .Y(D4700_Y), .B(D4678_Y), .A(D6329_Y));
KC_OR2_X1 D4699 ( .Y(D4699_Y), .B(D4702_Y), .A(D4766_Y));
KC_OR2_X1 D4698 ( .Y(D4698_Y), .B(D4844_Y), .A(D4700_Y));
KC_OR2_X1 D4526 ( .Y(D4526_Y), .B(D3069_Y), .A(D4566_Q));
KC_OR2_X1 D4363 ( .Y(D4363_Y), .B(D4292_Y), .A(D6034_Y));
KC_OR2_X1 D3339 ( .Y(D3339_Y), .B(D3306_Y), .A(D3308_Y));
KC_OR2_X1 D3253 ( .Y(D3253_Y), .B(D3283_Q), .A(D3281_Q));
KC_OR2_X1 D3249 ( .Y(D3249_Y), .B(D3263_Y), .A(D3224_Y));
KC_OR2_X1 D3242 ( .Y(D3242_Y), .B(D3291_Y), .A(D1469_Y));
KC_OR2_X1 D3155 ( .Y(D3155_Y), .B(D8152_Y), .A(D352_Y));
KC_OR2_X1 D2952 ( .Y(D2952_Y), .B(D2955_Y), .A(D2997_Y));
KC_OR2_X1 D2856 ( .Y(D2856_Y), .B(D2867_Y), .A(D2880_Y));
KC_OR2_X1 D2855 ( .Y(D2855_Y), .B(D2868_Y), .A(D2826_Y));
KC_OR2_X1 D2777 ( .Y(D2777_Y), .B(D2753_Y), .A(D2754_Y));
KC_OR2_X1 D2773 ( .Y(D2773_Y), .B(D2736_Y), .A(D2745_Y));
KC_OR2_X1 D2630 ( .Y(D2630_Y), .B(D15334_Y), .A(D15395_Y));
KC_OR2_X1 D2629 ( .Y(D2629_Y), .B(D15327_Y), .A(D2593_Y));
KC_OR2_X1 D2565 ( .Y(D2565_Y), .B(D2630_Y), .A(D15443_Y));
KC_OR2_X1 D2501 ( .Y(D2501_Y), .B(D2494_Y), .A(D14216_Y));
KC_OR2_X1 D2499 ( .Y(D2499_Y), .B(D2486_Y), .A(D14281_Y));
KC_OR2_X1 D1747 ( .Y(D1747_Y), .B(D6132_Y), .A(D6201_Y));
KC_OR2_X1 D1743 ( .Y(D1743_Y), .B(D8393_Y), .A(D7830_Y));
KC_OR2_X1 D1611 ( .Y(D1611_Y), .B(D309_Y), .A(D1667_Y));
KC_OR2_X1 D1459 ( .Y(D1459_Y), .B(D2821_Y), .A(D2885_Q));
KC_OR2_X1 D1457 ( .Y(D1457_Y), .B(D1432_Y), .A(D3187_Q));
KC_OR2_X1 D1404 ( .Y(D1404_Y), .B(D16588_Y), .A(D16585_Y));
KC_OR2_X1 D1188 ( .Y(D1188_Y), .B(D15091_Y), .A(D15966_Y));
KC_OR2_X1 D999 ( .Y(D999_Y), .B(D2493_Y), .A(D14221_Y));
KC_OR2_X1 D374 ( .Y(D374_Y), .B(D9148_Q), .A(D10108_Q));
KC_MXI2_X10 D327 ( .Y(D327_Y), .AN(D15250_Y), .B(D15276_Y),     .S0(D14586_Y));
KC_MXI2_X10 D16199 ( .Y(D16199_Y), .AN(D2658_Y), .B(D13345_Y),     .S0(D13268_Q));
KC_MXI2_X10 D16197 ( .Y(D16197_Y), .AN(D8352_Y), .B(D6786_Y),     .S0(D6773_Y));
KC_MXI2_X10 D16164 ( .Y(D16164_Y), .AN(D10753_Q), .B(D8111_Y),     .S0(D9426_Y));
KC_MXI2_X10 D16156 ( .Y(D16156_Y), .AN(D6313_Y), .B(D6343_Y),     .S0(D6355_Y));
KC_MXI2_X10 D16147 ( .Y(D16147_Y), .AN(D6267_Y), .B(D6224_Y),     .S0(D6266_Y));
KC_MXI2_X10 D16143 ( .Y(D16143_Y), .AN(D6086_Y), .B(D7531_Y),     .S0(D6100_Y));
KC_MXI2_X10 D16135 ( .Y(D16135_Y), .AN(D4123_Y), .B(D4103_Y),     .S0(D4104_Y));
KC_MXI2_X10 D16006 ( .Y(D16006_Y), .AN(D3458_Y), .B(D1531_Y),     .S0(D3598_Co));
KC_MXI2_X10 D15265 ( .Y(D15265_Y), .AN(D3314_Y), .B(D3377_Y),     .S0(D3315_Y));
KC_MXI2_X10 D13098 ( .Y(D13098_Y), .AN(D2896_Q), .B(D2766_Y),     .S0(D1477_Y));
KC_MXI2_X10 D10144 ( .Y(D10144_Y), .AN(D6475_Q), .B(D6416_Y),     .S0(D7935_Y));
KC_MXI2_X10 D9326 ( .Y(D9326_Y), .AN(D15534_Y), .B(D15567_Y),     .S0(D15362_Y));
KC_MXI2_X10 D8152 ( .Y(D8152_Y), .AN(D3161_Y), .B(D3181_Y),     .S0(D3171_S));
KC_AO21_X2 D16185 ( .B(D16124_Y), .A1(D16088_Y), .Y(D16185_Y),     .A0(D16066_Y));
KC_AO21_X2 D16174 ( .B(D16127_Y), .A1(D2673_Y), .Y(D16174_Y),     .A0(D16101_Y));
KC_AO21_X2 D16173 ( .B(D2682_Y), .A1(D16169_Y), .Y(D16173_Y),     .A0(D2652_Y));
KC_AO21_X2 D14908 ( .B(D13983_Y), .A1(D14169_Q), .Y(D14908_Y),     .A0(D14094_Q));
KC_AO21_X2 D14707 ( .B(D14661_Y), .A1(D13958_Y), .Y(D14707_Y),     .A0(D14662_Y));
KC_AO21_X2 D14599 ( .B(D14545_Y), .A1(D2570_Y), .Y(D14599_Y),     .A0(D2512_Y));
KC_AO21_X2 D13919 ( .B(D13878_Y), .A1(D8886_Y), .Y(D13919_Y),     .A0(D2509_Y));
KC_AO21_X2 D13917 ( .B(D13888_Y), .A1(D15438_Y), .Y(D13917_Y),     .A0(D2509_Y));
KC_AO21_X2 D13916 ( .B(D13885_Y), .A1(D9553_Y), .Y(D13916_Y),     .A0(D2509_Y));
KC_AO21_X2 D13915 ( .B(D13896_Y), .A1(D16139_Y), .Y(D13915_Y),     .A0(D2509_Y));
KC_AO21_X2 D13914 ( .B(D13893_Y), .A1(D16132_Y), .Y(D13914_Y),     .A0(D2509_Y));
KC_AO21_X2 D13913 ( .B(D13879_Y), .A1(D15437_Y), .Y(D13913_Y),     .A0(D2509_Y));
KC_AO21_X2 D12690 ( .B(D13216_Q), .A1(D396_Y), .Y(D12690_Y),     .A0(D6342_Y));
KC_AO21_X2 D11671 ( .B(D11645_Y), .A1(D11649_Y), .Y(D11671_Y),     .A0(D10181_Y));
KC_AO21_X2 D9386 ( .B(D9383_Y), .A1(D9367_Y), .Y(D9386_Y),     .A0(D9380_Y));
KC_AO21_X2 D8728 ( .B(D8717_Y), .A1(D8672_Y), .Y(D8728_Y),     .A0(D1977_Y));
KC_AO21_X2 D8353 ( .B(D8338_Y), .A1(D942_Y), .Y(D8353_Y),     .A0(D8281_Y));
KC_AO21_X2 D7983 ( .B(D7972_Y), .A1(D545_Y), .Y(D7983_Y),     .A0(D7935_Y));
KC_AO21_X2 D7982 ( .B(D7837_Y), .A1(D7978_Y), .Y(D7982_Y),     .A0(D7966_Q));
KC_AO21_X2 D7981 ( .B(D7837_Y), .A1(D7906_Y), .Y(D7981_Y),     .A0(D7968_Q));
KC_AO21_X2 D7748 ( .B(D7695_Y), .A1(D1865_Y), .Y(D7748_Y),     .A0(D7735_Q));
KC_AO21_X2 D7747 ( .B(D7694_Y), .A1(D1865_Y), .Y(D7747_Y),     .A0(D7745_Q));
KC_AO21_X2 D7746 ( .B(D7695_Y), .A1(D1865_Y), .Y(D7746_Y),     .A0(D7734_Q));
KC_AO21_X2 D7612 ( .B(D7582_Y), .A1(D7574_Y), .Y(D7612_Y),     .A0(D7555_Y));
KC_AO21_X2 D7487 ( .B(D7459_Y), .A1(D15448_Y), .Y(D7487_Y),     .A0(D7417_Y));
KC_AO21_X2 D7160 ( .B(D182_Y), .A1(D7114_Y), .Y(D7160_Y),     .A0(D7127_Y));
KC_AO21_X2 D6202 ( .B(D6253_Y), .A1(D6182_Y), .Y(D6202_Y),     .A0(D6117_Y));
KC_AO21_X2 D4250 ( .B(D4178_Y), .A1(D5973_Y), .Y(D4250_Y),     .A0(D5752_Y));
KC_AO21_X2 D4088 ( .B(D4032_Y), .A1(D4076_Y), .Y(D4088_Y),     .A0(D4078_Y));
KC_AO21_X2 D4068 ( .B(D4033_Y), .A1(D4078_Y), .Y(D4068_Y),     .A0(D4076_Y));
KC_AO21_X2 D3396 ( .B(D3390_Y), .A1(D3353_Y), .Y(D3396_Y),     .A0(D3352_Y));
KC_AO21_X2 D3194 ( .B(D3150_Y), .A1(D1468_Y), .Y(D3194_Y),     .A0(D3128_Y));
KC_AO21_X2 D3008 ( .B(D2990_Y), .A1(D2911_Y), .Y(D3008_Y),     .A0(D2989_Y));
KC_AO21_X2 D2899 ( .B(D2852_Y), .A1(D1440_Y), .Y(D2899_Y),     .A0(D2902_Q));
KC_AO21_X2 D2585 ( .B(D2565_Y), .A1(D15443_Y), .Y(D2585_Y),     .A0(D2630_Y));
KC_AO21_X2 D1967 ( .B(D1847_Y), .A1(D8030_Y), .Y(D1967_Y),     .A0(D7973_Q));
KC_AO21_X2 D1966 ( .B(D1770_Y), .A1(D1935_Y), .Y(D1966_Y),     .A0(D1935_Y));
KC_AO21_X2 D1965 ( .B(D7694_Y), .A1(D1865_Y), .Y(D1965_Y),     .A0(D7736_Q));
KC_AO21_X2 D366 ( .B(D4504_Y), .A1(D3169_Y), .Y(D366_Y), .A0(D4611_Y));
KC_NAND2_X4 D15955 ( .Y(D15955_Y), .B(D15954_Y), .A(D15953_Y));
KC_NAND2_X4 D15952 ( .Y(D15952_Y), .B(D15950_Y), .A(D15951_Y));
KC_NAND2_X4 D15877 ( .Y(D15877_Y), .B(D15876_Y), .A(D15875_Y));
KC_NAND2_X4 D15806 ( .Y(D15806_Y), .B(D15804_Y), .A(D15805_Y));
KC_NAND2_X4 D15803 ( .Y(D15803_Y), .B(D15802_Y), .A(D15801_Y));
KC_NAND2_X4 D15800 ( .Y(D15800_Y), .B(D15799_Y), .A(D15798_Y));
KC_NAND2_X4 D15680 ( .Y(D15680_Y), .B(D15679_Y), .A(D938_Y));
KC_NAND2_X4 D15678 ( .Y(D15678_Y), .B(D15677_Y), .A(D15676_Y));
KC_NAND2_X4 D15674 ( .Y(D15674_Y), .B(D937_Y), .A(D15675_Y));
KC_NAND2_X4 D15673 ( .Y(D15673_Y), .B(D15672_Y), .A(D15671_Y));
KC_NAND2_X4 D15581 ( .Y(D15581_Y), .B(D15579_Y), .A(D15578_Y));
KC_NAND2_X4 D15576 ( .Y(D15576_Y), .B(D15574_Y), .A(D15570_Y));
KC_NAND2_X4 D15575 ( .Y(D15575_Y), .B(D15573_Y), .A(D15571_Y));
KC_NAND2_X4 D15569 ( .Y(D15569_Y), .B(D832_Y), .A(D15572_Y));
KC_NAND2_X4 D15149 ( .Y(D15149_Y), .B(D15147_Y), .A(D15148_Y));
KC_NAND2_X4 D15146 ( .Y(D15146_Y), .B(D15145_Y), .A(D1239_Y));
KC_NAND2_X4 D15082 ( .Y(D15082_Y), .B(D15080_Y), .A(D15081_Y));
KC_NAND2_X4 D15079 ( .Y(D15079_Y), .B(D15077_Y), .A(D15078_Y));
KC_NAND2_X4 D15076 ( .Y(D15076_Y), .B(D15074_Y), .A(D15075_Y));
KC_NAND2_X4 D15003 ( .Y(D15003_Y), .B(D15001_Y), .A(D15002_Y));
KC_NAND2_X4 D15000 ( .Y(D15000_Y), .B(D14998_Y), .A(D14999_Y));
KC_NAND2_X4 D14902 ( .Y(D14902_Y), .B(D14900_Y), .A(D14901_Y));
KC_NAND2_X4 D14899 ( .Y(D14899_Y), .B(D14897_Y), .A(D14893_Y));
KC_NAND2_X4 D14898 ( .Y(D14898_Y), .B(D14896_Y), .A(D14894_Y));
KC_NAND2_X4 D14892 ( .Y(D14892_Y), .B(D14890_Y), .A(D14891_Y));
KC_NAND2_X4 D14889 ( .Y(D14889_Y), .B(D14888_Y), .A(D14887_Y));
KC_NAND2_X4 D14799 ( .Y(D14799_Y), .B(D14797_Y), .A(D14798_Y));
KC_NAND2_X4 D14796 ( .Y(D14796_Y), .B(D14795_Y), .A(D14794_Y));
KC_NAND2_X4 D14381 ( .Y(D14381_Y), .B(D14379_Y), .A(D14376_Y));
KC_NAND2_X4 D14396 ( .Y(D14396_Y), .B(D14393_Y), .A(D14395_Y));
KC_NAND2_X4 D14392 ( .Y(D14392_Y), .B(D14394_Y), .A(D14391_Y));
KC_NAND2_X4 D14390 ( .Y(D14390_Y), .B(D14389_Y), .A(D14388_Y));
KC_NAND2_X4 D14387 ( .Y(D14387_Y), .B(D14383_Y), .A(D14385_Y));
KC_NAND2_X4 D14386 ( .Y(D14386_Y), .B(D14382_Y), .A(D14384_Y));
KC_NAND2_X4 D14380 ( .Y(D14380_Y), .B(D14378_Y), .A(D14377_Y));
KC_NAND2_X4 D14314 ( .Y(D14314_Y), .B(D14312_Y), .A(D14313_Y));
KC_NAND2_X4 D14311 ( .Y(D14311_Y), .B(D14309_Y), .A(D14310_Y));
KC_NAND2_X4 D14262 ( .Y(D14262_Y), .B(D14260_Y), .A(D14261_Y));
KC_NAND2_X4 D14192 ( .Y(D14192_Y), .B(D14189_Y), .A(D939_Y));
KC_NAND2_X4 D14191 ( .Y(D14191_Y), .B(D14190_Y), .A(D14188_Y));
KC_NAND2_X4 D14187 ( .Y(D14187_Y), .B(D14185_Y), .A(D14186_Y));
KC_NAND2_X4 D14184 ( .Y(D14184_Y), .B(D14182_Y), .A(D14183_Y));
KC_NAND2_X4 D14181 ( .Y(D14181_Y), .B(D14179_Y), .A(D14180_Y));
KC_NAND2_X4 D11668 ( .Y(D11668_Y), .B(D11667_Y), .A(D11666_Y));
KC_NAND2_X4 D9334 ( .Y(D9334_Y), .B(D9335_Y), .A(D9329_Y));
KC_NAND2_X4 D9333 ( .Y(D9333_Y), .B(D9327_Y), .A(D9331_Y));
KC_NAND2_X4 D9332 ( .Y(D9332_Y), .B(D9330_Y), .A(D9328_Y));
KC_NAND2_X4 D9158 ( .Y(D9158_Y), .B(D9156_Y), .A(D9157_Y));
KC_NAND2_X4 D9155 ( .Y(D9155_Y), .B(D9153_Y), .A(D9154_Y));
KC_NAND2_X4 D8958 ( .Y(D8958_Y), .B(D8956_Y), .A(D8957_Y));
KC_NAND2_X4 D8721 ( .Y(D8721_Y), .B(D8720_Y), .A(D8719_Y));
KC_NAND2_X4 D8253 ( .Y(D8253_Y), .B(D8252_Y), .A(D8251_Y));
KC_NAND2_X4 D7666 ( .Y(D7666_Y), .B(D7665_Y), .A(D7664_Y));
KC_NAND2_X4 D7662 ( .Y(D7662_Y), .B(D7663_Y), .A(D7661_Y));
KC_NAND2_X4 D7608 ( .Y(D7608_Y), .B(D7606_Y), .A(D7607_Y));
KC_NAND2_X4 D7604 ( .Y(D7604_Y), .B(D7611_Y), .A(D7602_Y));
KC_NAND2_X4 D7603 ( .Y(D7603_Y), .B(D7600_Y), .A(D7601_Y));
KC_NAND2_X4 D7599 ( .Y(D7599_Y), .B(D7598_Y), .A(D7597_Y));
KC_NAND2_X4 D7595 ( .Y(D7595_Y), .B(D7593_Y), .A(D7594_Y));
KC_NAND2_X4 D7592 ( .Y(D7592_Y), .B(D7590_Y), .A(D7591_Y));
KC_NAND2_X4 D7158 ( .Y(D7158_Y), .B(D7157_Y), .A(D197_Y));
KC_NAND2_X4 D7156 ( .Y(D7156_Y), .B(D7155_Y), .A(D7154_Y));
KC_NAND2_X4 D6348 ( .Y(D6348_Y), .B(D6346_Y), .A(D6347_Y));
KC_NAND2_X4 D6271 ( .Y(D6271_Y), .B(D388_Y), .A(D6270_Y));
KC_NAND2_X4 D6194 ( .Y(D6194_Y), .B(D6192_Y), .A(D6193_Y));
KC_NAND2_X4 D6191 ( .Y(D6191_Y), .B(D359_Y), .A(D6190_Y));
KC_NAND2_X4 D6188 ( .Y(D6188_Y), .B(D357_Y), .A(D6187_Y));
KC_NAND2_X4 D4127 ( .Y(D4127_Y), .B(D4126_Y), .A(D4125_Y));
KC_NAND2_X4 D3582 ( .Y(D3582_Y), .B(D5081_Y), .A(D3581_Y));
KC_NAND2_X4 D3287 ( .Y(D3287_Y), .B(D3286_Y), .A(D3285_Y));
KC_NAND2_X4 D3086 ( .Y(D3086_Y), .B(D3089_Y), .A(D3088_Y));
KC_NAND2_X4 D2647 ( .Y(D2647_Y), .B(D2646_Y), .A(D2645_Y));
KC_NAND2_X4 D2644 ( .Y(D2644_Y), .B(D2642_Y), .A(D2643_Y));
KC_NAND2_X4 D2583 ( .Y(D2583_Y), .B(D2581_Y), .A(D2582_Y));
KC_NAND2_X4 D2579 ( .Y(D2579_Y), .B(D2580_Y), .A(D2577_Y));
KC_NAND2_X4 D2578 ( .Y(D2578_Y), .B(D2576_Y), .A(D2575_Y));
KC_NAND2_X4 D2521 ( .Y(D2521_Y), .B(D2520_Y), .A(D158_Y));
KC_NAND2_X4 D2098 ( .Y(D2098_Y), .B(D2097_Y), .A(D2096_Y));
KC_NAND2_X4 D1952 ( .Y(D1952_Y), .B(D1950_Y), .A(D1951_Y));
KC_NAND2_X4 D1949 ( .Y(D1949_Y), .B(D159_Y), .A(D1948_Y));
KC_NAND2_X4 D1804 ( .Y(D1804_Y), .B(D1802_Y), .A(D1803_Y));
KC_NAND2_X4 D940 ( .Y(D940_Y), .B(D14895_Y), .A(D15681_Y));
KC_NAND2_X4 D360 ( .Y(D360_Y), .B(D7605_Y), .A(D6195_Y));
KC_NAND2_X4 D358 ( .Y(D358_Y), .B(D7596_Y), .A(D6189_Y));
KC_XOR2_X3 D16736 ( .Y(D16736_Y), .B(D16772_Y), .A(D16709_Y));
KC_XOR2_X3 D16735 ( .Y(D16735_Y), .B(D16772_Y), .A(D16708_Y));
KC_XOR2_X3 D16734 ( .Y(D16734_Y), .B(D16715_Y), .A(D16730_Y));
KC_XOR2_X3 D16733 ( .Y(D16733_Y), .B(D16715_Y), .A(D16729_Y));
KC_XOR2_X3 D16397 ( .Y(D16397_Y), .B(D16588_Y), .A(D16591_Y));
KC_XOR2_X3 D16396 ( .Y(D16396_Y), .B(D16639_Y), .A(D16617_Y));
KC_XOR2_X3 D16395 ( .Y(D16395_Y), .B(D16588_Y), .A(D16583_Y));
KC_XOR2_X3 D16394 ( .Y(D16394_Y), .B(D16639_Y), .A(D16633_Y));
KC_XOR2_X3 D16328 ( .Y(D16328_Y), .B(D16341_Y), .A(D16330_Y));
KC_XOR2_X3 D16320 ( .Y(D16320_Y), .B(D16341_Y), .A(D16329_Y));
KC_XOR2_X3 D15139 ( .Y(D15139_Y), .B(D15159_Y), .A(D15151_Y));
KC_XOR2_X3 D15138 ( .Y(D15138_Y), .B(D15159_Y), .A(D15150_Y));
KC_XOR2_X3 D14694 ( .Y(D14694_Y), .B(D2585_Y), .A(D2585_Y));
KC_XOR2_X3 D14692 ( .Y(D14692_Y), .B(D14712_Y), .A(D14699_Y));
KC_XOR2_X3 D14690 ( .Y(D14690_Y), .B(D14712_Y), .A(D14700_Y));
KC_XOR2_X3 D13767 ( .Y(D13767_Y), .B(D13843_Y), .A(D13835_Y));
KC_XOR2_X3 D13766 ( .Y(D13766_Y), .B(D13843_Y), .A(D13834_Y));
KC_XOR2_X3 D13616 ( .Y(D13616_Y), .B(D1076_Y), .A(D13621_Y));
KC_XOR2_X3 D12547 ( .Y(D12547_Y), .B(D13094_Y), .A(D1241_Y));
KC_XOR2_X3 D12363 ( .Y(D12363_Y), .B(D12304_Y), .A(D12289_Y));
KC_XOR2_X3 D12286 ( .Y(D12286_Y), .B(D12304_Y), .A(D12290_Y));
KC_XOR2_X3 D12049 ( .Y(D12049_Y), .B(D11612_Y), .A(D1390_Y));
KC_XOR2_X3 D11540 ( .Y(D11540_Y), .B(D11612_Y), .A(D11605_Y));
KC_XOR2_X3 D11410 ( .Y(D11410_Y), .B(D11417_Y), .A(D11412_Y));
KC_XOR2_X3 D11409 ( .Y(D11409_Y), .B(D11417_Y), .A(D2262_Y));
KC_XOR2_X3 D11045 ( .Y(D11045_Y), .B(D11055_Y), .A(D11049_Y));
KC_XOR2_X3 D11039 ( .Y(D11039_Y), .B(D11055_Y), .A(D11048_Y));
KC_XOR2_X3 D9849 ( .Y(D9849_Y), .B(D8663_Y), .A(D9917_Y));
KC_XOR2_X3 D9223 ( .Y(D9223_Y), .B(D7691_Y), .A(D9259_Y));
KC_XOR2_X3 D9222 ( .Y(D9222_Y), .B(D2003_Y), .A(D9250_Y));
KC_XOR2_X3 D9025 ( .Y(D9025_Y), .B(D7490_Y), .A(D8701_Y));
KC_XOR2_X3 D8716 ( .Y(D8716_Y), .B(D8685_Y), .A(D8674_Y));
KC_XOR2_X3 D8602 ( .Y(D8602_Y), .B(D8607_Y), .A(D8604_Y));
KC_XOR2_X3 D8596 ( .Y(D8596_Y), .B(D8607_Y), .A(D8603_Y));
KC_XOR2_X3 D8164 ( .Y(D8164_Y), .B(D16753_Y), .A(D710_Y));
KC_XOR2_X3 D7589 ( .Y(D7589_Y), .B(D7555_Y), .A(D7559_Y));
KC_XOR2_X3 D7588 ( .Y(D7588_Y), .B(D7646_Y), .A(D7628_Y));
KC_XOR2_X3 D6556 ( .Y(D6556_Y), .B(D16696_Y), .A(D6562_Y));
KC_XOR2_X3 D6482 ( .Y(D6482_Y), .B(D6531_Y), .A(D6477_Y));
KC_XOR2_X3 D6392 ( .Y(D6392_Y), .B(D14591_Y), .A(D6400_Y));
KC_XOR2_X3 D6391 ( .Y(D6391_Y), .B(D14591_Y), .A(D6399_Y));
KC_XOR2_X3 D6267 ( .Y(D6267_Y), .B(D6247_Y), .A(D6221_Y));
KC_XOR2_X3 D6185 ( .Y(D6185_Y), .B(D4719_Y), .A(D7561_Y));
KC_XOR2_X3 D6123 ( .Y(D6123_Y), .B(D6128_Y), .A(D6125_Y));
KC_XOR2_X3 D5806 ( .Y(D5806_Y), .B(D6275_Y), .A(D5813_Y));
KC_XOR2_X3 D5485 ( .Y(D5485_Y), .B(D5489_Y), .A(D5488_Y));
KC_XOR2_X3 D5412 ( .Y(D5412_Y), .B(D5360_Y), .A(D5295_Y));
KC_XOR2_X3 D4645 ( .Y(D4645_Y), .B(D6197_Y), .A(D4653_Y));
KC_XOR2_X3 D4558 ( .Y(D4558_Y), .B(D6128_Y), .A(D329_Y));
KC_XOR2_X3 D4557 ( .Y(D4557_Y), .B(D3049_Y), .A(D3036_Y));
KC_XOR2_X3 D4060 ( .Y(D4060_Y), .B(D4072_Y), .A(D4064_Y));
KC_XOR2_X3 D4057 ( .Y(D4057_Y), .B(D4072_Y), .A(D4062_Y));
KC_XOR2_X3 D4019 ( .Y(D4019_Y), .B(D4571_Y), .A(D1522_Y));
KC_XOR2_X3 D4018 ( .Y(D4018_Y), .B(D4571_Y), .A(D4022_Y));
KC_XOR2_X3 D3755 ( .Y(D3755_Y), .B(D4406_Y), .A(D3764_Y));
KC_XOR2_X3 D3754 ( .Y(D3754_Y), .B(D4406_Y), .A(D3756_Y));
KC_XOR2_X3 D1974 ( .Y(D1974_Y), .B(D8478_Y), .A(D1061_Y));
KC_XOR2_X3 D1797 ( .Y(D1797_Y), .B(D16696_Y), .A(D6563_Y));
KC_XOR2_X3 D1658 ( .Y(D1658_Y), .B(D5489_Y), .A(D5414_Y));
KC_XOR2_X3 D1519 ( .Y(D1519_Y), .B(D1506_Y), .A(D1418_Y));
KC_XOR2_X3 D1237 ( .Y(D1237_Y), .B(D8663_Y), .A(D1391_Y));
KC_XOR2_X3 D1160 ( .Y(D1160_Y), .B(D13094_Y), .A(D2357_Y));
KC_XOR2_X3 D1057 ( .Y(D1057_Y), .B(D8478_Y), .A(D1060_Y));
KC_XOR2_X3 D1056 ( .Y(D1056_Y), .B(D1076_Y), .A(D13620_Y));
KC_XOR2_X3 D829 ( .Y(D829_Y), .B(D16082_Y), .A(D10825_Y));
KC_XOR2_X3 D828 ( .Y(D828_Y), .B(D16082_Y), .A(D10822_Y));
KC_XOR2_X3 D706 ( .Y(D706_Y), .B(D16753_Y), .A(D6681_Y));
KC_XOR2_X3 D705 ( .Y(D705_Y), .B(D14586_Y), .A(D15250_Y));
KC_XOR2_X3 D356 ( .Y(D356_Y), .B(D6197_Y), .A(D1664_Y));
KC_OR4_X2 D16661 ( .Y(D16661_Y), .C(D16656_Y), .B(D16655_Y),     .D(D1400_Q), .A(D16672_Y));
KC_OR4_X2 D16612 ( .Y(D16612_Y), .C(D16551_Y), .B(D16604_Y),     .D(D1342_Y), .A(D1400_Q));
KC_OR4_X2 D16127 ( .Y(D16127_Y), .C(D16101_Y), .B(D16178_Y),     .D(D16085_Y), .A(D16101_Y));
KC_OR4_X2 D15568 ( .Y(D15568_Y), .C(D15530_Y), .B(D15567_Y),     .D(D15515_Y), .A(D15567_Y));
KC_OR4_X2 D13763 ( .Y(D13763_Y), .C(D13730_Y), .B(D13769_Y),     .D(D10266_Y), .A(D13725_Y));
KC_OR4_X2 D12653 ( .Y(D12653_Y), .C(D12621_Y), .B(D12133_Y),     .D(D13152_Y), .A(D12622_Y));
KC_OR4_X2 D12362 ( .Y(D12362_Y), .C(D823_Q), .B(D821_Q), .D(D12355_Q),     .A(D822_Q));
KC_OR4_X2 D12361 ( .Y(D12361_Y), .C(D12368_Q), .B(D12358_Q),     .D(D12359_Q), .A(D12274_Q));
KC_OR4_X2 D12354 ( .Y(D12354_Y), .C(D12352_Q), .B(D12349_Q),     .D(D12353_Q), .A(D12350_Q));
KC_OR4_X2 D12347 ( .Y(D12347_Y), .C(D12346_Q), .B(D12351_Q),     .D(D12342_Q), .A(D12367_Q));
KC_OR4_X2 D12345 ( .Y(D12345_Y), .C(D12416_Q), .B(D12343_Q),     .D(D2355_Q), .A(D12348_Q));
KC_OR4_X2 D12276 ( .Y(D12276_Y), .C(D12360_Q), .B(D12275_Q),     .D(D12356_Q), .A(D12357_Q));
KC_OR4_X2 D10050 ( .Y(D10050_Y), .C(D10035_Y), .B(D10084_Y),     .D(D2121_Y), .A(D10034_Y));
KC_OR4_X2 D9383 ( .Y(D9383_Y), .C(D9367_Y), .B(D9376_Y), .D(D9794_Y),     .A(D9370_Y));
KC_OR4_X2 D9357 ( .Y(D9357_Y), .C(D4526_Y), .B(D9355_Q), .D(D7523_Y),     .A(D9564_Y));
KC_OR4_X2 D9022 ( .Y(D9022_Y), .C(D9011_Y), .B(D9091_Y), .D(D9010_Y),     .A(D9009_Y));
KC_OR4_X2 D9020 ( .Y(D9020_Y), .C(D7528_Y), .B(D7525_Y), .D(D9004_Y),     .A(D9008_Y));
KC_OR4_X2 D8710 ( .Y(D8710_Y), .C(D8683_Y), .B(D8707_Y), .D(D8707_Y),     .A(D8707_Y));
KC_OR4_X2 D7895 ( .Y(D7895_Y), .C(D7453_Y), .B(D6457_Y), .D(D9104_Y),     .A(D1941_Q));
KC_OR4_X2 D7792 ( .Y(D7792_Y), .C(D7775_Y), .B(D9254_Y), .D(D9254_Y),     .A(D1825_Y));
KC_OR4_X2 D7390 ( .Y(D7390_Y), .C(D7267_Y), .B(D1910_Y), .D(D7189_Y),     .A(D7347_Y));
KC_OR4_X2 D6266 ( .Y(D6266_Y), .C(D6263_Y), .B(D6219_Y), .D(D14498_Y),     .A(D6238_Y));
KC_OR4_X2 D4554 ( .Y(D4554_Y), .C(D4496_Y), .B(D1611_Y), .D(D4523_Y),     .A(D1579_Y));
KC_OR4_X2 D1939 ( .Y(D1939_Y), .C(D5703_Y), .B(D1905_Y), .D(D7507_Y),     .A(D5826_Y));
KC_OR4_X2 D1653 ( .Y(D1653_Y), .C(D4091_Y), .B(D2716_Y), .D(D2716_Y),     .A(D4111_Y));
KC_OR4_X2 D1513 ( .Y(D1513_Y), .C(D1433_Y), .B(D2955_Y), .D(D2954_Y),     .A(D2903_Y));
KC_OR4_X2 D1049 ( .Y(D1049_Y), .C(D16359_Q), .B(D16361_Q),     .D(D16360_Q), .A(D2516_Q));
KC_OR4_X2 D606 ( .Y(D606_Y), .C(D13920_Q), .B(D607_Q), .D(D619_Q),     .A(D13201_Q));
KC_OR4_X2 D355 ( .Y(D355_Y), .C(D9163_Q), .B(D363_Q), .D(D9160_Q),     .A(D60_Q));
KC_INV_X2 D16382 ( .Y(D16382_Y), .A(D7609_Y));
KC_INV_X2 D15789 ( .Y(D15789_Y), .A(D14821_Y));
KC_INV_X2 D14785 ( .Y(D14785_Y), .A(D16559_Y));
KC_INV_X2 D14295 ( .Y(D14295_Y), .A(D1382_Q));
KC_INV_X2 D13858 ( .Y(D13858_Y), .A(D13846_Y));
KC_INV_X2 D13392 ( .Y(D13392_Y), .A(D14057_Y));
KC_INV_X2 D12678 ( .Y(D12678_Y), .A(D12661_Y));
KC_INV_X2 D11476 ( .Y(D11476_Y), .A(D10861_Y));
KC_INV_X2 D11276 ( .Y(D11276_Y), .A(D464_Y));
KC_INV_X2 D10803 ( .Y(D10803_Y), .A(D7974_Y));
KC_INV_X2 D10356 ( .Y(D10356_Y), .A(D10242_Y));
KC_INV_X2 D10292 ( .Y(D10292_Y), .A(D10304_Q));
KC_INV_X2 D10162 ( .Y(D10162_Y), .A(D724_Y));
KC_INV_X2 D10161 ( .Y(D10161_Y), .A(D12863_Y));
KC_INV_X2 D10160 ( .Y(D10160_Y), .A(D12763_Y));
KC_INV_X2 D10159 ( .Y(D10159_Y), .A(D13288_Y));
KC_INV_X2 D10158 ( .Y(D10158_Y), .A(D12761_Y));
KC_INV_X2 D10142 ( .Y(D10142_Y), .A(D13171_Y));
KC_INV_X2 D10057 ( .Y(D10057_Y), .A(D5828_Y));
KC_INV_X2 D10045 ( .Y(D10045_Y), .A(D7_Y));
KC_INV_X2 D9794 ( .Y(D9794_Y), .A(D9772_Y));
KC_INV_X2 D9616 ( .Y(D9616_Y), .A(D9634_Q));
KC_INV_X2 D9469 ( .Y(D9469_Y), .A(D9489_Y));
KC_INV_X2 D9380 ( .Y(D9380_Y), .A(D8307_Y));
KC_INV_X2 D9354 ( .Y(D9354_Y), .A(D12301_Y));
KC_INV_X2 D9269 ( .Y(D9269_Y), .A(D13289_Y));
KC_INV_X2 D9268 ( .Y(D9268_Y), .A(D13280_Q));
KC_INV_X2 D9147 ( .Y(D9147_Y), .A(D2099_Y));
KC_INV_X2 D9018 ( .Y(D9018_Y), .A(D7553_Y));
KC_INV_X2 D8950 ( .Y(D8950_Y), .A(D151_Q));
KC_INV_X2 D8817 ( .Y(D8817_Y), .A(D4130_Y));
KC_INV_X2 D8816 ( .Y(D8816_Y), .A(D8923_Y));
KC_INV_X2 D8707 ( .Y(D8707_Y), .A(D8682_Y));
KC_INV_X2 D8706 ( .Y(D8706_Y), .A(D289_Y));
KC_INV_X2 D8705 ( .Y(D8705_Y), .A(D8861_Y));
KC_INV_X2 D8550 ( .Y(D8550_Y), .A(D2032_Y));
KC_INV_X2 D8465 ( .Y(D8465_Y), .A(D545_Y));
KC_INV_X2 D8331 ( .Y(D8331_Y), .A(D6792_Y));
KC_INV_X2 D8239 ( .Y(D8239_Y), .A(D8090_Y));
KC_INV_X2 D8056 ( .Y(D8056_Y), .A(D5142_Q));
KC_INV_X2 D7785 ( .Y(D7785_Y), .A(D725_Y));
KC_INV_X2 D7731 ( .Y(D7731_Y), .A(D7691_Y));
KC_INV_X2 D7730 ( .Y(D7730_Y), .A(D723_Q));
KC_INV_X2 D7657 ( .Y(D7657_Y), .A(D7692_Y));
KC_INV_X2 D7585 ( .Y(D7585_Y), .A(D7558_Y));
KC_INV_X2 D7532 ( .Y(D7532_Y), .A(D70_Y));
KC_INV_X2 D7531 ( .Y(D7531_Y), .A(D6258_QN));
KC_INV_X2 D7472 ( .Y(D7472_Y), .A(D7471_Y));
KC_INV_X2 D7471 ( .Y(D7471_Y), .A(D431_Y));
KC_INV_X2 D7142 ( .Y(D7142_Y), .A(D7098_Y));
KC_INV_X2 D6478 ( .Y(D6478_Y), .A(D533_Q));
KC_INV_X2 D6477 ( .Y(D6477_Y), .A(D7940_Y));
KC_INV_X2 D6340 ( .Y(D6340_Y), .A(D6308_Y));
KC_INV_X2 D6339 ( .Y(D6339_Y), .A(D9263_Y));
KC_INV_X2 D6264 ( .Y(D6264_Y), .A(D7563_Y));
KC_INV_X2 D6263 ( .Y(D6263_Y), .A(D6185_Y));
KC_INV_X2 D6184 ( .Y(D6184_Y), .A(D6173_Y));
KC_INV_X2 D6183 ( .Y(D6183_Y), .A(D10159_Y));
KC_INV_X2 D6182 ( .Y(D6182_Y), .A(D6307_Y));
KC_INV_X2 D6181 ( .Y(D6181_Y), .A(D4628_Y));
KC_INV_X2 D6180 ( .Y(D6180_Y), .A(D5949_Y));
KC_INV_X2 D6179 ( .Y(D6179_Y), .A(D16754_Y));
KC_INV_X2 D6178 ( .Y(D6178_Y), .A(D6185_Y));
KC_INV_X2 D6118 ( .Y(D6118_Y), .A(D6264_Y));
KC_INV_X2 D5932 ( .Y(D5932_Y), .A(D6163_Y));
KC_INV_X2 D5805 ( .Y(D5805_Y), .A(D1614_Y));
KC_INV_X2 D5804 ( .Y(D5804_Y), .A(D7376_Y));
KC_INV_X2 D5682 ( .Y(D5682_Y), .A(D4395_Y));
KC_INV_X2 D5481 ( .Y(D5481_Y), .A(D5455_Y));
KC_INV_X2 D5480 ( .Y(D5480_Y), .A(D5377_Y));
KC_INV_X2 D5479 ( .Y(D5479_Y), .A(D5376_Y));
KC_INV_X2 D5404 ( .Y(D5404_Y), .A(D1636_Q));
KC_INV_X2 D4962 ( .Y(D4962_Y), .A(D3488_Y));
KC_INV_X2 D4961 ( .Y(D4961_Y), .A(D399_Y));
KC_INV_X2 D4814 ( .Y(D4814_Y), .A(D7581_Y));
KC_INV_X2 D4813 ( .Y(D4813_Y), .A(D7692_Y));
KC_INV_X2 D4812 ( .Y(D4812_Y), .A(D1825_Y));
KC_INV_X2 D4633 ( .Y(D4633_Y), .A(D4817_Q));
KC_INV_X2 D4482 ( .Y(D4482_Y), .A(D1661_Y));
KC_INV_X2 D4481 ( .Y(D4481_Y), .A(D10006_Q));
KC_INV_X2 D4391 ( .Y(D4391_Y), .A(D172_Y));
KC_INV_X2 D4390 ( .Y(D4390_Y), .A(D4393_Y));
KC_INV_X2 D4233 ( .Y(D4233_Y), .A(D7376_Y));
KC_INV_X2 D3881 ( .Y(D3881_Y), .A(D6794_Y));
KC_INV_X2 D3634 ( .Y(D3634_Y), .A(D5133_Q));
KC_INV_X2 D3633 ( .Y(D3633_Y), .A(D5114_Y));
KC_INV_X2 D3377 ( .Y(D3377_Y), .A(D3358_Y));
KC_INV_X2 D3276 ( .Y(D3276_Y), .A(D3278_Y));
KC_INV_X2 D3182 ( .Y(D3182_Y), .A(D4807_Y));
KC_INV_X2 D3181 ( .Y(D3181_Y), .A(D3161_Y));
KC_INV_X2 D3180 ( .Y(D3180_Y), .A(D4807_Y));
KC_INV_X2 D3073 ( .Y(D3073_Y), .A(D377_Y));
KC_INV_X2 D3072 ( .Y(D3072_Y), .A(D38_Y));
KC_INV_X2 D3071 ( .Y(D3071_Y), .A(D321_Y));
KC_INV_X2 D2997 ( .Y(D2997_Y), .A(D2897_Y));
KC_INV_X2 D2996 ( .Y(D2996_Y), .A(D2846_Y));
KC_INV_X2 D2880 ( .Y(D2880_Y), .A(D2835_Y));
KC_INV_X2 D2353 ( .Y(D2353_Y), .A(D7669_Y));
KC_INV_X2 D2223 ( .Y(D2223_Y), .A(D8454_Y));
KC_INV_X2 D2162 ( .Y(D2162_Y), .A(D5828_Y));
KC_INV_X2 D1937 ( .Y(D1937_Y), .A(D101_Y));
KC_INV_X2 D1936 ( .Y(D1936_Y), .A(D7974_Y));
KC_INV_X2 D1935 ( .Y(D1935_Y), .A(D7549_Y));
KC_INV_X2 D1648 ( .Y(D1648_Y), .A(D6408_Y));
KC_INV_X2 D1506 ( .Y(D1506_Y), .A(D16754_Y));
KC_INV_X2 D1505 ( .Y(D1505_Y), .A(D3510_Y));
KC_INV_X2 D1504 ( .Y(D1504_Y), .A(D3773_Y));
KC_INV_X2 D1143 ( .Y(D1143_Y), .A(D6791_Y));
KC_INV_X2 D481 ( .Y(D481_Y), .A(D12764_Y));
KC_INV_X2 D447 ( .Y(D447_Y), .A(D7723_Y));
KC_INV_X2 D417 ( .Y(D417_Y), .A(D6075_Y));
KC_INV_X2 D383 ( .Y(D383_Y), .A(D7636_Y));
KC_INV_X2 D382 ( .Y(D382_Y), .A(D6075_Y));
KC_INV_X2 D352 ( .Y(D352_Y), .A(D1008_Y));
KC_AO21_X3 D332 ( .B(D1767_Y), .A1(D6198_Y), .Y(D332_Y), .A0(D6157_Y));
KC_SDFFRNHQ_X1 D16718 ( .Q(D16718_Q), .SI(D16734_Y), .SE(D16719_Y),     .D(D16718_Q), .RN(D16610_Y), .CK(D16716_Y));
KC_SDFFRNHQ_X1 D16717 ( .Q(D16717_Q), .SI(D16733_Y), .SE(D16719_Y),     .D(D16717_Q), .RN(D16610_Y), .CK(D2693_Y));
KC_SDFFRNHQ_X1 D16710 ( .Q(D16710_Q), .SI(D16736_Y), .SE(D16712_Y),     .D(D16710_Q), .RN(D16610_Y), .CK(D16705_Y));
KC_SDFFRNHQ_X1 D16635 ( .Q(D16635_Q), .SI(D16396_Y), .SE(D16645_Y),     .D(D16635_Q), .RN(D16610_Y), .CK(D2689_Y));
KC_SDFFRNHQ_X1 D16634 ( .Q(D16634_Q), .SI(D16394_Y), .SE(D16645_Y),     .D(D16634_Q), .RN(D16610_Y), .CK(D16629_Y));
KC_SDFFRNHQ_X1 D16566 ( .Q(D16566_Q), .SI(D16397_Y), .SE(D16568_Y),     .D(D16566_Q), .RN(D16579_Y), .CK(D2688_Y));
KC_SDFFRNHQ_X1 D16565 ( .Q(D16565_Q), .SI(D16395_Y), .SE(D16568_Y),     .D(D16565_Q), .RN(D16579_Y), .CK(D16567_Y));
KC_SDFFRNHQ_X1 D16332 ( .Q(D16332_Q), .SI(D16328_Y), .SE(D16337_Y),     .D(D16332_Q), .RN(D16267_Y), .CK(D16294_Y));
KC_SDFFRNHQ_X1 D16331 ( .Q(D16331_Q), .SI(D16320_Y), .SE(D16345_Y),     .D(D16331_Q), .RN(D16267_Y), .CK(D16321_Y));
KC_SDFFRNHQ_X1 D15153 ( .Q(D15153_Q), .SI(D15139_Y), .SE(D15158_Y),     .D(D15153_Q), .RN(D14291_Y), .CK(D15144_Y));
KC_SDFFRNHQ_X1 D15152 ( .Q(D15152_Q), .SI(D15138_Y), .SE(D15158_Y),     .D(D15152_Q), .RN(D14291_Y), .CK(D15143_Y));
KC_SDFFRNHQ_X1 D14702 ( .Q(D14702_Q), .SI(D14692_Y), .SE(D14713_Y),     .D(D14702_Q), .RN(D13265_Y), .CK(D14693_Y));
KC_SDFFRNHQ_X1 D14701 ( .Q(D14701_Q), .SI(D14690_Y), .SE(D14713_Y),     .D(D14701_Q), .RN(D13265_Y), .CK(D14691_Y));
KC_SDFFRNHQ_X1 D13837 ( .Q(D13837_Q), .SI(D13766_Y), .SE(D13842_Y),     .D(D13837_Q), .RN(D13757_Y), .CK(D13841_Y));
KC_SDFFRNHQ_X1 D13836 ( .Q(D13836_Q), .SI(D13767_Y), .SE(D13839_Y),     .D(D13836_Q), .RN(D13757_Y), .CK(D13840_Y));
KC_SDFFRNHQ_X1 D12366 ( .Q(D12366_Q), .SI(D12363_Y), .SE(D12369_Y),     .D(D12366_Q), .RN(D12838_Y), .CK(D12364_Y));
KC_SDFFRNHQ_X1 D12291 ( .Q(D12291_Q), .SI(D12286_Y), .SE(D12303_Y),     .D(D12291_Q), .RN(D12734_Y), .CK(D12281_Y));
KC_SDFFRNHQ_X1 D11606 ( .Q(D11606_Q), .SI(D11540_Y), .SE(D11609_Y),     .D(D11606_Q), .RN(D13757_Y), .CK(D11601_Y));
KC_SDFFRNHQ_X1 D11413 ( .Q(D11413_Q), .SI(D11410_Y), .SE(D11416_Y),     .D(D11413_Q), .RN(D12898_Y), .CK(D11411_Y));
KC_SDFFRNHQ_X1 D11051 ( .Q(D11051_Q), .SI(D11045_Y), .SE(D11057_Y),     .D(D11051_Q), .RN(D1934_Y), .CK(D11044_Y));
KC_SDFFRNHQ_X1 D11050 ( .Q(D11050_Q), .SI(D11039_Y), .SE(D11057_Y),     .D(D11050_Q), .RN(D1934_Y), .CK(D11043_Y));
KC_SDFFRNHQ_X1 D10828 ( .Q(D10828_Q), .SI(D829_Y), .SE(D10830_Y),     .D(D10828_Q), .RN(D10726_Y), .CK(D10815_Y));
KC_SDFFRNHQ_X1 D10826 ( .Q(D10826_Q), .SI(D828_Y), .SE(D10830_Y),     .D(D10826_Q), .RN(D10726_Y), .CK(D10811_Y));
KC_SDFFRNHQ_X1 D9918 ( .Q(D9918_Q), .SI(D1237_Y), .SE(D9921_Y),     .D(D9918_Q), .RN(D1934_Y), .CK(D1388_Y));
KC_SDFFRNHQ_X1 D8605 ( .Q(D8605_Q), .SI(D8596_Y), .SE(D8606_Y),     .D(D8605_Q), .RN(D1934_Y), .CK(D8597_Y));
KC_SDFFRNHQ_X1 D8159 ( .Q(D8159_Q), .SI(D8164_Y), .SE(D8166_Y),     .D(D8159_Q), .RN(D8300_Y), .CK(D8155_Y));
KC_SDFFRNHQ_X1 D8158 ( .Q(D8158_Q), .SI(D706_Y), .SE(D8166_Y),     .D(D8158_Q), .RN(D8300_Y), .CK(D8154_Y));
KC_SDFFRNHQ_X1 D6616 ( .Q(D6616_Q), .SI(D1797_Y), .SE(D6617_Y),     .D(D6616_Q), .RN(D9375_Y), .CK(D1799_Y));
KC_SDFFRNHQ_X1 D6402 ( .Q(D6402_Q), .SI(D6391_Y), .SE(D6414_Y),     .D(D6402_Q), .RN(D7786_Y), .CK(D6389_Y));
KC_SDFFRNHQ_X1 D6401 ( .Q(D6401_Q), .SI(D6392_Y), .SE(D6414_Y),     .D(D6401_Q), .RN(D7786_Y), .CK(D6390_Y));
KC_SDFFRNHQ_X1 D5815 ( .Q(D5815_Q), .SI(D5806_Y), .SE(D5823_Y),     .D(D5815_Q), .RN(D13757_Y), .CK(D5807_Y));
KC_SDFFRNHQ_X1 D5814 ( .Q(D5814_Q), .SI(D5707_Y), .SE(D5823_Y),     .D(D5814_Q), .RN(D13757_Y), .CK(D5808_Y));
KC_SDFFRNHQ_X1 D5416 ( .Q(D5416_Q), .SI(D1658_Y), .SE(D5419_Y),     .D(D5416_Q), .RN(D8300_Y), .CK(D5410_Y));
KC_SDFFRNHQ_X1 D5415 ( .Q(D5415_Q), .SI(D5485_Y), .SE(D1676_Y),     .D(D5415_Q), .RN(D8300_Y), .CK(D5411_Y));
KC_SDFFRNHQ_X1 D4647 ( .Q(D4647_Q), .SI(D4645_Y), .SE(D4652_Y),     .D(D4647_Q), .RN(D13757_Y), .CK(D4642_Y));
KC_SDFFRNHQ_X1 D4066 ( .Q(D4066_Q), .SI(D4060_Y), .SE(D4071_Y),     .D(D4066_Q), .RN(D1934_Y), .CK(D4061_Y));
KC_SDFFRNHQ_X1 D4065 ( .Q(D4065_Q), .SI(D4057_Y), .SE(D4071_Y),     .D(D4065_Q), .RN(D1934_Y), .CK(D4059_Y));
KC_SDFFRNHQ_X1 D4024 ( .Q(D4024_Q), .SI(D4018_Y), .SE(D4030_Y),     .D(D4024_Q), .RN(D1934_Y), .CK(D3983_Y));
KC_SDFFRNHQ_X1 D4023 ( .Q(D4023_Q), .SI(D4019_Y), .SE(D4030_Y),     .D(D4023_Q), .RN(D1934_Y), .CK(D1520_Y));
KC_SDFFRNHQ_X1 D3758 ( .Q(D3758_Q), .SI(D3755_Y), .SE(D3763_Y),     .D(D3758_Q), .RN(D3542_Y), .CK(D708_Y));
KC_SDFFRNHQ_X1 D3757 ( .Q(D3757_Q), .SI(D3754_Y), .SE(D3763_Y),     .D(D3757_Q), .RN(D3542_Y), .CK(D5248_Y));
KC_SDFFRNHQ_X1 D1806 ( .Q(D1806_Q), .SI(D6556_Y), .SE(D6617_Y),     .D(D1806_Q), .RN(D9375_Y), .CK(D1800_Y));
KC_SDFFRNHQ_X1 D1394 ( .Q(D1394_Q), .SI(D9849_Y), .SE(D9921_Y),     .D(D1394_Q), .RN(D1934_Y), .CK(D8661_Y));
KC_SDFFRNHQ_X1 D1393 ( .Q(D1393_Q), .SI(D12049_Y), .SE(D11609_Y),     .D(D1393_Q), .RN(D13757_Y), .CK(D11602_Y));
KC_SDFFRNHQ_X1 D1392 ( .Q(D1392_Q), .SI(D16735_Y), .SE(D16713_Y),     .D(D1392_Q), .RN(D16610_Y), .CK(D2692_Y));
KC_SDFFRNHQ_X1 D1243 ( .Q(D1243_Q), .SI(D8602_Y), .SE(D8606_Y),     .D(D1243_Q), .RN(D1934_Y), .CK(D8601_Y));
KC_SDFFRNHQ_X1 D1242 ( .Q(D1242_Q), .SI(D12547_Y), .SE(D2403_Y),     .D(D1242_Q), .RN(D13757_Y), .CK(D13091_Y));
KC_SDFFRNHQ_X1 D1162 ( .Q(D1162_Q), .SI(D1160_Y), .SE(D2403_Y),     .D(D1162_Q), .RN(D13757_Y), .CK(D13052_Y));
KC_SDFFRNHQ_X1 D1064 ( .Q(D1064_Q), .SI(D11409_Y), .SE(D11416_Y),     .D(D1064_Q), .RN(D12898_Y), .CK(D2263_Y));
KC_SDFFRNHQ_X1 D1063 ( .Q(D1063_Q), .SI(D13616_Y), .SE(D13639_Y),     .D(D1063_Q), .RN(D13757_Y), .CK(D1055_Y));
KC_SDFFRNHQ_X1 D1062 ( .Q(D1062_Q), .SI(D1056_Y), .SE(D13639_Y),     .D(D1062_Q), .RN(D13757_Y), .CK(D12998_Y));
KC_SDFFRNHQ_X1 D944 ( .Q(D944_Q), .SI(D1057_Y), .SE(D9722_Y),     .D(D944_Q), .RN(D8300_Y), .CK(D9626_Y));
KC_SDFFRNHQ_X1 D943 ( .Q(D943_Q), .SI(D1974_Y), .SE(D9722_Y),     .D(D943_Q), .RN(D8300_Y), .CK(D1946_Y));
KC_SDFFRNHQ_X1 D361 ( .Q(D361_Q), .SI(D356_Y), .SE(D6207_Y),     .D(D361_Q), .RN(D13757_Y), .CK(D6206_Y));
KC_SDFFRNHQ_X1 D331 ( .Q(D331_Q), .SI(D4558_Y), .SE(D33_Y), .D(D331_Q),     .RN(D1652_Y), .CK(D6122_Y));
KC_SDFFRNHQ_X1 D330 ( .Q(D330_Q), .SI(D6123_Y), .SE(D33_Y), .D(D330_Q),     .RN(D1652_Y), .CK(D6120_Y));
KC_MX2_X2 D16730 ( .Y(D16730_Y), .A(D16727_Y), .B(D16725_Y),     .S0(D16715_Y));
KC_MX2_X2 D16729 ( .Y(D16729_Y), .A(D2696_Y), .B(D16725_Y),     .S0(D16715_Y));
KC_MX2_X2 D16709 ( .Y(D16709_Y), .A(D16706_Y), .B(D16714_Y),     .S0(D16772_Y));
KC_MX2_X2 D16708 ( .Y(D16708_Y), .A(D1387_Y), .B(D16714_Y),     .S0(D16772_Y));
KC_MX2_X2 D16633 ( .Y(D16633_Y), .A(D16631_Y), .B(D16644_Y),     .S0(D16639_Y));
KC_MX2_X2 D16617 ( .Y(D16617_Y), .A(D16616_Y), .B(D16644_Y),     .S0(D16639_Y));
KC_MX2_X2 D16591 ( .Y(D16591_Y), .A(D16552_Y), .B(D16589_Y),     .S0(D16588_Y));
KC_MX2_X2 D16583 ( .Y(D16583_Y), .A(D1404_Y), .B(D16589_Y),     .S0(D16588_Y));
KC_MX2_X2 D16330 ( .Y(D16330_Y), .A(D16324_Y), .B(D16342_Y),     .S0(D16341_Y));
KC_MX2_X2 D16329 ( .Y(D16329_Y), .A(D16322_Y), .B(D16342_Y),     .S0(D16341_Y));
KC_MX2_X2 D15151 ( .Y(D15151_Y), .A(D15140_Y), .B(D15157_Y),     .S0(D15159_Y));
KC_MX2_X2 D15150 ( .Y(D15150_Y), .A(D15141_Y), .B(D15157_Y),     .S0(D15159_Y));
KC_MX2_X2 D14700 ( .Y(D14700_Y), .A(D14695_Y), .B(D14804_Y),     .S0(D14712_Y));
KC_MX2_X2 D14699 ( .Y(D14699_Y), .A(D14696_Y), .B(D14804_Y),     .S0(D14712_Y));
KC_MX2_X2 D13835 ( .Y(D13835_Y), .A(D13828_Y), .B(D13844_Y),     .S0(D13843_Y));
KC_MX2_X2 D13834 ( .Y(D13834_Y), .A(D13829_Y), .B(D13844_Y),     .S0(D13843_Y));
KC_MX2_X2 D13621 ( .Y(D13621_Y), .A(D13611_Y), .B(D13009_Y),     .S0(D1076_Y));
KC_MX2_X2 D13620 ( .Y(D13620_Y), .A(D13614_Y), .B(D13009_Y),     .S0(D1076_Y));
KC_MX2_X2 D12290 ( .Y(D12290_Y), .A(D12285_Y), .B(D12308_Y),     .S0(D12304_Y));
KC_MX2_X2 D12289 ( .Y(D12289_Y), .A(D12283_Y), .B(D12308_Y),     .S0(D12304_Y));
KC_MX2_X2 D11669 ( .Y(D11669_Y), .A(D12201_Y), .B(D11649_Y),     .S0(D10181_Y));
KC_MX2_X2 D11635 ( .Y(D11635_Y), .A(D11628_Y), .B(D11183_Y),     .S0(D12183_Y));
KC_MX2_X2 D11605 ( .Y(D11605_Y), .A(D11604_Y), .B(D11611_Y),     .S0(D11612_Y));
KC_MX2_X2 D11412 ( .Y(D11412_Y), .A(D11408_Y), .B(D11418_Y),     .S0(D11417_Y));
KC_MX2_X2 D11049 ( .Y(D11049_Y), .A(D11046_Y), .B(D11054_Y),     .S0(D11055_Y));
KC_MX2_X2 D11048 ( .Y(D11048_Y), .A(D11042_Y), .B(D11054_Y),     .S0(D11055_Y));
KC_MX2_X2 D10825 ( .Y(D10825_Y), .A(D10817_Y), .B(D10829_Y),     .S0(D16082_Y));
KC_MX2_X2 D10822 ( .Y(D10822_Y), .A(D10813_Y), .B(D10829_Y),     .S0(D16082_Y));
KC_MX2_X2 D9917 ( .Y(D9917_Y), .A(D9915_Y), .B(D8662_Y), .S0(D8663_Y));
KC_MX2_X2 D8722 ( .Y(D8722_Y), .A(D8732_Y), .B(D8665_Y), .S0(D8806_Y));
KC_MX2_X2 D8604 ( .Y(D8604_Y), .A(D7016_Y), .B(D8608_Y), .S0(D8607_Y));
KC_MX2_X2 D8603 ( .Y(D8603_Y), .A(D8598_Y), .B(D8608_Y), .S0(D8607_Y));
KC_MX2_X2 D7610 ( .Y(D7610_Y), .A(D7569_Y), .B(D7544_Y), .S0(D7572_Y));
KC_MX2_X2 D6681 ( .Y(D6681_Y), .A(D6676_Y), .B(D8165_Y),     .S0(D16753_Y));
KC_MX2_X2 D6563 ( .Y(D6563_Y), .A(D6557_Y), .B(D6567_Y),     .S0(D16696_Y));
KC_MX2_X2 D6562 ( .Y(D6562_Y), .A(D1798_Y), .B(D6567_Y),     .S0(D16696_Y));
KC_MX2_X2 D6400 ( .Y(D6400_Y), .A(D6397_Y), .B(D6413_Y),     .S0(D14591_Y));
KC_MX2_X2 D6399 ( .Y(D6399_Y), .A(D6394_Y), .B(D6413_Y),     .S0(D14591_Y));
KC_MX2_X2 D6349 ( .Y(D6349_Y), .A(D6339_Y), .B(D6339_Y), .S0(D6341_Y));
KC_MX2_X2 D6125 ( .Y(D6125_Y), .A(D6124_Y), .B(D30_Y), .S0(D6128_Y));
KC_MX2_X2 D5813 ( .Y(D5813_Y), .A(D5810_Y), .B(D5822_Y), .S0(D6275_Y));
KC_MX2_X2 D5699 ( .Y(D5699_Y), .A(D5694_Y), .B(D5822_Y), .S0(D6275_Y));
KC_MX2_X2 D5488 ( .Y(D5488_Y), .A(D5482_Y), .B(D5490_Y), .S0(D5489_Y));
KC_MX2_X2 D5414 ( .Y(D5414_Y), .A(D1659_Y), .B(D5490_Y), .S0(D5489_Y));
KC_MX2_X2 D4653 ( .Y(D4653_Y), .A(D4644_Y), .B(D1818_Y), .S0(D6197_Y));
KC_MX2_X2 D4064 ( .Y(D4064_Y), .A(D4058_Y), .B(D4073_Y), .S0(D4072_Y));
KC_MX2_X2 D4063 ( .Y(D4063_Y), .A(D4078_Y), .B(D4036_Y), .S0(D4076_Y));
KC_MX2_X2 D4062 ( .Y(D4062_Y), .A(D4054_Y), .B(D4073_Y), .S0(D4072_Y));
KC_MX2_X2 D4022 ( .Y(D4022_Y), .A(D4020_Y), .B(D1535_Y), .S0(D4571_Y));
KC_MX2_X2 D3756 ( .Y(D3756_Y), .A(D3753_Y), .B(D5253_Y), .S0(D4406_Y));
KC_MX2_X2 D3390 ( .Y(D3390_Y), .A(D3353_Y), .B(D3352_Y), .S0(D3337_Y));
KC_MX2_X2 D2893 ( .Y(D2893_Y), .A(D4310_Y), .B(D4366_Y), .S0(D2873_Y));
KC_MX2_X2 D2357 ( .Y(D2357_Y), .A(D2359_Y), .B(D13093_Y),     .S0(D13094_Y));
KC_MX2_X2 D2100 ( .Y(D2100_Y), .A(D2061_Y), .B(D9672_Y), .S0(D9495_Y));
KC_MX2_X2 D1664 ( .Y(D1664_Y), .A(D1657_Y), .B(D1818_Y), .S0(D6197_Y));
KC_MX2_X2 D1522 ( .Y(D1522_Y), .A(D3981_Y), .B(D1535_Y), .S0(D4571_Y));
KC_MX2_X2 D1391 ( .Y(D1391_Y), .A(D8659_Y), .B(D8662_Y), .S0(D8663_Y));
KC_MX2_X2 D1390 ( .Y(D1390_Y), .A(D11600_Y), .B(D11611_Y),     .S0(D11612_Y));
KC_MX2_X2 D1241 ( .Y(D1241_Y), .A(D12549_Y), .B(D13093_Y),     .S0(D13094_Y));
KC_MX2_X2 D1061 ( .Y(D1061_Y), .A(D9719_Y), .B(D9721_Y), .S0(D8478_Y));
KC_MX2_X2 D1060 ( .Y(D1060_Y), .A(D8467_Y), .B(D9721_Y), .S0(D8478_Y));
KC_MX2_X2 D710 ( .Y(D710_Y), .A(D6678_Y), .B(D8165_Y), .S0(D16753_Y));
KC_MX2_X2 D612 ( .Y(D612_Y), .A(D11646_Y), .B(D11653_Y),     .S0(D11653_Y));
KC_MX2_X2 D454 ( .Y(D454_Y), .A(D4940_Y), .B(D6370_Y), .S0(D4917_Y));
KC_MX2_X2 D329 ( .Y(D329_Y), .A(D156_Y), .B(D30_Y), .S0(D6128_Y));
KC_BUF_X6 D16614 ( .Y(D16614_Y), .A(D16639_Y));
KC_BUF_X6 D16610 ( .Y(D16610_Y), .A(D14858_Y));
KC_BUF_X6 D16594 ( .Y(D16594_Y), .A(D16588_Y));
KC_BUF_X6 D16579 ( .Y(D16579_Y), .A(D14858_Y));
KC_BUF_X6 D16469 ( .Y(D16469_Y), .A(D16474_Q));
KC_BUF_X6 D16384 ( .Y(D16384_Y), .A(D965_Y));
KC_BUF_X6 D16383 ( .Y(D16383_Y), .A(D965_Y));
KC_BUF_X6 D16352 ( .Y(D16352_Y), .A(D965_Y));
KC_BUF_X6 D15990 ( .Y(D15990_Y), .A(D16383_Y));
KC_BUF_X6 D15790 ( .Y(D15790_Y), .A(D14858_Y));
KC_BUF_X6 D14869 ( .Y(D14869_Y), .A(D14858_Y));
KC_BUF_X6 D14786 ( .Y(D14786_Y), .A(D14796_Y));
KC_BUF_X6 D14489 ( .Y(D14489_Y), .A(D14858_Y));
KC_BUF_X6 D14474 ( .Y(D14474_Y), .A(D14858_Y));
KC_BUF_X6 D14296 ( .Y(D14296_Y), .A(D14858_Y));
KC_BUF_X6 D14163 ( .Y(D14163_Y), .A(D2510_Y));
KC_BUF_X6 D13859 ( .Y(D13859_Y), .A(D13859_A));
KC_BUF_X6 D13825 ( .Y(D13825_Y), .A(D14858_Y));
KC_BUF_X6 D13758 ( .Y(D13758_Y), .A(D14858_Y));
KC_BUF_X6 D13394 ( .Y(D13394_Y), .A(D12697_Y));
KC_BUF_X6 D13266 ( .Y(D13266_Y), .A(D13242_Y));
KC_BUF_X6 D13265 ( .Y(D13265_Y), .A(D12280_Y));
KC_BUF_X6 D13194 ( .Y(D13194_Y), .A(D12280_Y));
KC_BUF_X6 D13171 ( .Y(D13171_Y), .A(D2469_Q));
KC_BUF_X6 D12846 ( .Y(D12846_Y), .A(D12280_Y));
KC_BUF_X6 D12679 ( .Y(D12679_Y), .A(D12280_Y));
KC_BUF_X6 D12339 ( .Y(D12339_Y), .A(D10725_Y));
KC_BUF_X6 D11990 ( .Y(D11990_Y), .A(D9555_Y));
KC_BUF_X6 D10726 ( .Y(D10726_Y), .A(D12280_Y));
KC_BUF_X6 D10725 ( .Y(D10725_Y), .A(D12280_Y));
KC_BUF_X6 D10358 ( .Y(D10358_Y), .A(D7757_Y));
KC_BUF_X6 D10357 ( .Y(D10357_Y), .A(D9538_Y));
KC_BUF_X6 D10143 ( .Y(D10143_Y), .A(D10146_Q));
KC_BUF_X6 D9617 ( .Y(D9617_Y), .A(D7756_Y));
KC_BUF_X6 D9381 ( .Y(D9381_Y), .A(D10726_Y));
KC_BUF_X6 D9271 ( .Y(D9271_Y), .A(D9358_Y));
KC_BUF_X6 D9214 ( .Y(D9214_Y), .A(D9358_Y));
KC_BUF_X6 D8894 ( .Y(D8894_Y), .A(D9358_Y));
KC_BUF_X6 D8818 ( .Y(D8818_Y), .A(D9358_Y));
KC_BUF_X6 D8466 ( .Y(D8466_Y), .A(D7991_Y));
KC_BUF_X6 D8336 ( .Y(D8336_Y), .A(D7824_Y));
KC_BUF_X6 D8240 ( .Y(D8240_Y), .A(D7990_Y));
KC_BUF_X6 D7893 ( .Y(D7893_Y), .A(D7795_Y));
KC_BUF_X6 D7892 ( .Y(D7892_Y), .A(D7893_Y));
KC_BUF_X6 D7788 ( .Y(D7788_Y), .A(D7795_Y));
KC_BUF_X6 D7786 ( .Y(D7786_Y), .A(D7795_Y));
KC_BUF_X6 D6759 ( .Y(D6759_Y), .A(D8177_Y));
KC_BUF_X6 D6342 ( .Y(D6342_Y), .A(D3225_Y));
KC_BUF_X6 D5683 ( .Y(D5683_Y), .A(D7795_Y));
KC_BUF_X6 D4634 ( .Y(D4634_Y), .A(D7795_Y));
KC_BUF_X6 D4553 ( .Y(D4553_Y), .A(D1934_Y));
KC_BUF_X6 D4483 ( .Y(D4483_Y), .A(D9358_Y));
KC_BUF_X6 D3577 ( .Y(D3577_Y), .A(D7795_Y));
KC_BUF_X6 D2882 ( .Y(D2882_Y), .A(D4483_Y));
KC_BUF_X6 D2677 ( .Y(D2677_Y), .A(D2627_Y));
KC_BUF_X6 D2676 ( .Y(D2676_Y), .A(D15700_Y));
KC_BUF_X6 D1652 ( .Y(D1652_Y), .A(D7795_Y));
KC_BUF_X6 D813 ( .Y(D813_Y), .A(D1976_Y));
KC_BUF_X6 D324 ( .Y(D324_Y), .A(D9358_Y));
KC_AOI22_X5 D488 ( .A1(D3516_Y), .B0(D5037_Y), .B1(D4913_Y),     .Y(D488_Y), .A0(D3446_Y));
KC_AOI22_X5 D461 ( .A1(D10142_Y), .B0(D1862_Y), .B1(D7819_Y),     .Y(D461_Y), .A0(D9237_Y));
KC_AOI22_X5 D460 ( .A1(D399_Y), .B0(D4914_Y), .B1(D3480_Y), .Y(D460_Y),     .A0(D3467_Y));
KC_AOI22_X5 D459 ( .A1(D7759_Y), .B0(D7779_Y), .B1(D12863_Y),     .Y(D459_Y), .A0(D9237_Y));
KC_AOI22_X5 D458 ( .A1(D9354_Y), .B0(D1862_Y), .B1(D7822_Y),     .Y(D458_Y), .A0(D9237_Y));
KC_AOI22_X5 D333 ( .A1(D7495_Y), .B0(D7361_Y), .B1(D8849_Y),     .Y(D333_Y), .A0(D9052_Y));
KC_AOI22_X5 D306 ( .A1(D318_Y), .B0(D6046_Y), .B1(D5936_Y), .Y(D306_Y),     .A0(D6043_Y));
KC_NOR2B_X2 D10117 ( .B(D10057_Y), .Y(D10117_Y), .AN(D10049_Q));
KC_NOR2B_X2 D2525 ( .B(D2330_Y), .Y(D2525_Y), .AN(D2408_Y));
KC_NOR2B_X2 D16 ( .B(D8952_Q), .Y(D16_Y), .AN(D149_Q));
KC_ADDF_X3 D16760 ( .Ci(D10864_Y), .B(D10863_Y), .Co(D16760_Co),     .A(D10870_Y));
KC_ADDF_X3 D16759 ( .Ci(D10220_Q), .B(D10221_Q), .Co(D16759_Co),     .A(D10223_Q));
KC_ADDF_X3 D16758 ( .Ci(D10219_Q), .B(D10217_Q), .Co(D16758_Co),     .A(D698_Q));
KC_ADDF_X3 D10240 ( .Ci(D10227_Q), .B(D10231_Q), .Co(D10240_Co),     .A(D10228_Q));
KC_ADDF_X3 D9230 ( .Ci(D9226_Y), .B(D9297_Y), .Co(D9230_Co),     .A(D7780_Y));
KC_ADDF_X3 D16756 ( .Ci(D8666_Y), .B(D8666_Y), .Co(D16756_Co),     .A(D8665_Y));
KC_ADDF_X3 D6208 ( .Ci(D6149_Y), .B(D1805_Y), .Co(D6208_Co),     .A(D6161_Y));
KC_ADDF_X3 D583 ( .Ci(D7381_Y), .B(D7381_Y), .Co(D583_Co),     .A(D7331_Y));
KC_ADDF_X3 D3598 ( .Ci(D3476_Y), .B(D3407_Y), .Co(D3598_Co),     .A(D3564_Y));
KC_ADDF_X3 D335 ( .Ci(D7531_Y), .B(D7515_Y), .Co(D335_Co),     .A(D7515_Y));
KC_ADDF_X3 D274 ( .Ci(D4394_Y), .B(D4390_Y), .Co(D274_Co),     .A(D4391_Y));
KC_TIELO_X1 D16725 ( .Y(D16725_Y));
KC_TIELO_X1 D16719 ( .Y(D16719_Y));
KC_TIELO_X1 D16714 ( .Y(D16714_Y));
KC_TIELO_X1 D16713 ( .Y(D16713_Y));
KC_TIELO_X1 D16712 ( .Y(D16712_Y));
KC_TIELO_X1 D16645 ( .Y(D16645_Y));
KC_TIELO_X1 D16644 ( .Y(D16644_Y));
KC_TIELO_X1 D16592 ( .Y(D16592_Y));
KC_TIELO_X1 D16589 ( .Y(D16589_Y));
KC_TIELO_X1 D16568 ( .Y(D16568_Y));
KC_TIELO_X1 D16525 ( .Y(D16525_Y));
KC_TIELO_X1 D16479 ( .Y(D16479_Y));
KC_TIELO_X1 D16345 ( .Y(D16345_Y));
KC_TIELO_X1 D16342 ( .Y(D16342_Y));
KC_TIELO_X1 D16337 ( .Y(D16337_Y));
KC_TIELO_X1 D16336 ( .Y(D16336_Y));
KC_TIELO_X1 D16298 ( .Y(D16298_Y));
KC_TIELO_X1 D15158 ( .Y(D15158_Y));
KC_TIELO_X1 D15157 ( .Y(D15157_Y));
KC_TIELO_X1 D14804 ( .Y(D14804_Y));
KC_TIELO_X1 D14713 ( .Y(D14713_Y));
KC_TIELO_X1 D16768 ( .Y(D16768_Y));
KC_TIELO_X1 D16766 ( .Y(D16766_Y));
KC_TIELO_X1 D14197 ( .Y(D14197_Y));
KC_TIELO_X1 D14110 ( .Y(D14110_Y));
KC_TIELO_X1 D14006 ( .Y(D14006_Y));
KC_TIELO_X1 D13867 ( .Y(D13867_Y));
KC_TIELO_X1 D13844 ( .Y(D13844_Y));
KC_TIELO_X1 D13842 ( .Y(D13842_Y));
KC_TIELO_X1 D13839 ( .Y(D13839_Y));
KC_TIELO_X1 D13639 ( .Y(D13639_Y));
KC_TIELO_X1 D13408 ( .Y(D13408_Y));
KC_TIELO_X1 D13290 ( .Y(D13290_Y));
KC_TIELO_X1 D13286 ( .Y(D13286_Y));
KC_TIELO_X1 D13215 ( .Y(D13215_Y));
KC_TIELO_X1 D13093 ( .Y(D13093_Y));
KC_TIELO_X1 D13009 ( .Y(D13009_Y));
KC_TIELO_X1 D12867 ( .Y(D12867_Y));
KC_TIELO_X1 D12758 ( .Y(D12758_Y));
KC_TIELO_X1 D12691 ( .Y(D12691_Y));
KC_TIELO_X1 D12369 ( .Y(D12369_Y));
KC_TIELO_X1 D12308 ( .Y(D12308_Y));
KC_TIELO_X1 D12303 ( .Y(D12303_Y));
KC_TIELO_X1 D12240 ( .Y(D12240_Y));
KC_TIELO_X1 D12183 ( .Y(D12183_Y));
KC_TIELO_X1 D12129 ( .Y(D12129_Y));
KC_TIELO_X1 D12128 ( .Y(D12128_Y));
KC_TIELO_X1 D11996 ( .Y(D11996_Y));
KC_TIELO_X1 D11933 ( .Y(D11933_Y));
KC_TIELO_X1 D11932 ( .Y(D11932_Y));
KC_TIELO_X1 D11931 ( .Y(D11931_Y));
KC_TIELO_X1 D11676 ( .Y(D11676_Y));
KC_TIELO_X1 D11613 ( .Y(D11613_Y));
KC_TIELO_X1 D11611 ( .Y(D11611_Y));
KC_TIELO_X1 D11610 ( .Y(D11610_Y));
KC_TIELO_X1 D11609 ( .Y(D11609_Y));
KC_TIELO_X1 D11608 ( .Y(D11608_Y));
KC_TIELO_X1 D11590 ( .Y(D11590_Y));
KC_TIELO_X1 D11589 ( .Y(D11589_Y));
KC_TIELO_X1 D11418 ( .Y(D11418_Y));
KC_TIELO_X1 D11416 ( .Y(D11416_Y));
KC_TIELO_X1 D11349 ( .Y(D11349_Y));
KC_TIELO_X1 D11279 ( .Y(D11279_Y));
KC_TIELO_X1 D11186 ( .Y(D11186_Y));
KC_TIELO_X1 D11185 ( .Y(D11185_Y));
KC_TIELO_X1 D11184 ( .Y(D11184_Y));
KC_TIELO_X1 D11135 ( .Y(D11135_Y));
KC_TIELO_X1 D11117 ( .Y(D11117_Y));
KC_TIELO_X1 D11113 ( .Y(D11113_Y));
KC_TIELO_X1 D11089 ( .Y(D11089_Y));
KC_TIELO_X1 D11088 ( .Y(D11088_Y));
KC_TIELO_X1 D11057 ( .Y(D11057_Y));
KC_TIELO_X1 D11054 ( .Y(D11054_Y));
KC_TIELO_X1 D10898 ( .Y(D10898_Y));
KC_TIELO_X1 D10897 ( .Y(D10897_Y));
KC_TIELO_X1 D10896 ( .Y(D10896_Y));
KC_TIELO_X1 D10895 ( .Y(D10895_Y));
KC_TIELO_X1 D10830 ( .Y(D10830_Y));
KC_TIELO_X1 D10829 ( .Y(D10829_Y));
KC_TIELO_X1 D10129 ( .Y(D10129_Y));
KC_TIELO_X1 D9953 ( .Y(D9953_Y));
KC_TIELO_X1 D9952 ( .Y(D9952_Y));
KC_TIELO_X1 D9951 ( .Y(D9951_Y));
KC_TIELO_X1 D9921 ( .Y(D9921_Y));
KC_TIELO_X1 D9722 ( .Y(D9722_Y));
KC_TIELO_X1 D9721 ( .Y(D9721_Y));
KC_TIELO_X1 D9591 ( .Y(D9591_Y));
KC_TIELO_X1 D9229 ( .Y(D9229_Y));
KC_TIELO_X1 D16757 ( .Y(D16757_Y));
KC_TIELO_X1 D9165 ( .Y(D9165_Y));
KC_TIELO_X1 D8837 ( .Y(D8837_Y));
KC_TIELO_X1 D8662 ( .Y(D8662_Y));
KC_TIELO_X1 D8608 ( .Y(D8608_Y));
KC_TIELO_X1 D8606 ( .Y(D8606_Y));
KC_TIELO_X1 D8263 ( .Y(D8263_Y));
KC_TIELO_X1 D8260 ( .Y(D8260_Y));
KC_TIELO_X1 D8167 ( .Y(D8167_Y));
KC_TIELO_X1 D8166 ( .Y(D8166_Y));
KC_TIELO_X1 D8165 ( .Y(D8165_Y));
KC_TIELO_X1 D7993 ( .Y(D7993_Y));
KC_TIELO_X1 D7754 ( .Y(D7754_Y));
KC_TIELO_X1 D35 ( .Y(D35_Y));
KC_TIELO_X1 D12 ( .Y(D12_Y));
KC_TIELO_X1 D4 ( .Y(D4_Y));
KC_TIELO_X1 D7162 ( .Y(D7162_Y));
KC_TIELO_X1 D7161 ( .Y(D7161_Y));
KC_TIELO_X1 D6910 ( .Y(D6910_Y));
KC_TIELO_X1 D6833 ( .Y(D6833_Y));
KC_TIELO_X1 D6832 ( .Y(D6832_Y));
KC_TIELO_X1 D6617 ( .Y(D6617_Y));
KC_TIELO_X1 D6567 ( .Y(D6567_Y));
KC_TIELO_X1 D6497 ( .Y(D6497_Y));
KC_TIELO_X1 D6493 ( .Y(D6493_Y));
KC_TIELO_X1 D6488 ( .Y(D6488_Y));
KC_TIELO_X1 D6414 ( .Y(D6414_Y));
KC_TIELO_X1 D6413 ( .Y(D6413_Y));
KC_TIELO_X1 D6409 ( .Y(D6409_Y));
KC_TIELO_X1 D6358 ( .Y(D6358_Y));
KC_TIELO_X1 D6207 ( .Y(D6207_Y));
KC_TIELO_X1 D33 ( .Y(D33_Y));
KC_TIELO_X1 D30 ( .Y(D30_Y));
KC_TIELO_X1 D5823 ( .Y(D5823_Y));
KC_TIELO_X1 D5822 ( .Y(D5822_Y));
KC_TIELO_X1 D5706 ( .Y(D5706_Y));
KC_TIELO_X1 D5701 ( .Y(D5701_Y));
KC_TIELO_X1 D5490 ( .Y(D5490_Y));
KC_TIELO_X1 D5419 ( .Y(D5419_Y));
KC_TIELO_X1 D5331 ( .Y(D5331_Y));
KC_TIELO_X1 D5253 ( .Y(D5253_Y));
KC_TIELO_X1 D5252 ( .Y(D5252_Y));
KC_TIELO_X1 D5251 ( .Y(D5251_Y));
KC_TIELO_X1 D5250 ( .Y(D5250_Y));
KC_TIELO_X1 D4979 ( .Y(D4979_Y));
KC_TIELO_X1 D4742 ( .Y(D4742_Y));
KC_TIELO_X1 D4652 ( .Y(D4652_Y));
KC_TIELO_X1 D4073 ( .Y(D4073_Y));
KC_TIELO_X1 D4071 ( .Y(D4071_Y));
KC_TIELO_X1 D4070 ( .Y(D4070_Y));
KC_TIELO_X1 D4069 ( .Y(D4069_Y));
KC_TIELO_X1 D4031 ( .Y(D4031_Y));
KC_TIELO_X1 D4030 ( .Y(D4030_Y));
KC_TIELO_X1 D4029 ( .Y(D4029_Y));
KC_TIELO_X1 D3892 ( .Y(D3892_Y));
KC_TIELO_X1 D3891 ( .Y(D3891_Y));
KC_TIELO_X1 D3890 ( .Y(D3890_Y));
KC_TIELO_X1 D3889 ( .Y(D3889_Y));
KC_TIELO_X1 D3763 ( .Y(D3763_Y));
KC_TIELO_X1 D3762 ( .Y(D3762_Y));
KC_TIELO_X1 D3701 ( .Y(D3701_Y));
KC_TIELO_X1 D3399 ( .Y(D3399_Y));
KC_TIELO_X1 D3297 ( .Y(D3297_Y));
KC_TIELO_X1 D3201 ( .Y(D3201_Y));
KC_TIELO_X1 D3196 ( .Y(D3196_Y));
KC_TIELO_X1 D38 ( .Y(D38_Y));
KC_TIELO_X1 D2811 ( .Y(D2811_Y));
KC_TIELO_X1 D2526 ( .Y(D2526_Y));
KC_TIELO_X1 D2403 ( .Y(D2403_Y));
KC_TIELO_X1 D2105 ( .Y(D2105_Y));
KC_TIELO_X1 D1973 ( .Y(D1973_Y));
KC_TIELO_X1 D1972 ( .Y(D1972_Y));
KC_TIELO_X1 D1819 ( .Y(D1819_Y));
KC_TIELO_X1 D1818 ( .Y(D1818_Y));
KC_TIELO_X1 D1676 ( .Y(D1676_Y));
KC_TIELO_X1 D1675 ( .Y(D1675_Y));
KC_TIELO_X1 D1673 ( .Y(D1673_Y));
KC_TIELO_X1 D1535 ( .Y(D1535_Y));
KC_TIELO_X1 D270 ( .Y(D270_Y));
KC_NOR2_X3 D14886 ( .Y(D14886_Y), .B(D14688_Q), .A(D14687_Q));
KC_NOR2_X3 D14885 ( .Y(D14885_Y), .B(D14643_Y), .A(D14532_Y));
KC_NOR2_X3 D14884 ( .Y(D14884_Y), .B(D14532_Y), .A(D14688_Q));
KC_NOR2_X3 D14883 ( .Y(D14883_Y), .B(D14643_Y), .A(D14687_Q));
KC_NOR2_X3 D14882 ( .Y(D14882_Y), .B(D14643_Y), .A(D14532_Y));
KC_NOR2_X3 D14881 ( .Y(D14881_Y), .B(D14643_Y), .A(D14687_Q));
KC_NOR2_X3 D14880 ( .Y(D14880_Y), .B(D14688_Q), .A(D14687_Q));
KC_NOR2_X3 D14879 ( .Y(D14879_Y), .B(D14532_Y), .A(D14688_Q));
KC_NOR2_X3 D14698 ( .Y(D14698_Y), .B(D14667_Y), .A(D14621_Y));
KC_NOR2_X3 D14259 ( .Y(D14259_Y), .B(D763_Y), .A(D2495_Y));
KC_NOR2_X3 D14258 ( .Y(D14258_Y), .B(D14141_Y), .A(D13304_Y));
KC_NOR2_X3 D14257 ( .Y(D14257_Y), .B(D14141_Y), .A(D2437_Y));
KC_NOR2_X3 D14256 ( .Y(D14256_Y), .B(D763_Y), .A(D13304_Y));
KC_NOR2_X3 D14255 ( .Y(D14255_Y), .B(D14141_Y), .A(D2495_Y));
KC_NOR2_X3 D14254 ( .Y(D14254_Y), .B(D763_Y), .A(D13291_Y));
KC_NOR2_X3 D14253 ( .Y(D14253_Y), .B(D763_Y), .A(D2437_Y));
KC_NOR2_X3 D14252 ( .Y(D14252_Y), .B(D14141_Y), .A(D13291_Y));
KC_NOR2_X3 D14251 ( .Y(D14251_Y), .B(D14133_Y), .A(D874_Y));
KC_NOR2_X3 D14250 ( .Y(D14250_Y), .B(D14134_Y), .A(D874_Y));
KC_NOR2_X3 D14249 ( .Y(D14249_Y), .B(D14132_Y), .A(D874_Y));
KC_NOR2_X3 D14248 ( .Y(D14248_Y), .B(D874_Y), .A(D14137_Y));
KC_NOR2_X3 D14176 ( .Y(D14176_Y), .B(D14141_Y), .A(D750_Y));
KC_NOR2_X3 D14175 ( .Y(D14175_Y), .B(D763_Y), .A(D13310_Y));
KC_NOR2_X3 D14174 ( .Y(D14174_Y), .B(D763_Y), .A(D87_Y));
KC_NOR2_X3 D14173 ( .Y(D14173_Y), .B(D763_Y), .A(D750_Y));
KC_NOR2_X3 D14172 ( .Y(D14172_Y), .B(D14141_Y), .A(D13310_Y));
KC_NOR2_X3 D14171 ( .Y(D14171_Y), .B(D763_Y), .A(D13303_Y));
KC_NOR2_X3 D13400 ( .Y(D13400_Y), .B(D12747_Y), .A(D7609_Y));
KC_NOR2_X3 D12052 ( .Y(D12052_Y), .B(D11963_Y), .A(D11957_Y));
KC_NOR2_X3 D11991 ( .Y(D11991_Y), .B(D11904_Y), .A(D11946_Y));
KC_NOR2_X3 D11014 ( .Y(D11014_Y), .B(D10983_Y), .A(D10963_Y));
KC_NOR2_X3 D11013 ( .Y(D11013_Y), .B(D10984_Y), .A(D10964_Y));
KC_NOR2_X3 D11012 ( .Y(D11012_Y), .B(D10982_Y), .A(D10964_Y));
KC_NOR2_X3 D11011 ( .Y(D11011_Y), .B(D10984_Y), .A(D10963_Y));
KC_NOR2_X3 D11010 ( .Y(D11010_Y), .B(D10982_Y), .A(D10963_Y));
KC_NOR2_X3 D10818 ( .Y(D10818_Y), .B(D10762_Y), .A(D10747_Y));
KC_NOR2_X3 D10727 ( .Y(D10727_Y), .B(D10768_Y), .A(D10664_Y));
KC_NOR2_X3 D10560 ( .Y(D10560_Y), .B(D10479_Y), .A(D10536_Y));
KC_NOR2_X3 D10190 ( .Y(D10190_Y), .B(D10043_Y), .A(D2162_Y));
KC_NOR2_X3 D10189 ( .Y(D10189_Y), .B(D10044_Y), .A(D2162_Y));
KC_NOR2_X3 D10188 ( .Y(D10188_Y), .B(D8948_Y), .A(D2162_Y));
KC_NOR2_X3 D10175 ( .Y(D10175_Y), .B(D9015_Y), .A(D2162_Y));
KC_NOR2_X3 D10174 ( .Y(D10174_Y), .B(D2160_Y), .A(D2162_Y));
KC_NOR2_X3 D10173 ( .Y(D10173_Y), .B(D8815_Y), .A(D2162_Y));
KC_NOR2_X3 D10172 ( .Y(D10172_Y), .B(D8950_Y), .A(D2162_Y));
KC_NOR2_X3 D10171 ( .Y(D10171_Y), .B(D9013_Y), .A(D2162_Y));
KC_NOR2_X3 D10170 ( .Y(D10170_Y), .B(D10039_Y), .A(D2162_Y));
KC_NOR2_X3 D10166 ( .Y(D10166_Y), .B(D8973_Y), .A(D2162_Y));
KC_NOR2_X3 D10165 ( .Y(D10165_Y), .B(D9017_Y), .A(D2162_Y));
KC_NOR2_X3 D10150 ( .Y(D10150_Y), .B(D8949_Y), .A(D2162_Y));
KC_NOR2_X3 D10114 ( .Y(D10114_Y), .B(D8972_Y), .A(D10057_Y));
KC_NOR2_X3 D10113 ( .Y(D10113_Y), .B(D10028_Y), .A(D10057_Y));
KC_NOR2_X3 D10112 ( .Y(D10112_Y), .B(D9118_Y), .A(D10057_Y));
KC_NOR2_X3 D10111 ( .Y(D10111_Y), .B(D10000_Y), .A(D10057_Y));
KC_NOR2_X3 D10110 ( .Y(D10110_Y), .B(D8904_Y), .A(D10057_Y));
KC_NOR2_X3 D9482 ( .Y(D9482_Y), .B(D9417_Y), .A(D9414_Y));
KC_NOR2_X3 D9481 ( .Y(D9481_Y), .B(D9417_Y), .A(D9422_Y));
KC_NOR2_X3 D9480 ( .Y(D9480_Y), .B(D9417_Y), .A(D9424_Y));
KC_NOR2_X3 D9479 ( .Y(D9479_Y), .B(D9417_Y), .A(D10196_Y));
KC_NOR2_X3 D9478 ( .Y(D9478_Y), .B(D9417_Y), .A(D9425_Y));
KC_NOR2_X3 D9477 ( .Y(D9477_Y), .B(D9417_Y), .A(D9415_Y));
KC_NOR2_X3 D9476 ( .Y(D9476_Y), .B(D9417_Y), .A(D1994_Y));
KC_NOR2_X3 D9475 ( .Y(D9475_Y), .B(D9417_Y), .A(D9423_Y));
KC_NOR2_X3 D9473 ( .Y(D9473_Y), .B(D714_Q), .A(D9419_Y));
KC_NOR2_X3 D8901 ( .Y(D8901_Y), .B(D7396_Y), .A(D7460_Y));
KC_NOR2_X3 D8900 ( .Y(D8900_Y), .B(D5825_Y), .A(D7460_Y));
KC_NOR2_X3 D8348 ( .Y(D8348_Y), .B(D8350_Y), .A(D8290_Y));
KC_NOR2_X3 D7394 ( .Y(D7394_Y), .B(D7376_Y), .A(D5656_Y));
KC_NOR2_X3 D7153 ( .Y(D7153_Y), .B(D5659_Y), .A(D5668_Y));
KC_NOR2_X3 D6483 ( .Y(D6483_Y), .B(D5021_Y), .A(D1564_Y));
KC_NOR2_X3 D6077 ( .Y(D6077_Y), .B(D5973_Y), .A(D8838_Y));
KC_NOR2_X3 D5698 ( .Y(D5698_Y), .B(D5662_Y), .A(D5675_Y));
KC_NOR2_X3 D5413 ( .Y(D5413_Y), .B(D5375_Y), .A(D5361_Y));
KC_NOR2_X3 D3284 ( .Y(D3284_Y), .B(D3350_Y), .A(D3245_Y));
KC_NOR2_X3 D2519 ( .Y(D2519_Y), .B(D14141_Y), .A(D13303_Y));
KC_NOR2_X3 D2171 ( .Y(D2171_Y), .B(D9016_Y), .A(D2162_Y));
KC_NOR2_X3 D2170 ( .Y(D2170_Y), .B(D10485_Y), .A(D10965_Y));
KC_NOR2_X3 D2095 ( .Y(D2095_Y), .B(D9417_Y), .A(D9406_Y));
KC_NOR2_X3 D936 ( .Y(D936_Y), .B(D14141_Y), .A(D87_Y));
KC_NOR2_X3 D831 ( .Y(D831_Y), .B(D1598_Y), .A(D5267_Y));
KC_NOR2_X3 D266 ( .Y(D266_Y), .B(D5876_Y), .A(D4301_Y));
KC_BUF_X4 D13757 ( .Y(D13757_Y), .A(D14858_Y));
KC_BUF_X4 D9939 ( .Y(D9939_Y), .A(D196_Y));
KC_BUF_X4 D9938 ( .Y(D9938_Y), .A(D10103_Y));
KC_BUF_X4 D9937 ( .Y(D9937_Y), .A(D9976_Y));
KC_BUF_X4 D9936 ( .Y(D9936_Y), .A(D8713_Y));
KC_BUF_X4 D9267 ( .Y(D9267_Y), .A(D9272_Q));
KC_BUF_X4 D1934 ( .Y(D1934_Y), .A(D9360_Y));
KC_BUF_X4 D263 ( .Y(D263_Y), .A(D8882_Y));
KC_DFFRNHQ_X2 D13280 ( .Q(D13280_Q), .D(D13260_Y), .RN(D13194_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X2 D7477 ( .Q(D7477_Q), .D(D10139_Y), .RN(D9271_Y),     .CK(D10107_QN));
KC_DFFRNHQ_X2 D13097 ( .Q(D13097_Q), .D(D9295_Y), .RN(D7892_Y),     .CK(D9212_QN));
KC_DFFRNHQ_X2 D9336 ( .Q(D9336_Q), .D(D9317_Y), .RN(D7893_Y),     .CK(D9212_QN));
KC_DFFRNHQ_X2 D8836 ( .Q(D8836_Q), .D(D8800_Y), .RN(D8818_Y),     .CK(D5931_QN));
KC_DFFRNHQ_X2 D8835 ( .Q(D8835_Q), .D(D8802_Y), .RN(D8818_Y),     .CK(D5931_QN));
KC_DFFRNHQ_X2 D8730 ( .Q(D8730_Q), .D(D8695_Y), .RN(D7795_Y),     .CK(D9140_QN));
KC_DFFRNHQ_X2 D10753 ( .Q(D10753_Q), .D(D16164_Y), .RN(D9375_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X2 D8073 ( .Q(D8073_Q), .D(D8020_Y), .RN(D9374_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X2 D40 ( .Q(D40_Q), .D(D8969_Y), .RN(D4483_Y),     .CK(D7466_QN));
KC_DFFRNHQ_X2 D4137 ( .Q(D4137_Q), .D(D7482_Y), .RN(D4483_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X2 D8313 ( .Q(D8313_Q), .D(D4232_Y), .RN(D4461_Y),     .CK(D5799_Y));
KC_DFFRNHQ_X2 D4149 ( .Q(D4149_Q), .D(D4223_Y), .RN(D4461_Y),     .CK(D5931_QN));
KC_DFFRNHQ_X2 D7647 ( .Q(D7647_Q), .D(D3210_Y), .RN(D4827_Y),     .CK(D3271_QN));
KC_DFFRNHQ_X2 D723 ( .Q(D723_Q), .D(D13979_Y), .RN(D13194_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X2 D6248 ( .Q(D6248_Q), .D(D8988_Y), .RN(D324_Y),     .CK(D7466_QN));
KC_DFFRNHQ_X2 D239 ( .Q(D239_Q), .D(D4214_Y), .RN(D4461_Y),     .CK(D5931_QN));
KC_OAI211B_X1 D16517 ( .B(D16502_Y), .C1N(D13966_Y), .C0(D16524_Y),     .A(D16498_Y), .Y(D16517_Y));
KC_OAI211B_X1 D16478 ( .B(D13394_Y), .C1N(D16510_Y), .C0(D16404_Y),     .A(D16523_Y), .Y(D16478_Y));
KC_OAI211B_X1 D16400 ( .B(D14057_Y), .C1N(D16460_Y), .C0(D16386_Q),     .A(D1276_Y), .Y(D16400_Y));
KC_OAI211B_X1 D16175 ( .B(D16108_Y), .C1N(D16066_Y), .C0(D16106_Y),     .A(D16088_Y), .Y(D16175_Y));
KC_OAI211B_X1 D15599 ( .B(D15555_Y), .C1N(D15517_Y), .C0(D15532_Y),     .A(D15561_Y), .Y(D15599_Y));
KC_OAI211B_X1 D15598 ( .B(D15547_Y), .C1N(D15637_Y), .C0(D15464_Y),     .A(D15560_Y), .Y(D15598_Y));
KC_OAI211B_X1 D15220 ( .B(D15941_Y), .C1N(D15217_Q), .C0(D15237_Q),     .A(D14419_Y), .Y(D15220_Y));
KC_OAI211B_X1 D14803 ( .B(D14751_Y), .C1N(D820_Q), .C0(D14115_Y),     .A(D14102_Y), .Y(D14803_Y));
KC_OAI211B_X1 D14600 ( .B(D14555_Y), .C1N(D14518_Q), .C0(D14530_Y),     .A(D14703_Y), .Y(D14600_Y));
KC_OAI211B_X1 D10518 ( .B(D10515_Q), .C1N(D10926_Y), .C0(D8363_Y),     .A(D1919_Y), .Y(D10518_Y));
KC_OAI211B_X1 D9485 ( .B(D9443_Y), .C1N(D9431_Y), .C0(D9395_Y),     .A(D9443_Y), .Y(D9485_Y));
KC_OAI211B_X1 D8732 ( .B(D16756_Co), .C1N(D8665_Y), .C0(D8806_Y),     .A(D8665_Y), .Y(D8732_Y));
KC_OAI211B_X1 D8356 ( .B(D8294_Y), .C1N(D8294_Y), .C0(D9616_Y),     .A(D8358_Y), .Y(D8356_Y));
KC_OAI211B_X1 D8163 ( .B(D674_Q), .C1N(D5174_Y), .C0(D8186_Y),     .A(D7974_Y), .Y(D8163_Y));
KC_OAI211B_X1 D8162 ( .B(D8136_Y), .C1N(D9390_Y), .C0(D8151_Q),     .A(D8089_Y), .Y(D8162_Y));
KC_OAI211B_X1 D7749 ( .B(D7704_Y), .C1N(D6328_Y), .C0(D7752_Y),     .A(D7738_Y), .Y(D7749_Y));
KC_OAI211B_X1 D6354 ( .B(D6330_Y), .C1N(D6315_Y), .C0(D6326_Y),     .A(D6348_Y), .Y(D6354_Y));
KC_OAI211B_X1 D6353 ( .B(D403_Y), .C1N(D7_Y), .C0(D3325_Y),     .A(D4655_Y), .Y(D6353_Y));
KC_OAI211B_X1 D6283 ( .B(D6231_Y), .C1N(D6227_Y), .C0(D1771_Y),     .A(D6282_Y), .Y(D6283_Y));
KC_OAI211B_X1 D6282 ( .B(D6244_Y), .C1N(D6229_Y), .C0(D6231_Y),     .A(D6231_Y), .Y(D6282_Y));
KC_OAI211B_X1 D5702 ( .B(D4216_Y), .C1N(D5645_Y), .C0(D4113_Y),     .A(D4089_Y), .Y(D5702_Y));
KC_OAI211B_X1 D4842 ( .B(D4697_Y), .C1N(D4818_Q), .C0(D3325_Y),     .A(D4757_Y), .Y(D4842_Y));
KC_OAI211B_X1 D4841 ( .B(D4754_Y), .C1N(D273_Y), .C0(D3325_Y),     .A(D4746_Y), .Y(D4841_Y));
KC_OAI211B_X1 D50 ( .B(D3012_Y), .C1N(D4595_Y), .C0(D4524_Y),     .A(D310_Y), .Y(D50_Y));
KC_OAI211B_X1 D4264 ( .B(D4189_Y), .C1N(D4242_Y), .C0(D5786_Y),     .A(D5824_Y), .Y(D4264_Y));
KC_OAI211B_X1 D4145 ( .B(D1538_Y), .C1N(D4091_Y), .C0(D4547_Y),     .A(D4547_Y), .Y(D4145_Y));
KC_OAI211B_X1 D4138 ( .B(D4104_Y), .C1N(D4099_Y), .C0(D16135_Y),     .A(D4110_Y), .Y(D4138_Y));
KC_OAI211B_X1 D3490 ( .B(D3403_Y), .C1N(D4873_Y), .C0(D1447_Y),     .A(D4968_Y), .Y(D3490_Y));
KC_OAI211B_X1 D3195 ( .B(D3155_Y), .C1N(D4607_Y), .C0(D3155_Y),     .A(D3180_Y), .Y(D3195_Y));
KC_OAI211B_X1 D43 ( .B(D3086_Y), .C1N(D3017_Y), .C0(D3042_Y),     .A(D42_Y), .Y(D43_Y));
KC_OAI211B_X1 D42 ( .B(D3022_Y), .C1N(D3042_Y), .C0(D3022_Y),     .A(D3087_Y), .Y(D42_Y));
KC_OAI211B_X1 D39 ( .B(D3064_Y), .C1N(D3071_Y), .C0(D3053_Y),     .A(D3053_Y), .Y(D39_Y));
KC_OAI211B_X1 D52 ( .B(D2004_Y), .C1N(D7958_Y), .C0(D7447_Y),     .A(D9071_Y), .Y(D52_Y));
KC_OAI211B_X1 D24 ( .B(D5966_Y), .C1N(D7533_Q), .C0(D7430_Y),     .A(D8952_Q), .Y(D24_Y));
KC_OAI211B_X1 D1817 ( .B(D4961_Y), .C1N(D6361_Y), .C0(D6465_Y),     .A(D1695_Y), .Y(D1817_Y));
KC_OAI211B_X1 D1671 ( .B(D4873_Y), .C1N(D4915_Y), .C0(D3400_Y),     .A(D3599_Y), .Y(D1671_Y));
KC_OAI211B_X1 D849 ( .B(D10264_Y), .C1N(D10239_Q), .C0(D1985_Y),     .A(D9546_Y), .Y(D849_Y));
KC_OAI211B_X1 D393 ( .B(D7618_Y), .C1N(D7649_Y), .C0(D7701_Y),     .A(D7731_Y), .Y(D393_Y));
KC_OAI211B_X1 D367 ( .B(D337_Y), .C1N(D369_Y), .C0(D3141_Y),     .A(D3158_Y), .Y(D367_Y));
KC_OAI211B_X1 D11 ( .B(D7426_Y), .C1N(D6057_Y), .C0(D9_Y), .A(D6035_Y),     .Y(D11_Y));
KC_OAI211B_X1 D236 ( .B(D5942_Y), .C1N(D4238_Y), .C0(D4186_Y),     .A(D4190_Y), .Y(D236_Y));
KC_NOR3_X1 D16658 ( .B(D1373_Q), .Y(D16658_Y), .C(D16661_Y),     .A(D16684_Q));
KC_NOR3_X1 D16657 ( .B(D16656_Y), .Y(D16657_Y), .C(D16653_Y),     .A(D16604_Y));
KC_NOR3_X1 D16647 ( .B(D16650_Q), .Y(D16647_Y), .C(D1395_Q),     .A(D16681_Q));
KC_NOR3_X1 D16503 ( .B(D16491_Y), .Y(D16503_Y), .C(D16519_Y),     .A(D16514_Y));
KC_NOR3_X1 D16502 ( .B(D16529_Y), .Y(D16502_Y), .C(D16518_Y),     .A(D1343_Y));
KC_NOR3_X1 D16453 ( .B(D15986_Y), .Y(D16453_Y), .C(D16442_Y),     .A(D16372_Y));
KC_NOR3_X1 D16449 ( .B(D16439_Y), .Y(D16449_Y), .C(D16432_Y),     .A(D16470_Q));
KC_NOR3_X1 D16380 ( .B(D1378_Q), .Y(D16380_Y), .C(D16375_Y),     .A(D16471_Q));
KC_NOR3_X1 D16379 ( .B(D16438_Y), .Y(D16379_Y), .C(D16457_Y),     .A(D16425_Y));
KC_NOR3_X1 D16277 ( .B(D16291_Q), .Y(D16277_Y), .C(D16286_Y),     .A(D2681_Q));
KC_NOR3_X1 D16276 ( .B(D7609_Y), .Y(D16276_Y), .C(D14017_Y),     .A(D16771_Y));
KC_NOR3_X1 D16275 ( .B(D16261_Y), .Y(D16275_Y), .C(D16286_Y),     .A(D16265_Y));
KC_NOR3_X1 D16274 ( .B(D16290_Q), .Y(D16274_Y), .C(D16289_Q),     .A(D16291_Q));
KC_NOR3_X1 D16273 ( .B(D16290_Q), .Y(D16273_Y), .C(D16261_Y),     .A(D2681_Q));
KC_NOR3_X1 D16271 ( .B(D16292_Q), .Y(D16271_Y), .C(D16250_Y),     .A(D2681_Q));
KC_NOR3_X1 D16270 ( .B(D16266_Y), .Y(D16270_Y), .C(D16247_Y),     .A(D16256_Y));
KC_NOR3_X1 D16269 ( .B(D16289_Q), .Y(D16269_Y), .C(D16247_Y),     .A(D16292_Q));
KC_NOR3_X1 D15986 ( .B(D1378_Q), .Y(D15986_Y), .C(D16416_Y),     .A(D1324_Q));
KC_NOR3_X1 D15985 ( .B(D16449_Y), .Y(D15985_Y), .C(D15986_Y),     .A(D15969_Y));
KC_NOR3_X1 D14861 ( .B(D14195_Y), .Y(D14861_Y), .C(D14842_Y),     .A(D14907_Y));
KC_NOR3_X1 D14668 ( .B(D14662_Y), .Y(D14668_Y), .C(D14661_Y),     .A(D16608_Y));
KC_NOR3_X1 D14664 ( .B(D637_Y), .Y(D14664_Y), .C(D14667_Y),     .A(D14686_Q));
KC_NOR3_X1 D14663 ( .B(D14621_Y), .Y(D14663_Y), .C(D14666_Y),     .A(D722_Q));
KC_NOR3_X1 D14662 ( .B(D637_Y), .Y(D14662_Y), .C(D635_Y), .A(D722_Q));
KC_NOR3_X1 D14661 ( .B(D14620_Y), .Y(D14661_Y), .C(D14666_Y),     .A(D14686_Q));
KC_NOR3_X1 D14571 ( .B(D14520_Q), .Y(D14571_Y), .C(D13905_Y),     .A(D2574_Q));
KC_NOR3_X1 D14570 ( .B(D14520_Q), .Y(D14570_Y), .C(D13905_Y),     .A(D2574_Q));
KC_NOR3_X1 D14569 ( .B(D14520_Q), .Y(D14569_Y), .C(D13905_Y),     .A(D2574_Q));
KC_NOR3_X1 D14562 ( .B(D2574_Q), .Y(D14562_Y), .C(D14556_Y),     .A(D14518_Q));
KC_NOR3_X1 D14292 ( .B(D14338_Y), .Y(D14292_Y), .C(D1179_Y),     .A(D14201_Y));
KC_NOR3_X1 D14286 ( .B(D14202_Y), .Y(D14286_Y), .C(D14340_Y),     .A(D14436_Y));
KC_NOR3_X1 D13848 ( .B(D770_Y), .Y(D13848_Y), .C(D13845_Y),     .A(D2866_Y));
KC_NOR3_X1 D13506 ( .B(D7669_Y), .Y(D13506_Y), .C(D13477_Y),     .A(D13338_Y));
KC_NOR3_X1 D13368 ( .B(D2658_Y), .Y(D13368_Y), .C(D13332_Y),     .A(D16203_Y));
KC_NOR3_X1 D13281 ( .B(D12191_Y), .Y(D13281_Y), .C(D2409_Y),     .A(D7609_Y));
KC_NOR3_X1 D13246 ( .B(D13344_Y), .Y(D13246_Y), .C(D13255_Y),     .A(D13360_Y));
KC_NOR3_X1 D13243 ( .B(D14003_Y), .Y(D13243_Y), .C(D13950_Y),     .A(D13270_Q));
KC_NOR3_X1 D12731 ( .B(D12296_Y), .Y(D12731_Y), .C(D12708_Y),     .A(D12250_Y));
KC_NOR3_X1 D12729 ( .B(D12753_Q), .Y(D12729_Y), .C(D12813_Y),     .A(D12756_Q));
KC_NOR3_X1 D12725 ( .B(D12756_Q), .Y(D12725_Y), .C(D13268_Q),     .A(D12703_Y));
KC_NOR3_X1 D12260 ( .B(D2358_Y), .Y(D12260_Y), .C(D14806_Y),     .A(D12203_Y));
KC_NOR3_X1 D12259 ( .B(D12276_Y), .Y(D12259_Y), .C(D12362_Y),     .A(D850_Y));
KC_NOR3_X1 D12257 ( .B(D12657_Y), .Y(D12257_Y), .C(D12801_Y),     .A(D12371_Y));
KC_NOR3_X1 D12137 ( .B(D11183_Y), .Y(D12137_Y), .C(D12178_Q),     .A(D12143_Q));
KC_NOR3_X1 D11958 ( .B(D5376_Y), .Y(D11958_Y), .C(D11941_Y),     .A(D5377_Y));
KC_NOR3_X1 D11650 ( .B(D11645_Y), .Y(D11650_Y), .C(D11646_Y),     .A(D10181_Y));
KC_NOR3_X1 D10860 ( .B(D2146_Y), .Y(D10860_Y), .C(D98_Y),     .A(D10321_Y));
KC_NOR3_X1 D10767 ( .B(D5376_Y), .Y(D10767_Y), .C(D10729_Y),     .A(D5377_Y));
KC_NOR3_X1 D10155 ( .B(D723_Q), .Y(D10155_Y), .C(D10153_Y),     .A(D13285_Y));
KC_NOR3_X1 D10095 ( .B(D10091_Y), .Y(D10095_Y), .C(D10096_Y),     .A(D10089_Y));
KC_NOR3_X1 D10090 ( .B(D10089_Y), .Y(D10090_Y), .C(D10087_Y),     .A(D10197_Y));
KC_NOR3_X1 D10089 ( .B(D419_Q), .Y(D10089_Y), .C(D10100_Y),     .A(D9218_Q));
KC_NOR3_X1 D10087 ( .B(D10076_Y), .Y(D10087_Y), .C(D374_Y),     .A(D10071_Y));
KC_NOR3_X1 D10086 ( .B(D10076_Y), .Y(D10086_Y), .C(D10100_Y),     .A(D10071_Y));
KC_NOR3_X1 D10085 ( .B(D419_Q), .Y(D10085_Y), .C(D368_Y), .A(D9218_Q));
KC_NOR3_X1 D9544 ( .B(D9574_Q), .Y(D9544_Y), .C(D9522_Y), .A(D9577_Q));
KC_NOR3_X1 D9439 ( .B(D9420_Y), .Y(D9439_Y), .C(D9490_Y), .A(D624_Y));
KC_NOR3_X1 D9245 ( .B(D9285_Y), .Y(D9245_Y), .C(D9285_Y), .A(D9234_Y));
KC_NOR3_X1 D8992 ( .B(D8977_Y), .Y(D8992_Y), .C(D8975_Y), .A(D8978_Y));
KC_NOR3_X1 D8991 ( .B(D9027_Y), .Y(D8991_Y), .C(D9020_Y), .A(D9022_Y));
KC_NOR3_X1 D8938 ( .B(D2076_Y), .Y(D8938_Y), .C(D8943_Y), .A(D8944_Y));
KC_NOR3_X1 D8937 ( .B(D7_Y), .Y(D8937_Y), .C(D272_Y), .A(D273_Y));
KC_NOR3_X1 D8787 ( .B(D8806_Y), .Y(D8787_Y), .C(D8732_Y), .A(D5733_Y));
KC_NOR3_X1 D8778 ( .B(D8751_Y), .Y(D8778_Y), .C(D9480_Y), .A(D7183_Y));
KC_NOR3_X1 D8772 ( .B(D8781_Y), .Y(D8772_Y), .C(D204_Y), .A(D8756_Y));
KC_NOR3_X1 D8221 ( .B(D8204_Y), .Y(D8221_Y), .C(D1840_Y), .A(D8250_Q));
KC_NOR3_X1 D8215 ( .B(D8183_Y), .Y(D8215_Y), .C(D8192_Y), .A(D8261_Y));
KC_NOR3_X1 D7953 ( .B(D7943_Y), .Y(D7953_Y), .C(D7919_Y), .A(D7921_Y));
KC_NOR3_X1 D7776 ( .B(D12301_Y), .Y(D7776_Y), .C(D12762_Y),     .A(D725_Y));
KC_NOR3_X1 D7697 ( .B(D7688_Y), .Y(D7697_Y), .C(D7685_Y), .A(D7675_Y));
KC_NOR3_X1 D7671 ( .B(D7622_Y), .Y(D7671_Y), .C(D7672_Y), .A(D7700_Y));
KC_NOR3_X1 D7512 ( .B(D7750_Y), .Y(D7512_Y), .C(D13280_Q),     .A(D10142_Y));
KC_NOR3_X1 D7456 ( .B(D5685_Y), .Y(D7456_Y), .C(D7429_Y), .A(D7361_Y));
KC_NOR3_X1 D7455 ( .B(D7184_Y), .Y(D7455_Y), .C(D268_Q), .A(D7470_Y));
KC_NOR3_X1 D7375 ( .B(D7153_Y), .Y(D7375_Y), .C(D7343_Y), .A(D7109_Y));
KC_NOR3_X1 D7374 ( .B(D7352_Y), .Y(D7374_Y), .C(D7384_Y), .A(D7344_Y));
KC_NOR3_X1 D7368 ( .B(D5908_Y), .Y(D7368_Y), .C(D583_Co), .A(D7382_Y));
KC_NOR3_X1 D7362 ( .B(D7318_Y), .Y(D7362_Y), .C(D7323_Y), .A(D7409_Q));
KC_NOR3_X1 D7307 ( .B(D5647_Y), .Y(D7307_Y), .C(D7308_Y), .A(D7219_Y));
KC_NOR3_X1 D7263 ( .B(D7247_Y), .Y(D7263_Y), .C(D7258_Y), .A(D7246_Y));
KC_NOR3_X1 D6883 ( .B(D6808_Y), .Y(D6883_Y), .C(D6854_Y), .A(D6809_Y));
KC_NOR3_X1 D6878 ( .B(D8222_Y), .Y(D6878_Y), .C(D1685_Y), .A(D5461_Y));
KC_NOR3_X1 D6452 ( .B(D6531_Y), .Y(D6452_Y), .C(D6422_Y), .A(D6422_Y));
KC_NOR3_X1 D6451 ( .B(D6431_Y), .Y(D6451_Y), .C(D6483_Y), .A(D7929_Y));
KC_NOR3_X1 D6311 ( .B(D6339_Y), .Y(D6311_Y), .C(D6339_Y), .A(D6318_Y));
KC_NOR3_X1 D6236 ( .B(D6240_Y), .Y(D6236_Y), .C(D9144_Y), .A(D6268_Y));
KC_NOR3_X1 D6163 ( .B(D6164_Y), .Y(D6163_Y), .C(D6194_Y), .A(D6162_Y));
KC_NOR3_X1 D6154 ( .B(D7657_Y), .Y(D6154_Y), .C(D7585_Y), .A(D378_Y));
KC_NOR3_X1 D6152 ( .B(D1741_Y), .Y(D6152_Y), .C(D1790_Y), .A(D1790_Y));
KC_NOR3_X1 D6104 ( .B(D6084_Y), .Y(D6104_Y), .C(D6165_Y), .A(D6118_Y));
KC_NOR3_X1 D6103 ( .B(D322_Y), .Y(D6103_Y), .C(D6165_Y), .A(D6084_Y));
KC_NOR3_X1 D6101 ( .B(D6102_Y), .Y(D6101_Y), .C(D6118_Y), .A(D322_Y));
KC_NOR3_X1 D6046 ( .B(D6011_Y), .Y(D6046_Y), .C(D284_Y), .A(D6044_Y));
KC_NOR3_X1 D5917 ( .B(D1592_Y), .Y(D5917_Y), .C(D5997_Y), .A(D5999_Y));
KC_NOR3_X1 D5903 ( .B(D5828_Y), .Y(D5903_Y), .C(D244_Y), .A(D5852_Y));
KC_NOR3_X1 D5899 ( .B(D1719_Y), .Y(D5899_Y), .C(D7103_Y), .A(D7164_Y));
KC_NOR3_X1 D5898 ( .B(D5877_Y), .Y(D5898_Y), .C(D5829_Y), .A(D7164_Y));
KC_NOR3_X1 D5671 ( .B(D5655_Y), .Y(D5671_Y), .C(D5662_Y), .A(D5664_Y));
KC_NOR3_X1 D5454 ( .B(D5376_Y), .Y(D5454_Y), .C(D5442_Y), .A(D5377_Y));
KC_NOR3_X1 D5450 ( .B(D760_Y), .Y(D5450_Y), .C(D5431_Y), .A(D1628_Y));
KC_NOR3_X1 D5369 ( .B(D5385_Y), .Y(D5369_Y), .C(D5295_Y), .A(D5393_Y));
KC_NOR3_X1 D5052 ( .B(D5053_Y), .Y(D5052_Y), .C(D4984_Y), .A(D5048_Y));
KC_NOR3_X1 D5051 ( .B(D475_Y), .Y(D5051_Y), .C(D4994_Y), .A(D5080_Y));
KC_NOR3_X1 D5047 ( .B(D6437_Y), .Y(D5047_Y), .C(D5055_Y), .A(D5094_Y));
KC_NOR3_X1 D4941 ( .B(D4886_Y), .Y(D4941_Y), .C(D4960_Y), .A(D5009_Y));
KC_NOR3_X1 D4938 ( .B(D6371_Y), .Y(D4938_Y), .C(D4910_Y), .A(D6381_Q));
KC_NOR3_X1 D4930 ( .B(D432_Y), .Y(D4930_Y), .C(D6427_Y), .A(D3540_Y));
KC_NOR3_X1 D4703 ( .B(D4680_Y), .Y(D4703_Y), .C(D4734_Y), .A(D4670_Y));
KC_NOR3_X1 D4609 ( .B(D4650_Y), .Y(D4609_Y), .C(D4589_Y), .A(D4594_Y));
KC_NOR3_X1 D47 ( .B(D3016_Y), .Y(D47_Y), .C(D46_Y), .A(D3080_Q));
KC_NOR3_X1 D4520 ( .B(D4499_Y), .Y(D4520_Y), .C(D1609_Y), .A(D4508_Y));
KC_NOR3_X1 D4457 ( .B(D4417_Y), .Y(D4457_Y), .C(D4453_Y), .A(D4149_Q));
KC_NOR3_X1 D4456 ( .B(D4453_Y), .Y(D4456_Y), .C(D4422_Y), .A(D4421_Y));
KC_NOR3_X1 D4455 ( .B(D4429_Y), .Y(D4455_Y), .C(D4177_Y), .A(D6009_Y));
KC_NOR3_X1 D4452 ( .B(D4416_Y), .Y(D4452_Y), .C(D4420_Y), .A(D8313_Q));
KC_NOR3_X1 D4373 ( .B(D4328_Y), .Y(D4373_Y), .C(D4349_Y), .A(D7737_Q));
KC_NOR3_X1 D4368 ( .B(D4425_Y), .Y(D4368_Y), .C(D239_Q), .A(D4422_Y));
KC_NOR3_X1 D4105 ( .B(D4100_Y), .Y(D4105_Y), .C(D4117_Y), .A(D4138_Y));
KC_NOR3_X1 D4077 ( .B(D4038_Y), .Y(D4077_Y), .C(D4035_Y), .A(D4079_Y));
KC_NOR3_X1 D3849 ( .B(D3832_Y), .Y(D3849_Y), .C(D3936_Q), .A(D1478_Y));
KC_NOR3_X1 D3545 ( .B(D3446_Y), .Y(D3545_Y), .C(D6478_Y), .A(D4882_Y));
KC_NOR3_X1 D3349 ( .B(D3332_Y), .Y(D3349_Y), .C(D3369_Y), .A(D3347_Y));
KC_NOR3_X1 D3348 ( .B(D3362_Y), .Y(D3348_Y), .C(D3330_Y), .A(D3346_Y));
KC_NOR3_X1 D3346 ( .B(D3369_Y), .Y(D3346_Y), .C(D3351_Y), .A(D3384_Q));
KC_NOR3_X1 D3345 ( .B(D15265_Y), .Y(D3345_Y), .C(D3359_Y),     .A(D3344_Y));
KC_NOR3_X1 D3343 ( .B(D3377_Y), .Y(D3343_Y), .C(D3315_Y), .A(D1454_Y));
KC_NOR3_X1 D3341 ( .B(D3352_Y), .Y(D3341_Y), .C(D3390_Y), .A(D3307_Y));
KC_NOR3_X1 D3336 ( .B(D3306_Y), .Y(D3336_Y), .C(D3521_Y), .A(D3375_Q));
KC_NOR3_X1 D3298 ( .B(D3270_Y), .Y(D3298_Y), .C(D3299_Y), .A(D3368_Y));
KC_NOR3_X1 D3256 ( .B(D3281_Q), .Y(D3256_Y), .C(D3283_Q), .A(D3282_Q));
KC_NOR3_X1 D3254 ( .B(D3232_Y), .Y(D3254_Y), .C(D1423_Y), .A(D1425_Y));
KC_NOR3_X1 D3252 ( .B(D4666_Y), .Y(D3252_Y), .C(D4682_Y), .A(D4592_Y));
KC_NOR3_X1 D3251 ( .B(D3154_Y), .Y(D3251_Y), .C(D3228_Y), .A(D3261_Y));
KC_NOR3_X1 D3250 ( .B(D3221_Y), .Y(D3250_Y), .C(D3350_Y), .A(D3273_Y));
KC_NOR3_X1 D3247 ( .B(D3270_Y), .Y(D3247_Y), .C(D3368_Y), .A(D3273_Y));
KC_NOR3_X1 D3165 ( .B(D1457_Y), .Y(D3165_Y), .C(D3145_Y), .A(D3132_Y));
KC_NOR3_X1 D3161 ( .B(D3123_Y), .Y(D3161_Y), .C(D3174_Y), .A(D3162_Y));
KC_NOR3_X1 D44 ( .B(D1515_Q), .Y(D44_Y), .C(D45_Y), .A(D3080_Q));
KC_NOR3_X1 D3042 ( .B(D3019_Y), .Y(D3042_Y), .C(D3027_Y), .A(D3062_Y));
KC_NOR3_X1 D3041 ( .B(D3023_Y), .Y(D3041_Y), .C(D3028_Y), .A(D3080_Q));
KC_NOR3_X1 D3040 ( .B(D3014_Y), .Y(D3040_Y), .C(D3043_Y), .A(D3028_Y));
KC_NOR3_X1 D3039 ( .B(D3084_Q), .Y(D3039_Y), .C(D3015_Y), .A(D1516_Q));
KC_NOR3_X1 D3038 ( .B(D3028_Y), .Y(D3038_Y), .C(D3013_Y), .A(D3084_Q));
KC_NOR3_X1 D3037 ( .B(D3020_Y), .Y(D3037_Y), .C(D3028_Y), .A(D1515_Q));
KC_NOR3_X1 D2782 ( .B(D2799_Q), .Y(D2782_Y), .C(D2798_Q), .A(D2797_Q));
KC_NOR3_X1 D2780 ( .B(D2796_Q), .Y(D2780_Y), .C(D2795_Q), .A(D2794_Q));
KC_NOR3_X1 D2628 ( .B(D16597_Y), .Y(D2628_Y), .C(D16264_Y),     .A(D2617_Y));
KC_NOR3_X1 D2454 ( .B(D12757_Y), .Y(D2454_Y), .C(D12720_Y),     .A(D12191_Y));
KC_NOR3_X1 D2330 ( .B(D6287_Y), .Y(D2330_Y), .C(D12186_Y),     .A(D2353_Y));
KC_NOR3_X1 D1617 ( .B(D4173_Y), .Y(D1617_Y), .C(D4234_Y), .A(D4119_Q));
KC_NOR3_X1 D1595 ( .B(D1653_Y), .Y(D1595_Y), .C(D2716_Y), .A(D4091_Y));
KC_NOR3_X1 D1456 ( .B(D3184_Q), .Y(D1456_Y), .C(D3234_Y), .A(D3117_Y));
KC_NOR3_X1 D1344 ( .B(D16535_Y), .Y(D1344_Y), .C(D16487_Y),     .A(D16536_Y));
KC_NOR3_X1 D647 ( .B(D721_Q), .Y(D647_Y), .C(D14620_Y), .A(D14689_Q));
KC_NOR3_X1 D646 ( .B(D16107_Y), .Y(D646_Y), .C(D16121_Y), .A(D650_Y));
KC_NOR3_X1 D643 ( .B(D703_Q), .Y(D643_Y), .C(D2063_Y), .A(D7655_Y));
KC_NOR3_X1 D573 ( .B(D608_Q), .Y(D573_Y), .C(D14540_Y), .A(D14519_Q));
KC_NOR3_X1 D436 ( .B(D4898_Y), .Y(D436_Y), .C(D4889_Y), .A(D3400_Y));
KC_NOR3_X1 D312 ( .B(D3084_Q), .Y(D312_Y), .C(D3020_Y), .A(D1516_Q));
KC_NOR3_X1 D291 ( .B(D4425_Y), .Y(D291_Y), .C(D4419_Y), .A(D6096_Y));
KC_NOR3_X1 D220 ( .B(D7183_Y), .Y(D220_Y), .C(D8783_Y), .A(D9481_Y));
KC_NAND3_X1 D16547 ( .Y(D16547_Y), .C(D1385_Q), .B(D16556_Q),     .A(D16493_Y));
KC_NAND3_X1 D16545 ( .Y(D16545_Y), .C(D16528_Y), .B(D1381_Q),     .A(D16556_Q));
KC_NAND3_X1 D16508 ( .Y(D16508_Y), .C(D16495_Y), .B(D16496_Y),     .A(D16382_Y));
KC_NAND3_X1 D16507 ( .Y(D16507_Y), .C(D16490_Y), .B(D16492_Y),     .A(D16559_Y));
KC_NAND3_X1 D16505 ( .Y(D16505_Y), .C(D16488_Y), .B(D16538_Y),     .A(D16539_Y));
KC_NAND3_X1 D16504 ( .Y(D16504_Y), .C(D13988_Y), .B(D16530_Y),     .A(D14651_Y));
KC_NAND3_X1 D16461 ( .Y(D16461_Y), .C(D16426_Y), .B(D16380_Y),     .A(D16436_Y));
KC_NAND3_X1 D16454 ( .Y(D16454_Y), .C(D16443_Y), .B(D16441_Y),     .A(D1324_Q));
KC_NAND3_X1 D16452 ( .Y(D16452_Y), .C(D16438_Y), .B(D16419_Y),     .A(D16436_Y));
KC_NAND3_X1 D16448 ( .Y(D16448_Y), .C(D16444_Y), .B(D16470_Q),     .A(D16459_Q));
KC_NAND3_X1 D16446 ( .Y(D16446_Y), .C(D16407_Y), .B(D16382_Y),     .A(D16430_Y));
KC_NAND3_X1 D16378 ( .Y(D16378_Y), .C(D14057_Y), .B(D16268_Y),     .A(D16374_Y));
KC_NAND3_X1 D16272 ( .Y(D16272_Y), .C(D16266_Y), .B(D16281_Y),     .A(D16293_Q));
KC_NAND3_X1 D16268 ( .Y(D16268_Y), .C(D16257_Y), .B(D16287_Q),     .A(D16279_Y));
KC_NAND3_X1 D16125 ( .Y(D16125_Y), .C(D16119_Y), .B(D16114_Y),     .A(D15311_Y));
KC_NAND3_X1 D16068 ( .Y(D16068_Y), .C(D16043_Y), .B(D16054_Y),     .A(D16094_Y));
KC_NAND3_X1 D16067 ( .Y(D16067_Y), .C(D16054_Y), .B(D16094_Y),     .A(D16059_Y));
KC_NAND3_X1 D15660 ( .Y(D15660_Y), .C(D15698_Y), .B(D2613_Y),     .A(D15641_Y));
KC_NAND3_X1 D15659 ( .Y(D15659_Y), .C(D2612_Y), .B(D15644_Y),     .A(D15643_Y));
KC_NAND3_X1 D15555 ( .Y(D15555_Y), .C(D8886_Y), .B(D15349_Y),     .A(D15522_Y));
KC_NAND3_X1 D15550 ( .Y(D15550_Y), .C(D14564_Y), .B(D2644_Y),     .A(D15563_Y));
KC_NAND3_X1 D15547 ( .Y(D15547_Y), .C(D2870_Y), .B(D2604_Y),     .A(D14813_Y));
KC_NAND3_X1 D15428 ( .Y(D15428_Y), .C(D2590_Y), .B(D15407_Y),     .A(D15409_Y));
KC_NAND3_X1 D15424 ( .Y(D15424_Y), .C(D15454_Y), .B(D15536_Y),     .A(D633_Y));
KC_NAND3_X1 D15423 ( .Y(D15423_Y), .C(D2590_Y), .B(D15407_Y),     .A(D15397_Y));
KC_NAND3_X1 D15422 ( .Y(D15422_Y), .C(D2590_Y), .B(D15408_Y),     .A(D15409_Y));
KC_NAND3_X1 D15421 ( .Y(D15421_Y), .C(D2590_Y), .B(D15408_Y),     .A(D15397_Y));
KC_NAND3_X1 D15420 ( .Y(D15420_Y), .C(D2590_Y), .B(D15408_Y),     .A(D15327_Y));
KC_NAND3_X1 D15419 ( .Y(D15419_Y), .C(D2590_Y), .B(D15407_Y),     .A(D15327_Y));
KC_NAND3_X1 D15418 ( .Y(D15418_Y), .C(D15564_Y), .B(D14531_Y),     .A(D816_Q));
KC_NAND3_X1 D15415 ( .Y(D15415_Y), .C(D15455_Y), .B(D15368_Y),     .A(D15343_Y));
KC_NAND3_X1 D15410 ( .Y(D15410_Y), .C(D15356_Y), .B(D15398_Y),     .A(D15347_Y));
KC_NAND3_X1 D15314 ( .Y(D15314_Y), .C(D2587_Y), .B(D15272_Y),     .A(D15326_Y));
KC_NAND3_X1 D15313 ( .Y(D15313_Y), .C(D2587_Y), .B(D15309_Y),     .A(D15272_Y));
KC_NAND3_X1 D15312 ( .Y(D15312_Y), .C(D2587_Y), .B(D15320_Y),     .A(D15273_Y));
KC_NAND3_X1 D15194 ( .Y(D15194_Y), .C(D16000_Y), .B(D14085_Y),     .A(D15164_Y));
KC_NAND3_X1 D15112 ( .Y(D15112_Y), .C(D15943_Y), .B(D13982_Y),     .A(D15099_Y));
KC_NAND3_X1 D15067 ( .Y(D15067_Y), .C(D2527_Y), .B(D15911_Y),     .A(D2528_Y));
KC_NAND3_X1 D15065 ( .Y(D15065_Y), .C(D15865_Y), .B(D13983_Y),     .A(D15032_Y));
KC_NAND3_X1 D15061 ( .Y(D15061_Y), .C(D15011_Y), .B(D15833_Y),     .A(D15041_Y));
KC_NAND3_X1 D15055 ( .Y(D15055_Y), .C(D15023_Y), .B(D15815_Y),     .A(D15024_Y));
KC_NAND3_X1 D14977 ( .Y(D14977_Y), .C(D1075_Y), .B(D14086_Y),     .A(D2537_Y));
KC_NAND3_X1 D14976 ( .Y(D14976_Y), .C(D14948_Y), .B(D14957_Y),     .A(D14958_Y));
KC_NAND3_X1 D14975 ( .Y(D14975_Y), .C(D14951_Y), .B(D15732_Y),     .A(D14954_Y));
KC_NAND3_X1 D14969 ( .Y(D14969_Y), .C(D15720_Y), .B(D14924_Y),     .A(D14933_Y));
KC_NAND3_X1 D14965 ( .Y(D14965_Y), .C(D14994_Y), .B(D1155_Q),     .A(D14021_Y));
KC_NAND3_X1 D14964 ( .Y(D14964_Y), .C(D14914_Y), .B(D15825_Y),     .A(D14920_Y));
KC_NAND3_X1 D14962 ( .Y(D14962_Y), .C(D14937_Y), .B(D15717_Y),     .A(D14932_Y));
KC_NAND3_X1 D14864 ( .Y(D14864_Y), .C(D14718_Y), .B(D14878_Q),     .A(D853_Q));
KC_NAND3_X1 D14857 ( .Y(D14857_Y), .C(D2584_Y), .B(D14002_Y),     .A(D2538_Y));
KC_NAND3_X1 D14670 ( .Y(D14670_Y), .C(D13988_Y), .B(D14662_Y),     .A(D14651_Y));
KC_NAND3_X1 D14669 ( .Y(D14669_Y), .C(D14662_Y), .B(D14651_Y),     .A(D14650_Y));
KC_NAND3_X1 D14666 ( .Y(D14666_Y), .C(D14622_Y), .B(D14630_Y),     .A(D721_Q));
KC_NAND3_X1 D14665 ( .Y(D14665_Y), .C(D637_Y), .B(D14619_Y),     .A(D13945_Y));
KC_NAND3_X1 D14572 ( .Y(D14572_Y), .C(D14539_Y), .B(D14708_Y),     .A(D608_Q));
KC_NAND3_X1 D14567 ( .Y(D14567_Y), .C(D14571_Y), .B(D14601_Q),     .A(D608_Q));
KC_NAND3_X1 D14564 ( .Y(D14564_Y), .C(D14570_Y), .B(D14601_Q),     .A(D608_Q));
KC_NAND3_X1 D14563 ( .Y(D14563_Y), .C(D14569_Y), .B(D14601_Q),     .A(D608_Q));
KC_NAND3_X1 D14369 ( .Y(D14369_Y), .C(D14471_Y), .B(D14090_Y),     .A(D14356_Y));
KC_NAND3_X1 D14366 ( .Y(D14366_Y), .C(D14470_Y), .B(D14089_Y),     .A(D14348_Y));
KC_NAND3_X1 D14361 ( .Y(D14361_Y), .C(D14476_Y), .B(D14082_Y),     .A(D14343_Y));
KC_NAND3_X1 D14289 ( .Y(D14289_Y), .C(D14294_Y), .B(D14293_Y),     .A(D14295_Y));
KC_NAND3_X1 D14149 ( .Y(D14149_Y), .C(D14030_Y), .B(D14170_Q),     .A(D14092_Q));
KC_NAND3_X1 D14148 ( .Y(D14148_Y), .C(D14134_Y), .B(D14008_Y),     .A(D13317_Y));
KC_NAND3_X1 D14143 ( .Y(D14143_Y), .C(D14193_Y), .B(D777_Y),     .A(D14127_Y));
KC_NAND3_X1 D14065 ( .Y(D14065_Y), .C(D14044_Y), .B(D14665_Y),     .A(D13977_Y));
KC_NAND3_X1 D14054 ( .Y(D14054_Y), .C(D14137_Y), .B(D14008_Y),     .A(D13478_Y));
KC_NAND3_X1 D13970 ( .Y(D13970_Y), .C(D13953_Y), .B(D13939_Y),     .A(D14785_Y));
KC_NAND3_X1 D13969 ( .Y(D13969_Y), .C(D14649_Y), .B(D13953_Y),     .A(D14664_Y));
KC_NAND3_X1 D13965 ( .Y(D13965_Y), .C(D13257_Y), .B(D16117_Y),     .A(D13184_Y));
KC_NAND3_X1 D13787 ( .Y(D13787_Y), .C(D13775_Y), .B(D14446_Y),     .A(D13810_Q));
KC_NAND3_X1 D13741 ( .Y(D13741_Y), .C(D13753_Y), .B(D13987_Y),     .A(D13729_Y));
KC_NAND3_X1 D13692 ( .Y(D13692_Y), .C(D13700_Y), .B(D778_Y),     .A(D2414_Y));
KC_NAND3_X1 D13603 ( .Y(D13603_Y), .C(D2435_Y), .B(D13578_Y),     .A(D13553_Y));
KC_NAND3_X1 D13602 ( .Y(D13602_Y), .C(D2438_Y), .B(D13578_Y),     .A(D13553_Y));
KC_NAND3_X1 D13601 ( .Y(D13601_Y), .C(D13007_Y), .B(D13599_Y),     .A(D13499_Y));
KC_NAND3_X1 D13599 ( .Y(D13599_Y), .C(D2371_Y), .B(D14246_Q),     .A(D12944_Y));
KC_NAND3_X1 D13503 ( .Y(D13503_Y), .C(D13521_Y), .B(D13492_Y),     .A(D13499_Y));
KC_NAND3_X1 D13499 ( .Y(D13499_Y), .C(D13323_Y), .B(D12905_Y),     .A(D13460_Y));
KC_NAND3_X1 D13498 ( .Y(D13498_Y), .C(D13520_Y), .B(D13491_Y),     .A(D13499_Y));
KC_NAND3_X1 D13492 ( .Y(D13492_Y), .C(D13467_Y), .B(D926_Q),     .A(D12944_Y));
KC_NAND3_X1 D13491 ( .Y(D13491_Y), .C(D13456_Y), .B(D12944_Y),     .A(D14166_Q));
KC_NAND3_X1 D13487 ( .Y(D13487_Y), .C(D13517_Y), .B(D13481_Y),     .A(D13499_Y));
KC_NAND3_X1 D13481 ( .Y(D13481_Y), .C(D13430_Y), .B(D14167_Q),     .A(D12944_Y));
KC_NAND3_X1 D13374 ( .Y(D13374_Y), .C(D13355_Y), .B(D12766_Y),     .A(D14066_Y));
KC_NAND3_X1 D13372 ( .Y(D13372_Y), .C(D13352_Y), .B(D13398_Q),     .A(D13333_Y));
KC_NAND3_X1 D13370 ( .Y(D13370_Y), .C(D13346_Y), .B(D13327_Y),     .A(D13395_Q));
KC_NAND3_X1 D13369 ( .Y(D13369_Y), .C(D13335_Y), .B(D13398_Q),     .A(D13397_Q));
KC_NAND3_X1 D13247 ( .Y(D13247_Y), .C(D13403_Y), .B(D13364_Y),     .A(D13234_Y));
KC_NAND3_X1 D13154 ( .Y(D13154_Y), .C(D13166_Y), .B(D13168_Y),     .A(D13165_Y));
KC_NAND3_X1 D12965 ( .Y(D12965_Y), .C(D13008_Y), .B(D997_Y),     .A(D13499_Y));
KC_NAND3_X1 D12964 ( .Y(D12964_Y), .C(D13006_Y), .B(D995_Y),     .A(D13499_Y));
KC_NAND3_X1 D12823 ( .Y(D12823_Y), .C(D12815_Y), .B(D12729_Y),     .A(D13268_Q));
KC_NAND3_X1 D12820 ( .Y(D12820_Y), .C(D12823_Y), .B(D12797_Y),     .A(D12856_Q));
KC_NAND3_X1 D12816 ( .Y(D12816_Y), .C(D12814_Y), .B(D13268_Q),     .A(D12754_Q));
KC_NAND3_X1 D12733 ( .Y(D12733_Y), .C(D12754_Q), .B(D12753_Q),     .A(D13268_Q));
KC_NAND3_X1 D12732 ( .Y(D12732_Y), .C(D658_Y), .B(D12729_Y),     .A(D12714_Y));
KC_NAND3_X1 D12261 ( .Y(D12261_Y), .C(D12206_Y), .B(D11657_Y),     .A(D11655_Y));
KC_NAND3_X1 D12210 ( .Y(D12210_Y), .C(D12255_Y), .B(D12273_Y),     .A(D12692_Y));
KC_NAND3_X1 D12032 ( .Y(D12032_Y), .C(D1143_Y), .B(D12028_Y),     .A(D6793_Y));
KC_NAND3_X1 D12031 ( .Y(D12031_Y), .C(D10514_Y), .B(D12028_Y),     .A(D6791_Y));
KC_NAND3_X1 D12030 ( .Y(D12030_Y), .C(D12028_Y), .B(D6793_Y),     .A(D6791_Y));
KC_NAND3_X1 D11965 ( .Y(D11965_Y), .C(D11421_Y), .B(D5376_Y),     .A(D5377_Y));
KC_NAND3_X1 D11964 ( .Y(D11964_Y), .C(D5479_Y), .B(D11421_Y),     .A(D5377_Y));
KC_NAND3_X1 D11963 ( .Y(D11963_Y), .C(D5480_Y), .B(D11421_Y),     .A(D5376_Y));
KC_NAND3_X1 D11962 ( .Y(D11962_Y), .C(D10514_Y), .B(D11954_Y),     .A(D6791_Y));
KC_NAND3_X1 D11961 ( .Y(D11961_Y), .C(D1143_Y), .B(D11954_Y),     .A(D6793_Y));
KC_NAND3_X1 D11960 ( .Y(D11960_Y), .C(D11954_Y), .B(D6793_Y),     .A(D6791_Y));
KC_NAND3_X1 D11959 ( .Y(D11959_Y), .C(D5480_Y), .B(D11421_Y),     .A(D5376_Y));
KC_NAND3_X1 D11904 ( .Y(D11904_Y), .C(D5479_Y), .B(D11421_Y),     .A(D5377_Y));
KC_NAND3_X1 D11566 ( .Y(D11566_Y), .C(D8331_Y), .B(D8473_Y),     .A(D5214_Y));
KC_NAND3_X1 D11565 ( .Y(D11565_Y), .C(D8331_Y), .B(D8473_Y),     .A(D5214_Y));
KC_NAND3_X1 D11564 ( .Y(D11564_Y), .C(D8331_Y), .B(D8472_Y),     .A(D5214_Y));
KC_NAND3_X1 D11563 ( .Y(D11563_Y), .C(D8331_Y), .B(D8472_Y),     .A(D5214_Y));
KC_NAND3_X1 D11379 ( .Y(D11379_Y), .C(D8331_Y), .B(D8302_Y),     .A(D5214_Y));
KC_NAND3_X1 D11377 ( .Y(D11377_Y), .C(D8331_Y), .B(D8302_Y),     .A(D5214_Y));
KC_NAND3_X1 D11305 ( .Y(D11305_Y), .C(D8331_Y), .B(D1961_Y),     .A(D5214_Y));
KC_NAND3_X1 D11154 ( .Y(D11154_Y), .C(D8331_Y), .B(D8258_Y),     .A(D5214_Y));
KC_NAND3_X1 D11153 ( .Y(D11153_Y), .C(D8331_Y), .B(D8258_Y),     .A(D5214_Y));
KC_NAND3_X1 D10989 ( .Y(D10989_Y), .C(D5480_Y), .B(D11421_Y),     .A(D5376_Y));
KC_NAND3_X1 D10988 ( .Y(D10988_Y), .C(D5479_Y), .B(D11421_Y),     .A(D5377_Y));
KC_NAND3_X1 D10987 ( .Y(D10987_Y), .C(D10514_Y), .B(D8540_Y),     .A(D6791_Y));
KC_NAND3_X1 D10986 ( .Y(D10986_Y), .C(D1143_Y), .B(D8540_Y),     .A(D6793_Y));
KC_NAND3_X1 D10984 ( .Y(D10984_Y), .C(D5479_Y), .B(D11421_Y),     .A(D5377_Y));
KC_NAND3_X1 D10983 ( .Y(D10983_Y), .C(D5480_Y), .B(D11421_Y),     .A(D5376_Y));
KC_NAND3_X1 D10982 ( .Y(D10982_Y), .C(D11421_Y), .B(D5376_Y),     .A(D5377_Y));
KC_NAND3_X1 D10937 ( .Y(D10937_Y), .C(D11421_Y), .B(D5376_Y),     .A(D5377_Y));
KC_NAND3_X1 D10862 ( .Y(D10862_Y), .C(D8331_Y), .B(D1961_Y),     .A(D5214_Y));
KC_NAND3_X1 D10771 ( .Y(D10771_Y), .C(D5403_Y), .B(D6793_Y),     .A(D6791_Y));
KC_NAND3_X1 D10768 ( .Y(D10768_Y), .C(D10514_Y), .B(D5403_Y),     .A(D6791_Y));
KC_NAND3_X1 D10764 ( .Y(D10764_Y), .C(D1143_Y), .B(D5403_Y),     .A(D6793_Y));
KC_NAND3_X1 D10763 ( .Y(D10763_Y), .C(D5480_Y), .B(D2206_Y),     .A(D5376_Y));
KC_NAND3_X1 D10762 ( .Y(D10762_Y), .C(D5479_Y), .B(D2206_Y),     .A(D5377_Y));
KC_NAND3_X1 D10761 ( .Y(D10761_Y), .C(D2206_Y), .B(D5376_Y),     .A(D5377_Y));
KC_NAND3_X1 D10487 ( .Y(D10487_Y), .C(D10464_Y), .B(D8498_Y),     .A(D10926_Y));
KC_NAND3_X1 D10486 ( .Y(D10486_Y), .C(D10514_Y), .B(D8540_Y),     .A(D6791_Y));
KC_NAND3_X1 D10485 ( .Y(D10485_Y), .C(D1143_Y), .B(D8540_Y),     .A(D6793_Y));
KC_NAND3_X1 D10483 ( .Y(D10483_Y), .C(D10451_Y), .B(D10470_Y),     .A(D8498_Y));
KC_NAND3_X1 D10479 ( .Y(D10479_Y), .C(D8540_Y), .B(D6793_Y),     .A(D6791_Y));
KC_NAND3_X1 D10478 ( .Y(D10478_Y), .C(D10452_Y), .B(D10531_Y),     .A(D8498_Y));
KC_NAND3_X1 D10473 ( .Y(D10473_Y), .C(D10447_Y), .B(D10579_Y),     .A(D8498_Y));
KC_NAND3_X1 D10410 ( .Y(D10410_Y), .C(D10466_Y), .B(D8498_Y),     .A(D10908_Y));
KC_NAND3_X1 D10409 ( .Y(D10409_Y), .C(D10460_Y), .B(D10901_Y),     .A(D8498_Y));
KC_NAND3_X1 D10154 ( .Y(D10154_Y), .C(D10161_Y), .B(D10159_Y),     .A(D10162_Y));
KC_NAND3_X1 D10055 ( .Y(D10055_Y), .C(D338_Y), .B(D9147_Y),     .A(D10059_Q));
KC_NAND3_X1 D9770 ( .Y(D9770_Y), .C(D9726_Y), .B(D9874_Y),     .A(D8499_Y));
KC_NAND3_X1 D9759 ( .Y(D9759_Y), .C(D9741_Y), .B(D10585_Y),     .A(D8498_Y));
KC_NAND3_X1 D9758 ( .Y(D9758_Y), .C(D9740_Y), .B(D10521_Y),     .A(D8498_Y));
KC_NAND3_X1 D9756 ( .Y(D9756_Y), .C(D9742_Y), .B(D9820_Y),     .A(D8499_Y));
KC_NAND3_X1 D9755 ( .Y(D9755_Y), .C(D9727_Y), .B(D9870_Y),     .A(D8499_Y));
KC_NAND3_X1 D9754 ( .Y(D9754_Y), .C(D9736_Y), .B(D9823_Y),     .A(D8499_Y));
KC_NAND3_X1 D9753 ( .Y(D9753_Y), .C(D9733_Y), .B(D10591_Y),     .A(D8499_Y));
KC_NAND3_X1 D9691 ( .Y(D9691_Y), .C(D9643_Y), .B(D10384_Y),     .A(D8498_Y));
KC_NAND3_X1 D9690 ( .Y(D9690_Y), .C(D9682_Y), .B(D10400_Y),     .A(D8498_Y));
KC_NAND3_X1 D9689 ( .Y(D9689_Y), .C(D9681_Y), .B(D9671_Y),     .A(D8498_Y));
KC_NAND3_X1 D9688 ( .Y(D9688_Y), .C(D9750_Y), .B(D10935_Y),     .A(D8498_Y));
KC_NAND3_X1 D9687 ( .Y(D9687_Y), .C(D9752_Y), .B(D9667_Y),     .A(D8498_Y));
KC_NAND3_X1 D9552 ( .Y(D9552_Y), .C(D9590_Y), .B(D2073_Y),     .A(D9394_Y));
KC_NAND3_X1 D9551 ( .Y(D9551_Y), .C(D9528_Y), .B(D9526_Y),     .A(D9575_Q));
KC_NAND3_X1 D9550 ( .Y(D9550_Y), .C(D9528_Y), .B(D9520_Y),     .A(D9575_Q));
KC_NAND3_X1 D9547 ( .Y(D9547_Y), .C(D9514_Y), .B(D9522_Y),     .A(D9513_Y));
KC_NAND3_X1 D9546 ( .Y(D9546_Y), .C(D9535_Y), .B(D1983_Y),     .A(D10300_Q));
KC_NAND3_X1 D9545 ( .Y(D9545_Y), .C(D9536_Y), .B(D9579_Q),     .A(D9544_Y));
KC_NAND3_X1 D9543 ( .Y(D9543_Y), .C(D2039_Y), .B(D9506_Y),     .A(D9576_Q));
KC_NAND3_X1 D9437 ( .Y(D9437_Y), .C(D9421_Y), .B(D9416_Y),     .A(D9439_Y));
KC_NAND3_X1 D9436 ( .Y(D9436_Y), .C(D9403_Y), .B(D9403_Y),     .A(D9395_Y));
KC_NAND3_X1 D9435 ( .Y(D9435_Y), .C(D1982_Y), .B(D9409_Y),     .A(D9407_Y));
KC_NAND3_X1 D9309 ( .Y(D9309_Y), .C(D9288_Y), .B(D9338_Y),     .A(D2002_Y));
KC_NAND3_X1 D9308 ( .Y(D9308_Y), .C(D9339_Y), .B(D9337_Y),     .A(D9167_Y));
KC_NAND3_X1 D9250 ( .Y(D9250_Y), .C(D2120_Y), .B(D2003_Y), .A(D407_Y));
KC_NAND3_X1 D9248 ( .Y(D9248_Y), .C(D7816_Y), .B(D9291_Y),     .A(D9240_Y));
KC_NAND3_X1 D9244 ( .Y(D9244_Y), .C(D9287_Y), .B(D9289_Y),     .A(D9180_Y));
KC_NAND3_X1 D8783 ( .Y(D8783_Y), .C(D8741_Y), .B(D2095_Y),     .A(D9480_Y));
KC_NAND3_X1 D8782 ( .Y(D8782_Y), .C(D8789_Y), .B(D7755_Y),     .A(D8793_Y));
KC_NAND3_X1 D8781 ( .Y(D8781_Y), .C(D9482_Y), .B(D9479_Y),     .A(D9477_Y));
KC_NAND3_X1 D8776 ( .Y(D8776_Y), .C(D8756_Y), .B(D9481_Y),     .A(D9479_Y));
KC_NAND3_X1 D8568 ( .Y(D8568_Y), .C(D8482_Y), .B(D9822_Y),     .A(D8499_Y));
KC_NAND3_X1 D8567 ( .Y(D8567_Y), .C(D8564_Y), .B(D10565_Y),     .A(D8499_Y));
KC_NAND3_X1 D8517 ( .Y(D8517_Y), .C(D8501_Y), .B(D6859_Y),     .A(D8499_Y));
KC_NAND3_X1 D8513 ( .Y(D8513_Y), .C(D8503_Y), .B(D9660_Y),     .A(D8498_Y));
KC_NAND3_X1 D8510 ( .Y(D8510_Y), .C(D8492_Y), .B(D1255_Y),     .A(D8499_Y));
KC_NAND3_X1 D8508 ( .Y(D8508_Y), .C(D8494_Y), .B(D9871_Y),     .A(D8499_Y));
KC_NAND3_X1 D8297 ( .Y(D8297_Y), .C(D7669_Y), .B(D6702_Y),     .A(D2343_Y));
KC_NAND3_X1 D8207 ( .Y(D8207_Y), .C(D8296_Y), .B(D8300_Y),     .A(D7895_Y));
KC_NAND3_X1 D8128 ( .Y(D8128_Y), .C(D7782_Y), .B(D6014_Y),     .A(D8105_Y));
KC_NAND3_X1 D8125 ( .Y(D8125_Y), .C(D8128_Y), .B(D8116_Y),     .A(D1839_Y));
KC_NAND3_X1 D8030 ( .Y(D8030_Y), .C(D8017_Y), .B(D9385_Q),     .A(D8016_Y));
KC_NAND3_X1 D7955 ( .Y(D7955_Y), .C(D7949_Y), .B(D7941_Y),     .A(D1940_Q));
KC_NAND3_X1 D7954 ( .Y(D7954_Y), .C(D7987_Y), .B(D7934_Y),     .A(D7944_Y));
KC_NAND3_X1 D7871 ( .Y(D7871_Y), .C(D1860_Y), .B(D7899_Y),     .A(D7874_Y));
KC_NAND3_X1 D7870 ( .Y(D7870_Y), .C(D7903_Y), .B(D7874_Y),     .A(D7939_Y));
KC_NAND3_X1 D7867 ( .Y(D7867_Y), .C(D7898_Y), .B(D7904_Y),     .A(D7866_Y));
KC_NAND3_X1 D7866 ( .Y(D7866_Y), .C(D7862_Y), .B(D7888_Q),     .A(D7953_Y));
KC_NAND3_X1 D7862 ( .Y(D7862_Y), .C(D1853_Y), .B(D152_Q), .A(D1940_Q));
KC_NAND3_X1 D7777 ( .Y(D7777_Y), .C(D7817_Y), .B(D461_Y), .A(D9175_Y));
KC_NAND3_X1 D7774 ( .Y(D7774_Y), .C(D458_Y), .B(D7820_Y), .A(D434_Y));
KC_NAND3_X1 D7773 ( .Y(D7773_Y), .C(D459_Y), .B(D7815_Y), .A(D7683_Y));
KC_NAND3_X1 D7700 ( .Y(D7700_Y), .C(D9269_Y), .B(D10142_Y),     .A(D12863_Y));
KC_NAND3_X1 D7699 ( .Y(D7699_Y), .C(D9164_Y), .B(D9101_Y),     .A(D7693_Y));
KC_NAND3_X1 D7698 ( .Y(D7698_Y), .C(D9164_Y), .B(D7683_Y),     .A(D7619_Y));
KC_NAND3_X1 D7644 ( .Y(D7644_Y), .C(D235_Y), .B(D8838_Y), .A(D1787_Y));
KC_NAND3_X1 D7643 ( .Y(D7643_Y), .C(D4150_Y), .B(D8838_Y), .A(D20_Y));
KC_NAND3_X1 D7457 ( .Y(D7457_Y), .C(D6038_Y), .B(D1875_Y),     .A(D7374_Y));
KC_NAND3_X1 D7452 ( .Y(D7452_Y), .C(D9_Y), .B(D7426_Y), .A(D726_Y));
KC_NAND3_X1 D7450 ( .Y(D7450_Y), .C(D7478_Q), .B(D285_Y), .A(D7452_Y));
KC_NAND3_X1 D7447 ( .Y(D7447_Y), .C(D6022_Y), .B(D5684_Y),     .A(D6001_Y));
KC_NAND3_X1 D7377 ( .Y(D7377_Y), .C(D7359_Y), .B(D268_Q), .A(D7337_Y));
KC_NAND3_X1 D7372 ( .Y(D7372_Y), .C(D7409_Q), .B(D9478_Y),     .A(D7193_Y));
KC_NAND3_X1 D7371 ( .Y(D7371_Y), .C(D7317_Y), .B(D7193_Y),     .A(D9478_Y));
KC_NAND3_X1 D7365 ( .Y(D7365_Y), .C(D7436_Y), .B(D7984_Y),     .A(D5863_Y));
KC_NAND3_X1 D7279 ( .Y(D7279_Y), .C(D7101_Y), .B(D6334_Y),     .A(D6333_Y));
KC_NAND3_X1 D7274 ( .Y(D7274_Y), .C(D7242_Y), .B(D7241_Y),     .A(D7256_Y));
KC_NAND3_X1 D7273 ( .Y(D7273_Y), .C(D6470_Y), .B(D7140_Y),     .A(D7256_Y));
KC_NAND3_X1 D7271 ( .Y(D7271_Y), .C(D8749_Y), .B(D8876_Y),     .A(D7304_Y));
KC_NAND3_X1 D7268 ( .Y(D7268_Y), .C(D8876_Y), .B(D7183_Y), .A(D209_Y));
KC_NAND3_X1 D7267 ( .Y(D7267_Y), .C(D202_Y), .B(D7175_Y), .A(D7171_Y));
KC_NAND3_X1 D7266 ( .Y(D7266_Y), .C(D7185_Y), .B(D8822_Q),     .A(D7184_Y));
KC_NAND3_X1 D7264 ( .Y(D7264_Y), .C(D7227_Y), .B(D7214_Y),     .A(D7171_Y));
KC_NAND3_X1 D7126 ( .Y(D7126_Y), .C(D7144_Q), .B(D7146_Q), .A(D192_Q));
KC_NAND3_X1 D7124 ( .Y(D7124_Y), .C(D8861_Y), .B(D192_Q), .A(D7116_Y));
KC_NAND3_X1 D7120 ( .Y(D7120_Y), .C(D7101_Y), .B(D7255_Y),     .A(D6334_Y));
KC_NAND3_X1 D7119 ( .Y(D7119_Y), .C(D7099_Y), .B(D174_Y), .A(D189_Y));
KC_NAND3_X1 D6944 ( .Y(D6944_Y), .C(D10514_Y), .B(D8540_Y),     .A(D6791_Y));
KC_NAND3_X1 D6943 ( .Y(D6943_Y), .C(D8540_Y), .B(D6793_Y),     .A(D6791_Y));
KC_NAND3_X1 D6942 ( .Y(D6942_Y), .C(D1143_Y), .B(D8540_Y),     .A(D6793_Y));
KC_NAND3_X1 D6882 ( .Y(D6882_Y), .C(D8540_Y), .B(D6808_Y),     .A(D6809_Y));
KC_NAND3_X1 D6881 ( .Y(D6881_Y), .C(D1143_Y), .B(D8540_Y),     .A(D6808_Y));
KC_NAND3_X1 D6795 ( .Y(D6795_Y), .C(D5403_Y), .B(D6808_Y),     .A(D6809_Y));
KC_NAND3_X1 D6457 ( .Y(D6457_Y), .C(D471_Y), .B(D6442_Y), .A(D5071_Y));
KC_NAND3_X1 D6164 ( .Y(D6164_Y), .C(D6151_Y), .B(D6151_Y),     .A(D6184_Y));
KC_NAND3_X1 D6061 ( .Y(D6061_Y), .C(D6060_Y), .B(D5841_Y),     .A(D5646_Y));
KC_NAND3_X1 D6060 ( .Y(D6060_Y), .C(D5831_Y), .B(D6032_Y),     .A(D6036_Y));
KC_NAND3_X1 D6057 ( .Y(D6057_Y), .C(D6061_Y), .B(D7242_Y),     .A(D4402_Y));
KC_NAND3_X1 D6054 ( .Y(D6054_Y), .C(D5986_Y), .B(D5988_Y),     .A(D5989_Y));
KC_NAND3_X1 D6048 ( .Y(D6048_Y), .C(D20_Y), .B(D5986_Y), .A(D4150_Y));
KC_NAND3_X1 D6047 ( .Y(D6047_Y), .C(D6099_Y), .B(D5988_Y),     .A(D6008_Y));
KC_NAND3_X1 D6045 ( .Y(D6045_Y), .C(D5987_Y), .B(D6002_Y),     .A(D5641_Y));
KC_NAND3_X1 D6044 ( .Y(D6044_Y), .C(D4416_Y), .B(D1713_Y), .A(D277_Y));
KC_NAND3_X1 D6043 ( .Y(D6043_Y), .C(D6099_Y), .B(D6011_Y),     .A(D5993_Y));
KC_NAND3_X1 D6040 ( .Y(D6040_Y), .C(D5958_Y), .B(D4417_Y),     .A(D4408_Y));
KC_NAND3_X1 D5918 ( .Y(D5918_Y), .C(D1592_Y), .B(D5771_Y),     .A(D5651_Y));
KC_NAND3_X1 D5912 ( .Y(D5912_Y), .C(D5840_Y), .B(D5846_Y),     .A(D7315_Y));
KC_NAND3_X1 D5909 ( .Y(D5909_Y), .C(D5908_Y), .B(D7368_Y),     .A(D7335_Y));
KC_NAND3_X1 D5907 ( .Y(D5907_Y), .C(D5925_Y), .B(D5851_Y),     .A(D5755_Y));
KC_NAND3_X1 D5905 ( .Y(D5905_Y), .C(D213_Y), .B(D5898_Y), .A(D5831_Y));
KC_NAND3_X1 D5904 ( .Y(D5904_Y), .C(D213_Y), .B(D6032_Y), .A(D5899_Y));
KC_NAND3_X1 D5793 ( .Y(D5793_Y), .C(D7092_Y), .B(D7257_Y),     .A(D5642_Y));
KC_NAND3_X1 D5792 ( .Y(D5792_Y), .C(D7242_Y), .B(D7254_Y),     .A(D7256_Y));
KC_NAND3_X1 D5789 ( .Y(D5789_Y), .C(D5744_Y), .B(D5743_Y),     .A(D1726_Y));
KC_NAND3_X1 D5788 ( .Y(D5788_Y), .C(D5744_Y), .B(D5743_Y),     .A(D5704_Y));
KC_NAND3_X1 D5783 ( .Y(D5783_Y), .C(D5885_Y), .B(D5884_Y),     .A(D1732_Y));
KC_NAND3_X1 D5775 ( .Y(D5775_Y), .C(D5774_Y), .B(D5804_Y), .A(D217_Y));
KC_NAND3_X1 D5676 ( .Y(D5676_Y), .C(D5665_Y), .B(D5686_Q),     .A(D5690_Q));
KC_NAND3_X1 D5675 ( .Y(D5675_Y), .C(D5670_Y), .B(D5664_Y),     .A(D5686_Q));
KC_NAND3_X1 D5674 ( .Y(D5674_Y), .C(D4135_Y), .B(D4216_Y),     .A(D4090_Y));
KC_NAND3_X1 D5673 ( .Y(D5673_Y), .C(D5664_Y), .B(D5666_Y),     .A(D5691_Q));
KC_NAND3_X1 D5672 ( .Y(D5672_Y), .C(D5653_Y), .B(D5664_Y),     .A(D5660_Y));
KC_NAND3_X1 D5523 ( .Y(D5523_Y), .C(D5480_Y), .B(D5432_Y),     .A(D5389_Y));
KC_NAND3_X1 D5521 ( .Y(D5521_Y), .C(D5479_Y), .B(D5432_Y),     .A(D5388_Y));
KC_NAND3_X1 D5453 ( .Y(D5453_Y), .C(D5480_Y), .B(D5432_Y),     .A(D5376_Y));
KC_NAND3_X1 D5452 ( .Y(D5452_Y), .C(D5479_Y), .B(D5432_Y),     .A(D5377_Y));
KC_NAND3_X1 D5451 ( .Y(D5451_Y), .C(D5432_Y), .B(D5376_Y),     .A(D5377_Y));
KC_NAND3_X1 D5378 ( .Y(D5378_Y), .C(D5432_Y), .B(D5389_Y),     .A(D5388_Y));
KC_NAND3_X1 D5375 ( .Y(D5375_Y), .C(D1143_Y), .B(D5403_Y),     .A(D6808_Y));
KC_NAND3_X1 D5374 ( .Y(D5374_Y), .C(D5403_Y), .B(D6808_Y),     .A(D6809_Y));
KC_NAND3_X1 D5373 ( .Y(D5373_Y), .C(D10514_Y), .B(D5403_Y),     .A(D6809_Y));
KC_NAND3_X1 D5372 ( .Y(D5372_Y), .C(D1143_Y), .B(D5403_Y),     .A(D6808_Y));
KC_NAND3_X1 D5371 ( .Y(D5371_Y), .C(D5480_Y), .B(D5432_Y),     .A(D5389_Y));
KC_NAND3_X1 D5370 ( .Y(D5370_Y), .C(D5479_Y), .B(D5432_Y),     .A(D5388_Y));
KC_NAND3_X1 D5294 ( .Y(D5294_Y), .C(D5432_Y), .B(D5389_Y),     .A(D5388_Y));
KC_NAND3_X1 D5066 ( .Y(D5066_Y), .C(D1562_Y), .B(D3509_Y),     .A(D3499_Y));
KC_NAND3_X1 D5062 ( .Y(D5062_Y), .C(D4900_Y), .B(D3498_Y),     .A(D3484_Q));
KC_NAND3_X1 D5058 ( .Y(D5058_Y), .C(D3446_Y), .B(D4877_Y),     .A(D4897_Y));
KC_NAND3_X1 D5057 ( .Y(D5057_Y), .C(D4867_Y), .B(D4875_Y),     .A(D4874_Y));
KC_NAND3_X1 D5054 ( .Y(D5054_Y), .C(D3371_Y), .B(D1565_Y),     .A(D4877_Y));
KC_NAND3_X1 D4949 ( .Y(D4949_Y), .C(D4985_Y), .B(D1567_Y),     .A(D3498_Y));
KC_NAND3_X1 D4946 ( .Y(D4946_Y), .C(D3429_Y), .B(D4926_Y),     .A(D7968_Q));
KC_NAND3_X1 D4945 ( .Y(D4945_Y), .C(D4907_Y), .B(D7966_Q),     .A(D3498_Y));
KC_NAND3_X1 D4935 ( .Y(D4935_Y), .C(D3430_Y), .B(D4891_Y),     .A(D3499_Y));
KC_NAND3_X1 D4933 ( .Y(D4933_Y), .C(D4925_Y), .B(D3416_Y),     .A(D3509_Y));
KC_NAND3_X1 D4932 ( .Y(D4932_Y), .C(D5012_Y), .B(D4891_Y), .A(D445_Q));
KC_NAND3_X1 D4789 ( .Y(D4789_Y), .C(D4614_Y), .B(D4770_Y),     .A(D3163_Y));
KC_NAND3_X1 D4788 ( .Y(D4788_Y), .C(D4811_Y), .B(D4821_Q),     .A(D4822_Q));
KC_NAND3_X1 D4787 ( .Y(D4787_Y), .C(D6329_Y), .B(D4778_Y),     .A(D4816_Y));
KC_NAND3_X1 D4783 ( .Y(D4783_Y), .C(D4806_Y), .B(D4753_Y),     .A(D4792_Y));
KC_NAND3_X1 D4706 ( .Y(D4706_Y), .C(D4575_Y), .B(D1574_Y),     .A(D4694_Y));
KC_NAND3_X1 D4701 ( .Y(D4701_Y), .C(D4699_Y), .B(D4714_Y),     .A(D4711_Y));
KC_NAND3_X1 D4617 ( .Y(D4617_Y), .C(D4606_Y), .B(D4567_Q),     .A(D1706_Y));
KC_NAND3_X1 D4614 ( .Y(D4614_Y), .C(D7984_Y), .B(D3131_Y),     .A(D4528_Y));
KC_NAND3_X1 D4612 ( .Y(D4612_Y), .C(D4604_Y), .B(D3250_Y),     .A(D3135_Y));
KC_NAND3_X1 D4524 ( .Y(D4524_Y), .C(D312_Y), .B(D1515_Q), .A(D3080_Q));
KC_NAND3_X1 D4523 ( .Y(D4523_Y), .C(D4505_Y), .B(D1576_Y), .A(D309_Y));
KC_NAND3_X1 D4522 ( .Y(D4522_Y), .C(D1577_Y), .B(D310_Y), .A(D4524_Y));
KC_NAND3_X1 D4521 ( .Y(D4521_Y), .C(D1577_Y), .B(D3018_Y),     .A(D4524_Y));
KC_NAND3_X1 D4454 ( .Y(D4454_Y), .C(D4452_Y), .B(D228_Q), .A(D5969_Y));
KC_NAND3_X1 D4453 ( .Y(D4453_Y), .C(D239_Q), .B(D4294_Y), .A(D1787_Y));
KC_NAND3_X1 D4451 ( .Y(D4451_Y), .C(D5907_Y), .B(D5985_Y),     .A(D7337_Y));
KC_NAND3_X1 D4377 ( .Y(D4377_Y), .C(D4391_Y), .B(D7280_Y),     .A(D4390_Y));
KC_NAND3_X1 D4374 ( .Y(D4374_Y), .C(D5868_Y), .B(D4338_Y),     .A(D7243_Y));
KC_NAND3_X1 D4369 ( .Y(D4369_Y), .C(D4390_Y), .B(D4330_Y),     .A(D4394_Y));
KC_NAND3_X1 D4217 ( .Y(D4217_Y), .C(D5747_Y), .B(D4180_Y),     .A(D4195_Y));
KC_NAND3_X1 D4216 ( .Y(D4216_Y), .C(D4233_Y), .B(D5752_Y),     .A(D5841_Y));
KC_NAND3_X1 D4212 ( .Y(D4212_Y), .C(D5747_Y), .B(D4156_Y),     .A(D4194_Y));
KC_NAND3_X1 D4211 ( .Y(D4211_Y), .C(D5747_Y), .B(D4163_Y),     .A(D4192_Y));
KC_NAND3_X1 D4102 ( .Y(D4102_Y), .C(D5649_Y), .B(D4094_Y),     .A(D4092_Y));
KC_NAND3_X1 D4078 ( .Y(D4078_Y), .C(D4076_Y), .B(D4035_Y),     .A(D4077_Y));
KC_NAND3_X1 D3851 ( .Y(D3851_Y), .C(D8331_Y), .B(D8309_Y), .A(D497_Y));
KC_NAND3_X1 D3850 ( .Y(D3850_Y), .C(D8331_Y), .B(D8309_Y), .A(D497_Y));
KC_NAND3_X1 D3717 ( .Y(D3717_Y), .C(D8331_Y), .B(D561_Y), .A(D5214_Y));
KC_NAND3_X1 D3716 ( .Y(D3716_Y), .C(D8331_Y), .B(D561_Y), .A(D5214_Y));
KC_NAND3_X1 D3544 ( .Y(D3544_Y), .C(D124_Q), .B(D3508_Y), .A(D3370_Y));
KC_NAND3_X1 D3465 ( .Y(D3465_Y), .C(D4926_Y), .B(D3426_Y),     .A(D3372_Q));
KC_NAND3_X1 D3460 ( .Y(D3460_Y), .C(D3371_Y), .B(D4887_Y),     .A(D3431_Y));
KC_NAND3_X1 D3453 ( .Y(D3453_Y), .C(D3538_Y), .B(D3539_Y),     .A(D4923_Y));
KC_NAND3_X1 D3452 ( .Y(D3452_Y), .C(D3576_Q), .B(D5012_Y),     .A(D3365_Y));
KC_NAND3_X1 D3351 ( .Y(D3351_Y), .C(D3208_Y), .B(D3205_Y),     .A(D3387_Q));
KC_NAND3_X1 D3350 ( .Y(D3350_Y), .C(D3318_Y), .B(D3317_Y),     .A(D3275_Y));
KC_NAND3_X1 D3347 ( .Y(D3347_Y), .C(D3384_Q), .B(D3275_Y),     .A(D3208_Y));
KC_NAND3_X1 D3338 ( .Y(D3338_Y), .C(D3306_Y), .B(D3305_Y),     .A(D3303_Y));
KC_NAND3_X1 D3248 ( .Y(D3248_Y), .C(D3219_Y), .B(D3380_Y),     .A(D3214_Y));
KC_NAND3_X1 D3245 ( .Y(D3245_Y), .C(D3215_Y), .B(D3368_Y),     .A(D3273_Y));
KC_NAND3_X1 D3244 ( .Y(D3244_Y), .C(D3290_Y), .B(D3291_Y),     .A(D3290_Y));
KC_NAND3_X1 D3243 ( .Y(D3243_Y), .C(D3322_Y), .B(D3368_Y),     .A(D3270_Y));
KC_NAND3_X1 D3163 ( .Y(D3163_Y), .C(D3129_Y), .B(D3139_Y),     .A(D1430_Y));
KC_NAND3_X1 D3162 ( .Y(D3162_Y), .C(D3121_Y), .B(D3182_Y),     .A(D3170_Y));
KC_NAND3_X1 D3157 ( .Y(D3157_Y), .C(D3163_Y), .B(D4570_Y),     .A(D3126_Y));
KC_NAND3_X1 D3156 ( .Y(D3156_Y), .C(D336_Y), .B(D3163_Y), .A(D1429_Y));
KC_NAND3_X1 D3043 ( .Y(D3043_Y), .C(D3023_Y), .B(D3084_Q),     .A(D3080_Q));
KC_NAND3_X1 D2858 ( .Y(D2858_Y), .C(D2844_Y), .B(D268_Q), .A(D2902_Q));
KC_NAND3_X1 D2778 ( .Y(D2778_Y), .C(D2747_Y), .B(D2799_Q),     .A(D2798_Q));
KC_NAND3_X1 D2775 ( .Y(D2775_Y), .C(D2741_Y), .B(D2795_Q),     .A(D2796_Q));
KC_NAND3_X1 D2564 ( .Y(D2564_Y), .C(D2547_Y), .B(D2548_Y),     .A(D14501_Y));
KC_NAND3_X1 D2503 ( .Y(D2503_Y), .C(D14132_Y), .B(D14008_Y),     .A(D14019_Y));
KC_NAND3_X1 D2455 ( .Y(D2455_Y), .C(D7670_Y), .B(D2343_Y),     .A(D12659_Y));
KC_NAND3_X1 D2447 ( .Y(D2447_Y), .C(D2396_Y), .B(D2446_Y),     .A(D13499_Y));
KC_NAND3_X1 D2446 ( .Y(D2446_Y), .C(D2401_Y), .B(D14164_Q),     .A(D12944_Y));
KC_NAND3_X1 D2140 ( .Y(D2140_Y), .C(D10458_Y), .B(D10962_Y),     .A(D8498_Y));
KC_NAND3_X1 D2139 ( .Y(D2139_Y), .C(D10459_Y), .B(D2200_Y),     .A(D8498_Y));
KC_NAND3_X1 D2054 ( .Y(D2054_Y), .C(D8749_Y), .B(D9476_Y),     .A(D9482_Y));
KC_NAND3_X1 D2053 ( .Y(D2053_Y), .C(D9481_Y), .B(D2095_Y),     .A(D8749_Y));
KC_NAND3_X1 D2045 ( .Y(D2045_Y), .C(D9217_Q), .B(D7631_Y),     .A(D9068_Y));
KC_NAND3_X1 D2043 ( .Y(D2043_Y), .C(D2000_Y), .B(D9303_Y),     .A(D9239_Y));
KC_NAND3_X1 D2042 ( .Y(D2042_Y), .C(D7669_Y), .B(D7670_Y),     .A(D7668_Y));
KC_NAND3_X1 D2041 ( .Y(D2041_Y), .C(D9536_Y), .B(D10239_Q),     .A(D8105_Y));
KC_NAND3_X1 D2038 ( .Y(D2038_Y), .C(D8424_Y), .B(D9661_Y),     .A(D8498_Y));
KC_NAND3_X1 D2033 ( .Y(D2033_Y), .C(D1832_Y), .B(D10569_Y),     .A(D8499_Y));
KC_NAND3_X1 D3 ( .Y(D3_Y), .C(D6038_Y), .B(D1874_Y), .A(D7374_Y));
KC_NAND3_X1 D1910 ( .Y(D1910_Y), .C(D8777_Y), .B(D207_Y), .A(D172_Y));
KC_NAND3_X1 D1907 ( .Y(D1907_Y), .C(D7317_Y), .B(D177_Y), .A(D7318_Y));
KC_NAND3_X1 D1904 ( .Y(D1904_Y), .C(D235_Y), .B(D1787_Y), .A(D1713_Y));
KC_NAND3_X1 D1902 ( .Y(D1902_Y), .C(D7940_Y), .B(D7832_Y),     .A(D7955_Y));
KC_NAND3_X1 D1899 ( .Y(D1899_Y), .C(D7974_Y), .B(D7921_Y), .A(D727_Y));
KC_NAND3_X1 D1897 ( .Y(D1897_Y), .C(D1915_Y), .B(D8249_Q),     .A(D8247_Q));
KC_NAND3_X1 D1892 ( .Y(D1892_Y), .C(D8504_Y), .B(D6847_Y),     .A(D8499_Y));
KC_NAND3_X1 D1749 ( .Y(D1749_Y), .C(D6043_Y), .B(D6093_Y), .A(D723_Q));
KC_NAND3_X1 D1746 ( .Y(D1746_Y), .C(D1696_Y), .B(D1695_Y),     .A(D1696_Y));
KC_NAND3_X1 D1744 ( .Y(D1744_Y), .C(D4864_Y), .B(D4926_Y),     .A(D7935_Y));
KC_NAND3_X1 D1612 ( .Y(D1612_Y), .C(D5988_Y), .B(D4235_Q), .A(D228_Q));
KC_NAND3_X1 D1607 ( .Y(D1607_Y), .C(D4589_Y), .B(D4638_Q),     .A(D4636_Q));
KC_NAND3_X1 D1606 ( .Y(D1606_Y), .C(D4581_Y), .B(D4575_Y),     .A(D4578_Y));
KC_NAND3_X1 D1599 ( .Y(D1599_Y), .C(D5479_Y), .B(D5432_Y),     .A(D5388_Y));
KC_NAND3_X1 D1598 ( .Y(D1598_Y), .C(D5480_Y), .B(D5432_Y),     .A(D5389_Y));
KC_NAND3_X1 D1597 ( .Y(D1597_Y), .C(D5432_Y), .B(D5389_Y),     .A(D5388_Y));
KC_NAND3_X1 D1458 ( .Y(D1458_Y), .C(D3144_Y), .B(D3190_Q),     .A(D3187_Q));
KC_NAND3_X1 D1450 ( .Y(D1450_Y), .C(D3576_Q), .B(D3540_Y),     .A(D3477_Y));
KC_NAND3_X1 D1445 ( .Y(D1445_Y), .C(D8331_Y), .B(D8471_Y), .A(D497_Y));
KC_NAND3_X1 D1444 ( .Y(D1444_Y), .C(D8331_Y), .B(D8471_Y), .A(D497_Y));
KC_NAND3_X1 D1108 ( .Y(D1108_Y), .C(D11421_Y), .B(D5376_Y),     .A(D5377_Y));
KC_NAND3_X1 D1107 ( .Y(D1107_Y), .C(D8540_Y), .B(D6793_Y),     .A(D6791_Y));
KC_NAND3_X1 D1104 ( .Y(D1104_Y), .C(D9744_Y), .B(D2131_Y),     .A(D8498_Y));
KC_NAND3_X1 D997 ( .Y(D997_Y), .C(D12950_Y), .B(D14239_Q),     .A(D12944_Y));
KC_NAND3_X1 D995 ( .Y(D995_Y), .C(D2372_Y), .B(D14241_Q),     .A(D12944_Y));
KC_NAND3_X1 D992 ( .Y(D992_Y), .C(D10514_Y), .B(D8540_Y), .A(D6809_Y));
KC_NAND3_X1 D991 ( .Y(D991_Y), .C(D8366_Y), .B(D10376_Y), .A(D8498_Y));
KC_NAND3_X1 D990 ( .Y(D990_Y), .C(D9645_Y), .B(D10391_Y), .A(D8498_Y));
KC_NAND3_X1 D879 ( .Y(D879_Y), .C(D15697_Y), .B(D15646_Y), .A(D88_Y));
KC_NAND3_X1 D878 ( .Y(D878_Y), .C(D14563_Y), .B(D15079_Y),     .A(D15562_Y));
KC_NAND3_X1 D875 ( .Y(D875_Y), .C(D10514_Y), .B(D5403_Y), .A(D6809_Y));
KC_NAND3_X1 D765 ( .Y(D765_Y), .C(D10775_Y), .B(D10863_Y),     .A(D10819_Y));
KC_NAND3_X1 D764 ( .Y(D764_Y), .C(D15958_Y), .B(D14665_Y),     .A(D13947_Y));
KC_NAND3_X1 D763 ( .Y(D763_Y), .C(D14026_Y), .B(D13328_Y),     .A(D12856_Q));
KC_NAND3_X1 D648 ( .Y(D648_Y), .C(D12279_Q), .B(D12729_Y), .A(D699_Q));
KC_NAND3_X1 D645 ( .Y(D645_Y), .C(D14619_Y), .B(D647_Y), .A(D14685_Q));
KC_NAND3_X1 D435 ( .Y(D435_Y), .C(D1603_Y), .B(D444_Q), .A(D4930_Y));
KC_NAND3_X1 D347 ( .Y(D347_Y), .C(D9057_Y), .B(D9147_Y), .A(D10062_Q));
KC_NAND3_X1 D346 ( .Y(D346_Y), .C(D1787_Y), .B(D235_Y), .A(D6114_Y));
KC_NAND3_X1 D314 ( .Y(D314_Y), .C(D5641_Y), .B(D6028_Y), .A(D7496_Y));
KC_NAND3_X1 D310 ( .Y(D310_Y), .C(D3016_Y), .B(D3037_Y), .A(D3080_Q));
KC_NAND3_X1 D293 ( .Y(D293_Y), .C(D4437_Y), .B(D5982_Y), .A(D286_Y));
KC_NAND3_X1 D290 ( .Y(D290_Y), .C(D4417_Y), .B(D4421_Y), .A(D4235_Q));
KC_NAND3_X1 D257 ( .Y(D257_Y), .C(D5864_Y), .B(D243_Y), .A(D5866_Y));
KC_NAND3_X1 D222 ( .Y(D222_Y), .C(D8756_Y), .B(D8760_Y), .A(D9480_Y));
KC_NAND3_X1 D219 ( .Y(D219_Y), .C(D4168_Y), .B(D5754_Y), .A(D5980_Y));
KC_XOR2_X4 D15435 ( .Y(D15435_Y), .A(D16677_Q), .B(D16693_Y));
KC_XOR2_X4 D15434 ( .Y(D15434_Y), .A(D16216_Y), .B(D16219_Y));
KC_XOR2_X4 D15330 ( .Y(D15330_Y), .A(D16205_Y), .B(D16209_Y));
KC_XOR2_X4 D15329 ( .Y(D15329_Y), .A(D15331_Y), .B(D16109_Y));
KC_XOR2_X4 D15323 ( .Y(D15323_Y), .A(D16173_Y), .B(D2674_Y));
KC_XOR2_X4 D15322 ( .Y(D15322_Y), .A(D16154_Y), .B(D16165_Y));
KC_XOR2_X4 D15319 ( .Y(D15319_Y), .A(D659_Y), .B(D16152_Y));
KC_XOR2_X4 D15316 ( .Y(D15316_Y), .A(D16098_Y), .B(D2152_Y));
KC_XOR2_X4 D15257 ( .Y(D15257_Y), .A(D15266_Y), .B(D2669_Y));
KC_XOR2_X4 D15256 ( .Y(D15256_Y), .A(D16024_Y), .B(D16074_Y));
KC_XOR2_X4 D15255 ( .Y(D15255_Y), .A(D16091_Y), .B(D16075_Y));
KC_XOR2_X4 D15254 ( .Y(D15254_Y), .A(D16076_Y), .B(D16081_Y));
KC_XOR2_X4 D15253 ( .Y(D15253_Y), .A(D16061_Y), .B(D16046_Y));
KC_XOR2_X4 D14586 ( .Y(D14586_Y), .A(D15306_Y), .B(D12637_Y));
KC_XOR2_X4 D14517 ( .Y(D14517_Y), .A(D16171_Y), .B(D15332_Y));
KC_XOR2_X4 D14515 ( .Y(D14515_Y), .A(D15456_Y), .B(D2683_Y));
KC_XOR2_X4 D14373 ( .Y(D14373_Y), .A(D15390_Y), .B(D16035_Y));
KC_XOR2_X4 D13857 ( .Y(D13857_Y), .A(D16034_Y), .B(D16019_Y));
KC_XOR2_X4 D13754 ( .Y(D13754_Y), .A(D505_Y), .B(D16021_Y));
KC_XOR2_X4 D13411 ( .Y(D13411_Y), .A(D16023_Y), .B(D16030_Y));
KC_XOR2_X4 D13170 ( .Y(D13170_Y), .A(D16036_Y), .B(D16039_Y));
KC_XOR2_X4 D12637 ( .Y(D12637_Y), .A(D16022_Y), .B(D16020_Y));
KC_XOR2_X4 D12238 ( .Y(D12238_Y), .A(D15252_Y), .B(D15251_Y));
KC_XOR2_X4 D12218 ( .Y(D12218_Y), .A(D2574_Q), .B(D13923_Y));
KC_XOR2_X4 D12214 ( .Y(D12214_Y), .A(D13866_Y), .B(D7819_Y));
KC_XOR2_X4 D12140 ( .Y(D12140_Y), .A(D541_Y), .B(D7819_Y));
KC_XOR2_X4 D11100 ( .Y(D11100_Y), .A(D1245_Y), .B(D14284_Y));
KC_XOR2_X4 D770 ( .Y(D770_Y), .A(D13862_Y), .B(D2506_Y));
KC_XOR2_X4 D10266 ( .Y(D10266_Y), .A(D13747_Y), .B(D13738_Y));
KC_XOR2_X4 D10207 ( .Y(D10207_Y), .A(D13376_Y), .B(D13320_Y));
KC_XOR2_X4 D10206 ( .Y(D10206_Y), .A(D16764_Y), .B(D529_Q));
KC_XOR2_X4 D9457 ( .Y(D9457_Y), .A(D12180_Y), .B(D7822_Y));
KC_XOR2_X4 D9379 ( .Y(D9379_Y), .A(D12226_Y), .B(D11668_Y));
KC_XOR2_X4 D9265 ( .Y(D9265_Y), .A(D9030_Y), .B(D1364_Q));
KC_XOR2_X4 D9030 ( .Y(D9030_Y), .A(D11090_Y), .B(D11091_Y));
KC_XOR2_X4 D9006 ( .Y(D9006_Y), .A(D9434_Y), .B(D9493_Q));
KC_XOR2_X4 D8946 ( .Y(D8946_Y), .A(D9376_Y), .B(D9366_Y));
KC_XOR2_X4 D8893 ( .Y(D8893_Y), .A(D7626_Y), .B(D1787_Y));
KC_XOR2_X4 D8703 ( .Y(D8703_Y), .A(D8987_Y), .B(D7549_Y));
KC_XOR2_X4 D8701 ( .Y(D8701_Y), .A(D9018_Y), .B(D2016_Y));
KC_XOR2_X4 D8237 ( .Y(D8237_Y), .A(D2025_Y), .B(D303_Q));
KC_XOR2_X4 D8050 ( .Y(D8050_Y), .A(D267_Q), .B(D8829_Y));
KC_XOR2_X4 D7882 ( .Y(D7882_Y), .A(D8727_Y), .B(D8721_Y));
KC_XOR2_X4 D7781 ( .Y(D7781_Y), .A(D8676_Y), .B(D180_Y));
KC_XOR2_X4 D7655 ( .Y(D7655_Y), .A(D8150_Q), .B(D8253_Y));
KC_XOR2_X4 D7653 ( .Y(D7653_Y), .A(D8058_Q), .B(D9377_S));
KC_XOR2_X4 D7580 ( .Y(D7580_Y), .A(D6485_Y), .B(D7861_Y));
KC_XOR2_X4 D7523 ( .Y(D7523_Y), .A(D1942_Q), .B(D4801_S));
KC_XOR2_X4 D7136 ( .Y(D7136_Y), .A(D7692_Y), .B(D6258_QN));
KC_XOR2_X4 D7135 ( .Y(D7135_Y), .A(D1863_Y), .B(D7583_QN));
KC_XOR2_X4 D7134 ( .Y(D7134_Y), .A(D7550_Y), .B(D7589_Y));
KC_XOR2_X4 D6813 ( .Y(D6813_Y), .A(D6198_Y), .B(D7489_Y));
KC_XOR2_X4 D6470 ( .Y(D6470_Y), .A(D195_Q), .B(D2055_Y));
KC_XOR2_X4 D6334 ( .Y(D6334_Y), .A(D7149_Q), .B(D7431_Y));
KC_XOR2_X4 D6333 ( .Y(D6333_Y), .A(D7151_Q), .B(D7487_Y));
KC_XOR2_X4 D6260 ( .Y(D6260_Y), .A(D1762_Y), .B(D6887_S));
KC_XOR2_X4 D6259 ( .Y(D6259_Y), .A(D6451_Y), .B(D6469_Y));
KC_XOR2_X4 D6176 ( .Y(D6176_Y), .A(D6319_Y), .B(D6297_Y));
KC_XOR2_X4 D6175 ( .Y(D6175_Y), .A(D6130_Y), .B(D6232_Y));
KC_XOR2_X4 D6173 ( .Y(D6173_Y), .A(D6230_Y), .B(D6223_Y));
KC_XOR2_X4 D6172 ( .Y(D6172_Y), .A(D6166_Y), .B(D6160_Y));
KC_XOR2_X4 D6117 ( .Y(D6117_Y), .A(D6253_Y), .B(D6184_Y));
KC_XOR2_X4 D5930 ( .Y(D5930_Y), .A(D6140_Y), .B(D6203_Y));
KC_XOR2_X4 D4807 ( .Y(D4807_Y), .A(D6158_Y), .B(D6307_Y));
KC_XOR2_X4 D4804 ( .Y(D4804_Y), .A(D6127_Y), .B(D6142_Y));
KC_XOR2_X4 D4721 ( .Y(D4721_Y), .A(D7331_Y), .B(D7330_Y));
KC_XOR2_X4 D4720 ( .Y(D4720_Y), .A(D3355_Y), .B(D7623_Y));
KC_XOR2_X4 D4550 ( .Y(D4550_Y), .A(D1654_Q), .B(D4857_Y));
KC_XOR2_X4 D4549 ( .Y(D4549_Y), .A(D4661_Y), .B(D4665_Y));
KC_XOR2_X4 D4468 ( .Y(D4468_Y), .A(D4569_Q), .B(D4554_Y));
KC_XOR2_X4 D4467 ( .Y(D4467_Y), .A(D43_Y), .B(D4556_Q));
KC_XOR2_X4 D4389 ( .Y(D4389_Y), .A(D4309_Y), .B(D4450_Y));
KC_XOR2_X4 D4116 ( .Y(D4116_Y), .A(D4487_Q), .B(D1580_Y));
KC_XOR2_X4 D4115 ( .Y(D4115_Y), .A(D2956_Y), .B(D255_Y));
KC_XOR2_X4 D4111 ( .Y(D4111_Y), .A(D5678_Y), .B(D4106_Y));
KC_XOR2_X4 D3573 ( .Y(D3573_Y), .A(D4118_Q), .B(D4144_Y));
KC_XOR2_X4 D3572 ( .Y(D3572_Y), .A(D8313_Q), .B(D4151_Y));
KC_XOR2_X4 D3571 ( .Y(D3571_Y), .A(D4882_Y), .B(D3552_Y));
KC_XOR2_X4 D3370 ( .Y(D3370_Y), .A(D3543_Y), .B(D3504_Y));
KC_XOR2_X4 D3364 ( .Y(D3364_Y), .A(D3481_Q), .B(D3586_Y));
KC_XOR2_X4 D3275 ( .Y(D3275_Y), .A(D3326_Y), .B(D3287_Y));
KC_XOR2_X4 D3067 ( .Y(D3067_Y), .A(D1527_Q), .B(D4966_Y));
KC_XOR2_X4 D2995 ( .Y(D2995_Y), .A(D3267_Y), .B(D6174_Y));
KC_XOR2_X4 D2948 ( .Y(D2948_Y), .A(D4616_Y), .B(D4525_Y));
KC_XOR2_X4 D2878 ( .Y(D2878_Y), .A(D271_Y), .B(D304_Q));
KC_XOR2_X4 D2792 ( .Y(D2792_Y), .A(D2877_Y), .B(D2889_Q));
KC_XOR2_X4 D2672 ( .Y(D2672_Y), .A(D2785_Y), .B(D2800_Q));
KC_XOR2_X4 D2669 ( .Y(D2669_Y), .A(D16031_Y), .B(D2670_Y));
KC_XOR2_X4 D2152 ( .Y(D2152_Y), .A(D16026_Y), .B(D16032_Y));
KC_XOR2_X4 D1921 ( .Y(D1921_Y), .A(D8670_Y), .B(D10064_Y));
KC_XOR2_X4 D1920 ( .Y(D1920_Y), .A(D8034_Y), .B(D7980_Y));
KC_XOR2_X4 D1770 ( .Y(D1770_Y), .A(D105_Y), .B(D7617_Y));
KC_XOR2_X4 D1008 ( .Y(D1008_Y), .A(D6308_Y), .B(D1747_Y));
KC_XOR2_X4 D781 ( .Y(D781_Y), .A(D8456_Y), .B(D6889_Y));
KC_XOR2_X4 D779 ( .Y(D779_Y), .A(D10775_Y), .B(D10864_Y));
KC_XOR2_X4 D616 ( .Y(D616_Y), .A(D765_Y), .B(D16760_Co));
KC_XOR2_X4 D584 ( .Y(D584_Y), .A(D16038_Y), .B(D16027_Y));
KC_XOR2_X4 D508 ( .Y(D508_Y), .A(D528_Y), .B(D2637_Y));
KC_XOR2_X4 D504 ( .Y(D504_Y), .A(D12239_Y), .B(D11624_Y));
KC_XOR2_X4 D381 ( .Y(D381_Y), .A(D4740_Y), .B(D4730_Y));
KC_XOR2_X4 D378 ( .Y(D378_Y), .A(D370_Y), .B(D7627_Y));
KC_XOR2_X4 D323 ( .Y(D323_Y), .A(D4555_Q), .B(D3033_Y));
KC_XOR2_X4 D321 ( .Y(D321_Y), .A(D3092_Y), .B(D4562_Q));
KC_XOR2_X4 D190 ( .Y(D190_Y), .A(D7142_Y), .B(D7133_Y));
KC_BUF_X7 D16745 ( .Y(D16745_Y), .A(D4085_Y));
KC_BUF_X7 D16744 ( .Y(D16744_Y), .A(D8715_Y));
KC_BUF_X7 D16743 ( .Y(D16743_Y), .A(D12267_Y));
KC_BUF_X7 D13204 ( .Y(D13204_Y), .A(D13273_Q));
KC_BUF_X7 D13172 ( .Y(D13172_Y), .A(D535_Y));
KC_BUF_X7 D12655 ( .Y(D12655_Y), .A(D10145_Q));
KC_BUF_X7 D12654 ( .Y(D12654_Y), .A(D9362_Y));
KC_BUF_X7 D12280 ( .Y(D12280_Y), .A(D9360_Y));
KC_BUF_X7 D10660 ( .Y(D10660_Y), .A(D10132_Y));
KC_BUF_X7 D10373 ( .Y(D10373_Y), .A(D10372_Y));
KC_BUF_X7 D10164 ( .Y(D10164_Y), .A(D2167_Q));
KC_BUF_X7 D10163 ( .Y(D10163_Y), .A(D9227_Q));
KC_BUF_X7 D10149 ( .Y(D10149_Y), .A(D9217_Q));
KC_BUF_X7 D10148 ( .Y(D10148_Y), .A(D9279_Q));
KC_BUF_X7 D9945 ( .Y(D9945_Y), .A(D9977_Y));
KC_BUF_X7 D9944 ( .Y(D9944_Y), .A(D9977_Y));
KC_BUF_X7 D9943 ( .Y(D9943_Y), .A(D9935_Y));
KC_BUF_X7 D9942 ( .Y(D9942_Y), .A(D9942_A));
KC_BUF_X7 D9358 ( .Y(D9358_Y), .A(D9360_Y));
KC_BUF_X7 D8715 ( .Y(D8715_Y), .A(D8790_Y));
KC_BUF_X7 D8714 ( .Y(D8714_Y), .A(D8692_Y));
KC_BUF_X7 D8713 ( .Y(D8713_Y), .A(D9003_Y));
KC_BUF_X7 D7795 ( .Y(D7795_Y), .A(D9358_Y));
KC_BUF_X7 D4086 ( .Y(D4086_Y), .A(D2728_Y));
KC_BUF_X7 D4085 ( .Y(D4085_Y), .A(D16743_Y));
KC_BUF_X7 D2728 ( .Y(D2728_Y), .A(D4535_Y));
KC_BUF_X7 D2727 ( .Y(D2727_Y), .A(D8714_Y));
KC_BUF_X7 D2470 ( .Y(D2470_Y), .A(D13207_Q));
KC_BUF_X7 D453 ( .Y(D453_Y), .A(D10147_Q));
KC_BUF_X7 D196 ( .Y(D196_Y), .A(D9000_Y));
KC_NAND2B_X1 D16656 ( .Y(D16656_Y), .AN(D1320_Q), .B(D16681_Q));
KC_NAND2B_X1 D16604 ( .Y(D16604_Y), .AN(D1396_Q), .B(D16599_Q));
KC_NAND2B_X1 D16108 ( .Y(D16108_Y), .AN(D16106_Y), .B(D16104_Y));
KC_NAND2B_X1 D15740 ( .Y(D15740_Y), .AN(D15795_Q), .B(D145_Q));
KC_NAND2B_X1 D15498 ( .Y(D15498_Y), .AN(D16272_Y), .B(D15500_Y));
KC_NAND2B_X1 D15396 ( .Y(D15396_Y), .AN(D15267_Y), .B(D2589_Y));
KC_NAND2B_X1 D15268 ( .Y(D15268_Y), .AN(D15289_Y), .B(D15272_Y));
KC_NAND2B_X1 D14852 ( .Y(D14852_Y), .AN(D14094_Q), .B(D14725_Y));
KC_NAND2B_X1 D14730 ( .Y(D14730_Y), .AN(D16272_Y), .B(D15505_Y));
KC_NAND2B_X1 D14644 ( .Y(D14644_Y), .AN(D14635_Y), .B(D14641_Y));
KC_NAND2B_X1 D14632 ( .Y(D14632_Y), .AN(D15499_Y), .B(D14673_Y));
KC_NAND2B_X1 D14544 ( .Y(D14544_Y), .AN(D2512_Y), .B(D14556_Y));
KC_NAND2B_X1 D14536 ( .Y(D14536_Y), .AN(D14736_Y), .B(D14802_Y));
KC_NAND2B_X1 D14282 ( .Y(D14282_Y), .AN(D2435_Y), .B(D13419_Y));
KC_NAND2B_X1 D14277 ( .Y(D14277_Y), .AN(D14295_Y), .B(D14275_Y));
KC_NAND2B_X1 D14045 ( .Y(D14045_Y), .AN(D13973_Y), .B(D13975_Y));
KC_NAND2B_X1 D13725 ( .Y(D13725_Y), .AN(D13738_Y), .B(D13752_Y));
KC_NAND2B_X1 D13724 ( .Y(D13724_Y), .AN(D13718_Y), .B(D13723_Y));
KC_NAND2B_X1 D13641 ( .Y(D13641_Y), .AN(D2438_Y), .B(D13419_Y));
KC_NAND2B_X1 D13462 ( .Y(D13462_Y), .AN(D2432_Y), .B(D10216_Y));
KC_NAND2B_X1 D13340 ( .Y(D13340_Y), .AN(D13369_Y), .B(D13352_Y));
KC_NAND2B_X1 D13222 ( .Y(D13222_Y), .AN(D13340_Y), .B(D14785_Y));
KC_NAND2B_X1 D12955 ( .Y(D12955_Y), .AN(D12931_Y), .B(D12995_Q));
KC_NAND2B_X1 D12705 ( .Y(D12705_Y), .AN(D699_Q), .B(D12729_Y));
KC_NAND2B_X1 D12241 ( .Y(D12241_Y), .AN(D12195_Y), .B(D12212_Y));
KC_NAND2B_X1 D10100 ( .Y(D10100_Y), .AN(D10108_Q), .B(D9148_Q));
KC_NAND2B_X1 D9523 ( .Y(D9523_Y), .AN(D9590_Y), .B(D9519_Y));
KC_NAND2B_X1 D9497 ( .Y(D9497_Y), .AN(D9542_Y), .B(D9540_Y));
KC_NAND2B_X1 D9496 ( .Y(D9496_Y), .AN(D10241_Y), .B(D9503_Y));
KC_NAND2B_X1 D9409 ( .Y(D9409_Y), .AN(D9551_Y), .B(D8079_Y));
KC_NAND2B_X1 D9367 ( .Y(D9367_Y), .AN(D8056_Y), .B(D9794_Y));
KC_NAND2B_X1 D9238 ( .Y(D9238_Y), .AN(D70_Y), .B(D9101_Y));
KC_NAND2B_X1 D9176 ( .Y(D9176_Y), .AN(D9179_Y), .B(D9180_Y));
KC_NAND2B_X1 D9116 ( .Y(D9116_Y), .AN(D9117_Y), .B(D2122_Y));
KC_NAND2B_X1 D9103 ( .Y(D9103_Y), .AN(D9112_Y), .B(D2122_Y));
KC_NAND2B_X1 D8866 ( .Y(D8866_Y), .AN(D8895_Q), .B(D8869_Y));
KC_NAND2B_X1 D8771 ( .Y(D8771_Y), .AN(D8664_Y), .B(D8761_Y));
KC_NAND2B_X1 D8770 ( .Y(D8770_Y), .AN(D8745_Y), .B(D8761_Y));
KC_NAND2B_X1 D8678 ( .Y(D8678_Y), .AN(D8672_Y), .B(D8718_Y));
KC_NAND2B_X1 D8672 ( .Y(D8672_Y), .AN(D2056_Y), .B(D2030_Y));
KC_NAND2B_X1 D8371 ( .Y(D8371_Y), .AN(D6889_Y), .B(D11024_Y));
KC_NAND2B_X1 D8295 ( .Y(D8295_Y), .AN(D8326_Y), .B(D7895_Y));
KC_NAND2B_X1 D8294 ( .Y(D8294_Y), .AN(D6773_Y), .B(D8171_Y));
KC_NAND2B_X1 D8020 ( .Y(D8020_Y), .AN(D8212_Y), .B(D8017_Y));
KC_NAND2B_X1 D7928 ( .Y(D7928_Y), .AN(D7830_Y), .B(D7829_Y));
KC_NAND2B_X1 D7859 ( .Y(D7859_Y), .AN(D7890_Q), .B(D7855_Y));
KC_NAND2B_X1 D7772 ( .Y(D7772_Y), .AN(D6345_Q), .B(D6291_Y));
KC_NAND2B_X1 D7559 ( .Y(D7559_Y), .AN(D7574_Y), .B(D7612_Y));
KC_NAND2B_X1 D7507 ( .Y(D7507_Y), .AN(D5826_Y), .B(D7532_Y));
KC_NAND2B_X1 D7431 ( .Y(D7431_Y), .AN(D7483_Y), .B(D7463_Y));
KC_NAND2B_X1 D7319 ( .Y(D7319_Y), .AN(D8050_Y), .B(D149_Q));
KC_NAND2B_X1 D7240 ( .Y(D7240_Y), .AN(D8772_Y), .B(D7176_Y));
KC_NAND2B_X1 D7113 ( .Y(D7113_Y), .AN(D5682_Y), .B(D7125_Y));
KC_NAND2B_X1 D6784 ( .Y(D6784_Y), .AN(D5214_Y), .B(D6800_Y));
KC_NAND2B_X1 D6439 ( .Y(D6439_Y), .AN(D6479_Y), .B(D6435_Y));
KC_NAND2B_X1 D6419 ( .Y(D6419_Y), .AN(D6513_Y), .B(D6473_Q));
KC_NAND2B_X1 D6300 ( .Y(D6300_Y), .AN(D6322_Y), .B(D6338_Y));
KC_NAND2B_X1 D6299 ( .Y(D6299_Y), .AN(D6350_Q), .B(D6291_Y));
KC_NAND2B_X1 D6295 ( .Y(D6295_Y), .AN(D6340_Y), .B(D428_Y));
KC_NAND2B_X1 D6294 ( .Y(D6294_Y), .AN(D6356_Y), .B(D6312_Y));
KC_NAND2B_X1 D6293 ( .Y(D6293_Y), .AN(D6357_Q), .B(D6291_Y));
KC_NAND2B_X1 D6292 ( .Y(D6292_Y), .AN(D7741_Q), .B(D6291_Y));
KC_NAND2B_X1 D6222 ( .Y(D6222_Y), .AN(D384_Q), .B(D6291_Y));
KC_NAND2B_X1 D6219 ( .Y(D6219_Y), .AN(D6280_Y), .B(D6247_Y));
KC_NAND2B_X1 D6214 ( .Y(D6214_Y), .AN(D364_Q), .B(D6291_Y));
KC_NAND2B_X1 D6213 ( .Y(D6213_Y), .AN(D6351_Q), .B(D6291_Y));
KC_NAND2B_X1 D6150 ( .Y(D6150_Y), .AN(D395_Q), .B(D6291_Y));
KC_NAND2B_X1 D6027 ( .Y(D6027_Y), .AN(D6054_Y), .B(D5871_Y));
KC_NAND2B_X1 D5868 ( .Y(D5868_Y), .AN(D5999_Y), .B(D5848_Y));
KC_NAND2B_X1 D5858 ( .Y(D5858_Y), .AN(D5849_Y), .B(D5927_Y));
KC_NAND2B_X1 D5717 ( .Y(D5717_Y), .AN(D7195_Y), .B(D5761_Y));
KC_NAND2B_X1 D5656 ( .Y(D5656_Y), .AN(D5654_Y), .B(D5653_Y));
KC_NAND2B_X1 D5045 ( .Y(D5045_Y), .AN(D4893_Y), .B(D1562_Y));
KC_NAND2B_X1 D4763 ( .Y(D4763_Y), .AN(D7764_Y), .B(D7766_Y));
KC_NAND2B_X1 D4686 ( .Y(D4686_Y), .AN(D1606_Y), .B(D4737_Y));
KC_NAND2B_X1 D4685 ( .Y(D4685_Y), .AN(D4690_Y), .B(D4574_Y));
KC_NAND2B_X1 D4669 ( .Y(D4669_Y), .AN(D1622_Y), .B(D4668_Y));
KC_NAND2B_X1 D4668 ( .Y(D4668_Y), .AN(D4619_Y), .B(D3243_Y));
KC_NAND2B_X1 D4573 ( .Y(D4573_Y), .AN(D7787_Y), .B(D4576_Y));
KC_NAND2B_X1 D4519 ( .Y(D4519_Y), .AN(D4517_Y), .B(D1593_Y));
KC_NAND2B_X1 D4512 ( .Y(D4512_Y), .AN(D323_Y), .B(D6291_Y));
KC_NAND2B_X1 D4511 ( .Y(D4511_Y), .AN(D4561_Q), .B(D6291_Y));
KC_NAND2B_X1 D4510 ( .Y(D4510_Y), .AN(D321_Y), .B(D6291_Y));
KC_NAND2B_X1 D4507 ( .Y(D4507_Y), .AN(D328_Q), .B(D6291_Y));
KC_NAND2B_X1 D4422 ( .Y(D4422_Y), .AN(D6096_Y), .B(D4408_Y));
KC_NAND2B_X1 D4341 ( .Y(D4341_Y), .AN(D4335_Y), .B(D4374_Y));
KC_NAND2B_X1 D4329 ( .Y(D4329_Y), .AN(D4298_Y), .B(D7243_Y));
KC_NAND2B_X1 D4285 ( .Y(D4285_Y), .AN(D7316_Y), .B(D4414_Y));
KC_NAND2B_X1 D4206 ( .Y(D4206_Y), .AN(D4222_Y), .B(D4202_Y));
KC_NAND2B_X1 D4174 ( .Y(D4174_Y), .AN(D1751_Y), .B(D213_Y));
KC_NAND2B_X1 D4091 ( .Y(D4091_Y), .AN(D2716_Y), .B(D4547_Y));
KC_NAND2B_X1 D3833 ( .Y(D3833_Y), .AN(D3863_Y), .B(D3848_Y));
KC_NAND2B_X1 D3327 ( .Y(D3327_Y), .AN(D3362_Y), .B(D3331_Y));
KC_NAND2B_X1 D3313 ( .Y(D3313_Y), .AN(D3353_Y), .B(D3341_Y));
KC_NAND2B_X1 D3225 ( .Y(D3225_Y), .AN(D3350_Y), .B(D3247_Y));
KC_NAND2B_X1 D3034 ( .Y(D3034_Y), .AN(D316_Y), .B(D32_Y));
KC_NAND2B_X1 D3017 ( .Y(D3017_Y), .AN(D3027_Y), .B(D3019_Y));
KC_NAND2B_X1 D2937 ( .Y(D2937_Y), .AN(D2823_Y), .B(D2854_Y));
KC_NAND2B_X1 D2911 ( .Y(D2911_Y), .AN(D2989_Y), .B(D2991_Y));
KC_NAND2B_X1 D2742 ( .Y(D2742_Y), .AN(D2771_Y), .B(D2773_Y));
KC_NAND2B_X1 D2410 ( .Y(D2410_Y), .AN(D11228_Y), .B(D13236_Y));
KC_NAND2B_X1 D2135 ( .Y(D2135_Y), .AN(D10304_Q), .B(D98_Y));
KC_NAND2B_X1 D2120 ( .Y(D2120_Y), .AN(D9193_Y), .B(D10105_Y));
KC_NAND2B_X1 D1977 ( .Y(D1977_Y), .AN(D2030_Y), .B(D8698_Y));
KC_NAND2B_X1 D1861 ( .Y(D1861_Y), .AN(D167_Q), .B(D6291_Y));
KC_NAND2B_X1 D1860 ( .Y(D1860_Y), .AN(D7925_Y), .B(D7963_Y));
KC_NAND2B_X1 D1705 ( .Y(D1705_Y), .AN(D1766_Y), .B(D1790_Y));
KC_NAND2B_X1 D1694 ( .Y(D1694_Y), .AN(D6473_Q), .B(D6513_Y));
KC_NAND2B_X1 D1579 ( .Y(D1579_Y), .AN(D1667_Y), .B(D1667_Y));
KC_NAND2B_X1 D1578 ( .Y(D1578_Y), .AN(D6150_Y), .B(D6408_Y));
KC_NAND2B_X1 D468 ( .Y(D468_Y), .AN(D4982_Y), .B(D5093_Y));
KC_NAND2B_X1 D401 ( .Y(D401_Y), .AN(D418_Q), .B(D6291_Y));
KC_NAND2B_X1 D368 ( .Y(D368_Y), .AN(D9148_Q), .B(D10108_Q));
KC_NAND2B_X1 D182 ( .Y(D182_Y), .AN(D8708_Y), .B(D7114_Y));
KC_NAND2B_X1 D180 ( .Y(D180_Y), .AN(D9931_Y), .B(D9932_Y));
KC_NAND2B_X1 D179 ( .Y(D179_Y), .AN(D5659_Y), .B(D5667_Y));
KC_OAI22BB_X1 D14867 ( .Y(D14867_Y), .D(D14854_Y), .B(D15003_Y),     .C(D8998_Y), .A(D15562_Y));
KC_OAI22BB_X1 D14293 ( .Y(D14293_Y), .D(D14295_Y), .B(D14295_Y),     .C(D14204_Y), .A(D14294_Y));
KC_OAI22BB_X1 D13972 ( .Y(D13972_Y), .D(D14665_Y), .B(D14005_Y),     .C(D13220_Y), .A(D13939_Y));
KC_OAI22BB_X1 D12904 ( .Y(D12904_Y), .D(D12748_Q), .B(D12886_Y),     .C(D12951_Y), .A(D961_Y));
KC_OAI22BB_X1 D12834 ( .Y(D12834_Y), .D(D12314_Y), .B(D12794_Y),     .C(D12855_Q), .A(D12849_Q));
KC_OAI22BB_X1 D12396 ( .Y(D12396_Y), .D(D12888_Y), .B(D12414_Q),     .C(D12318_Y), .A(D12312_Y));
KC_OAI22BB_X1 D12395 ( .Y(D12395_Y), .D(D12888_Y), .B(D12415_Q),     .C(D2327_Y), .A(D2325_Y));
KC_OAI22BB_X1 D12394 ( .Y(D12394_Y), .D(D12770_Y), .B(D12418_Q),     .C(D12318_Y), .A(D12312_Y));
KC_OAI22BB_X1 D12393 ( .Y(D12393_Y), .D(D12770_Y), .B(D12419_Q),     .C(D2327_Y), .A(D2325_Y));
KC_OAI22BB_X1 D12333 ( .Y(D12333_Y), .D(D12771_Y), .B(D12348_Q),     .C(D12318_Y), .A(D12312_Y));
KC_OAI22BB_X1 D12332 ( .Y(D12332_Y), .D(D12888_Y), .B(D12340_Q),     .C(D2328_Y), .A(D2326_Y));
KC_OAI22BB_X1 D12331 ( .Y(D12331_Y), .D(D12869_Y), .B(D2355_Q),     .C(D2327_Y), .A(D2325_Y));
KC_OAI22BB_X1 D12330 ( .Y(D12330_Y), .D(D12869_Y), .B(D12367_Q),     .C(D2328_Y), .A(D2326_Y));
KC_OAI22BB_X1 D12329 ( .Y(D12329_Y), .D(D12869_Y), .B(D12343_Q),     .C(D12318_Y), .A(D12312_Y));
KC_OAI22BB_X1 D12039 ( .Y(D12039_Y), .D(D8461_Y), .B(D12040_Y),     .C(D6406_Y), .A(D8430_Y));
KC_OAI22BB_X1 D12038 ( .Y(D12038_Y), .D(D8461_Y), .B(D12034_Y),     .C(D10192_Y), .A(D8430_Y));
KC_OAI22BB_X1 D12036 ( .Y(D12036_Y), .D(D8461_Y), .B(D1195_Y),     .C(D1964_Y), .A(D8430_Y));
KC_OAI22BB_X1 D12035 ( .Y(D12035_Y), .D(D8461_Y), .B(D12037_Y),     .C(D463_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11853 ( .Y(D11853_Y), .D(D8464_Y), .B(D11845_Y),     .C(D813_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11850 ( .Y(D11850_Y), .D(D8464_Y), .B(D890_Y),     .C(D1814_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11844 ( .Y(D11844_Y), .D(D8464_Y), .B(D11319_Y),     .C(D6410_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11843 ( .Y(D11843_Y), .D(D8464_Y), .B(D11320_Y),     .C(D10358_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11782 ( .Y(D11782_Y), .D(D8470_Y), .B(D11249_Y),     .C(D6410_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11781 ( .Y(D11781_Y), .D(D8470_Y), .B(D11780_Y),     .C(D8336_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11777 ( .Y(D11777_Y), .D(D8470_Y), .B(D11240_Y),     .C(D813_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11532 ( .Y(D11532_Y), .D(D8461_Y), .B(D11530_Y),     .C(D8336_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11531 ( .Y(D11531_Y), .D(D8461_Y), .B(D11528_Y),     .C(D6405_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11478 ( .Y(D11478_Y), .D(D8464_Y), .B(D2237_Y),     .C(D6407_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11458 ( .Y(D11458_Y), .D(D8461_Y), .B(D11527_Y),     .C(D813_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11456 ( .Y(D11456_Y), .D(D8464_Y), .B(D11448_Y),     .C(D462_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11455 ( .Y(D11455_Y), .D(D8464_Y), .B(D11457_Y),     .C(D10192_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11451 ( .Y(D11451_Y), .D(D8464_Y), .B(D11452_Y),     .C(D10191_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11449 ( .Y(D11449_Y), .D(D8464_Y), .B(D11450_Y),     .C(D463_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11447 ( .Y(D11447_Y), .D(D8461_Y), .B(D11463_Y),     .C(D1814_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11446 ( .Y(D11446_Y), .D(D8461_Y), .B(D11460_Y),     .C(D9617_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11445 ( .Y(D11445_Y), .D(D8461_Y), .B(D11462_Y),     .C(D1813_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11444 ( .Y(D11444_Y), .D(D8461_Y), .B(D11459_Y),     .C(D464_Y), .A(D8430_Y));
KC_OAI22BB_X1 D11317 ( .Y(D11317_Y), .D(D8464_Y), .B(D11318_Y),     .C(D6406_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11248 ( .Y(D11248_Y), .D(D8470_Y), .B(D11250_Y),     .C(D6406_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11247 ( .Y(D11247_Y), .D(D8470_Y), .B(D11251_Y),     .C(D1813_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11244 ( .Y(D11244_Y), .D(D8470_Y), .B(D11245_Y),     .C(D10191_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11243 ( .Y(D11243_Y), .D(D8470_Y), .B(D772_Y),     .C(D463_Y), .A(D10788_Y));
KC_OAI22BB_X1 D11241 ( .Y(D11241_Y), .D(D8470_Y), .B(D10780_Y),     .C(D10192_Y), .A(D10788_Y));
KC_OAI22BB_X1 D10869 ( .Y(D10869_Y), .D(D8470_Y), .B(D2212_Y),     .C(D6405_Y), .A(D8431_Y));
KC_OAI22BB_X1 D10785 ( .Y(D10785_Y), .D(D8470_Y), .B(D10779_Y),     .C(D462_Y), .A(D8013_Y));
KC_OAI22BB_X1 D10782 ( .Y(D10782_Y), .D(D8470_Y), .B(D10777_Y),     .C(D1964_Y), .A(D8013_Y));
KC_OAI22BB_X1 D10781 ( .Y(D10781_Y), .D(D8470_Y), .B(D10778_Y),     .C(D6407_Y), .A(D10788_Y));
KC_OAI22BB_X1 D10506 ( .Y(D10506_Y), .D(D813_Y), .B(D10456_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10504 ( .Y(D10504_Y), .D(D8336_Y), .B(D10462_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10501 ( .Y(D10501_Y), .D(D10358_Y), .B(D10463_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10500 ( .Y(D10500_Y), .D(D10358_Y), .B(D10450_Y),     .C(D8370_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10499 ( .Y(D10499_Y), .D(D1814_Y), .B(D10520_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10497 ( .Y(D10497_Y), .D(D8336_Y), .B(D10448_Y),     .C(D8370_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10495 ( .Y(D10495_Y), .D(D6410_Y), .B(D10457_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10493 ( .Y(D10493_Y), .D(D8370_Y), .B(D10449_Y),     .C(D9617_Y), .A(D8533_Y));
KC_OAI22BB_X1 D10413 ( .Y(D10413_Y), .D(D8464_Y), .B(D8405_Y),     .C(D8336_Y), .A(D8455_Y));
KC_OAI22BB_X1 D10093 ( .Y(D10093_Y), .D(D10082_Y), .B(D12176_Y),     .C(D9943_Y), .A(D10078_Y));
KC_OAI22BB_X1 D9831 ( .Y(D9831_Y), .D(D8370_Y), .B(D9732_Y),     .C(D6405_Y), .A(D8533_Y));
KC_OAI22BB_X1 D9798 ( .Y(D9798_Y), .D(D8370_Y), .B(D9731_Y),     .C(D1814_Y), .A(D8533_Y));
KC_OAI22BB_X1 D9779 ( .Y(D9779_Y), .D(D462_Y), .B(D9747_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D9778 ( .Y(D9778_Y), .D(D8370_Y), .B(D9730_Y),     .C(D6407_Y), .A(D8533_Y));
KC_OAI22BB_X1 D9776 ( .Y(D9776_Y), .D(D464_Y), .B(D9745_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D9775 ( .Y(D9775_Y), .D(D6406_Y), .B(D9749_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D9774 ( .Y(D9774_Y), .D(D463_Y), .B(D9748_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D9773 ( .Y(D9773_Y), .D(D1813_Y), .B(D9751_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D9772 ( .Y(D9772_Y), .D(D8370_Y), .B(D9729_Y),     .C(D1964_Y), .A(D8533_Y));
KC_OAI22BB_X1 D9771 ( .Y(D9771_Y), .D(D8370_Y), .B(D9734_Y),     .C(D462_Y), .A(D8533_Y));
KC_OAI22BB_X1 D9694 ( .Y(D9694_Y), .D(D6407_Y), .B(D1980_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D9693 ( .Y(D9693_Y), .D(D1964_Y), .B(D65_Y), .C(D1836_Y),     .A(D8533_Y));
KC_OAI22BB_X1 D9692 ( .Y(D9692_Y), .D(D6405_Y), .B(D1981_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D9258 ( .Y(D9258_Y), .D(D9249_Y), .B(D9200_Y),     .C(D7626_Y), .A(D9242_Y));
KC_OAI22BB_X1 D9132 ( .Y(D9132_Y), .D(D2099_Y), .B(D5966_Y),     .C(D8971_Y), .A(D8711_Q));
KC_OAI22BB_X1 D9131 ( .Y(D9131_Y), .D(D2099_Y), .B(D5966_Y),     .C(D9014_Y), .A(D10109_Q));
KC_OAI22BB_X1 D8999 ( .Y(D8999_Y), .D(D9012_Y), .B(D9067_Y),     .C(D8980_Y), .A(D7430_Y));
KC_OAI22BB_X1 D8802 ( .Y(D8802_Y), .D(D8764_Y), .B(D8835_Q),     .C(D211_Y), .A(D215_Y));
KC_OAI22BB_X1 D8800 ( .Y(D8800_Y), .D(D8764_Y), .B(D8836_Q),     .C(D8758_Y), .A(D215_Y));
KC_OAI22BB_X1 D8687 ( .Y(D8687_Y), .D(D8722_Y), .B(D8732_Y),     .C(D2098_Y), .A(D8665_Y));
KC_OAI22BB_X1 D8575 ( .Y(D8575_Y), .D(D8378_Y), .B(D8582_Y),     .C(D464_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8574 ( .Y(D8574_Y), .D(D8370_Y), .B(D8563_Y),     .C(D10191_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8531 ( .Y(D8531_Y), .D(D8370_Y), .B(D8495_Y),     .C(D464_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8530 ( .Y(D8530_Y), .D(D8378_Y), .B(D8577_Y),     .C(D6407_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8529 ( .Y(D8529_Y), .D(D8378_Y), .B(D8578_Y),     .C(D10191_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8527 ( .Y(D8527_Y), .D(D8378_Y), .B(D8528_Y),     .C(D462_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8526 ( .Y(D8526_Y), .D(D8370_Y), .B(D8490_Y),     .C(D1813_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8525 ( .Y(D8525_Y), .D(D8370_Y), .B(D8489_Y),     .C(D6410_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8524 ( .Y(D8524_Y), .D(D8378_Y), .B(D8491_Y),     .C(D463_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8523 ( .Y(D8523_Y), .D(D8370_Y), .B(D8483_Y),     .C(D6406_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8522 ( .Y(D8522_Y), .D(D8378_Y), .B(D8486_Y),     .C(D1964_Y), .A(D8533_Y));
KC_OAI22BB_X1 D8454 ( .Y(D8454_Y), .D(D10192_Y), .B(D8367_Y),     .C(D1836_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8452 ( .Y(D8452_Y), .D(D8280_Y), .B(D8414_Y),     .C(D6407_Y), .A(D8227_Y));
KC_OAI22BB_X1 D8451 ( .Y(D8451_Y), .D(D8280_Y), .B(D8306_Y),     .C(D10191_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8450 ( .Y(D8450_Y), .D(D8280_Y), .B(D8448_Y),     .C(D1964_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8449 ( .Y(D8449_Y), .D(D8386_Y), .B(D8400_Y),     .C(D8383_Y), .A(D8387_Y));
KC_OAI22BB_X1 D8447 ( .Y(D8447_Y), .D(D8464_Y), .B(D8387_Y),     .C(D6405_Y), .A(D8455_Y));
KC_OAI22BB_X1 D8446 ( .Y(D8446_Y), .D(D10191_Y), .B(D8372_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D8445 ( .Y(D8445_Y), .D(D1846_Y), .B(D8376_Y),     .C(D9617_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8444 ( .Y(D8444_Y), .D(D8464_Y), .B(D8388_Y),     .C(D1964_Y), .A(D8455_Y));
KC_OAI22BB_X1 D8443 ( .Y(D8443_Y), .D(D8464_Y), .B(D8394_Y),     .C(D464_Y), .A(D8455_Y));
KC_OAI22BB_X1 D8442 ( .Y(D8442_Y), .D(D9617_Y), .B(D8440_Y),     .C(D1836_Y), .A(D8455_Y));
KC_OAI22BB_X1 D8316 ( .Y(D8316_Y), .D(D6772_Y), .B(D6693_Y),     .C(D8355_Y), .A(D6759_Y));
KC_OAI22BB_X1 D8315 ( .Y(D8315_Y), .D(D8356_Y), .B(D16197_Y),     .C(D8321_Y), .A(D16096_Y));
KC_OAI22BB_X1 D8314 ( .Y(D8314_Y), .D(D6772_Y), .B(D6698_Y),     .C(D8325_Y), .A(D6759_Y));
KC_OAI22BB_X1 D8311 ( .Y(D8311_Y), .D(D8280_Y), .B(D2210_Y),     .C(D464_Y), .A(D8431_Y));
KC_OAI22BB_X1 D8308 ( .Y(D8308_Y), .D(D8280_Y), .B(D8304_Y),     .C(D462_Y), .A(D8227_Y));
KC_OAI22BB_X1 D8307 ( .Y(D8307_Y), .D(D8280_Y), .B(D880_Y), .C(D463_Y),     .A(D8227_Y));
KC_OAI22BB_X1 D8303 ( .Y(D8303_Y), .D(D8280_Y), .B(D8305_Y),     .C(D10192_Y), .A(D8227_Y));
KC_OAI22BB_X1 D8134 ( .Y(D8134_Y), .D(D6490_Y), .B(D8141_Y),     .C(D1964_Y), .A(D8212_Y));
KC_OAI22BB_X1 D8132 ( .Y(D8132_Y), .D(D8259_Y), .B(D5213_Y),     .C(D6772_Y), .A(D6759_Y));
KC_OAI22BB_X1 D8131 ( .Y(D8131_Y), .D(D8130_Y), .B(D8246_Q),     .C(D8076_Y), .A(D8147_Q));
KC_OAI22BB_X1 D8046 ( .Y(D8046_Y), .D(D6490_Y), .B(D8036_Y),     .C(D10191_Y), .A(D8212_Y));
KC_OAI22BB_X1 D8042 ( .Y(D8042_Y), .D(D6490_Y), .B(D8041_Y),     .C(D6407_Y), .A(D8212_Y));
KC_OAI22BB_X1 D8039 ( .Y(D8039_Y), .D(D6490_Y), .B(D8040_Y),     .C(D10192_Y), .A(D8212_Y));
KC_OAI22BB_X1 D8035 ( .Y(D8035_Y), .D(D6490_Y), .B(D8037_Y),     .C(D6405_Y), .A(D8212_Y));
KC_OAI22BB_X1 D8032 ( .Y(D8032_Y), .D(D6490_Y), .B(D8043_Y),     .C(D462_Y), .A(D8212_Y));
KC_OAI22BB_X1 D7956 ( .Y(D7956_Y), .D(D7910_Y), .B(D6544_Q),     .C(D6517_Y), .A(D7911_Y));
KC_OAI22BB_X1 D7778 ( .Y(D7778_Y), .D(D4770_Y), .B(D8062_Y),     .C(D9354_Y), .A(D7771_Y));
KC_OAI22BB_X1 D7517 ( .Y(D7517_Y), .D(D9269_Y), .B(D7608_Y),     .C(D1709_Y), .A(D266_Y));
KC_OAI22BB_X1 D7386 ( .Y(D7386_Y), .D(D5864_Y), .B(D7358_Y),     .C(D5656_Y), .A(D7153_Y));
KC_OAI22BB_X1 D7384 ( .Y(D7384_Y), .D(D5710_Y), .B(D7984_Y),     .C(D5846_Y), .A(D5684_Y));
KC_OAI22BB_X1 D7287 ( .Y(D7287_Y), .D(D7211_Y), .B(D7408_Y),     .C(D7119_Y), .A(D5671_Y));
KC_OAI22BB_X1 D7285 ( .Y(D7285_Y), .D(D8877_Y), .B(D5783_Y),     .C(D7204_Y), .A(D7_Y));
KC_OAI22BB_X1 D6955 ( .Y(D6955_Y), .D(D8378_Y), .B(D6926_Y),     .C(D6410_Y), .A(D8431_Y));
KC_OAI22BB_X1 D6950 ( .Y(D6950_Y), .D(D8378_Y), .B(D6948_Y),     .C(D1813_Y), .A(D8431_Y));
KC_OAI22BB_X1 D6949 ( .Y(D6949_Y), .D(D8378_Y), .B(D6920_Y),     .C(D1814_Y), .A(D8431_Y));
KC_OAI22BB_X1 D6947 ( .Y(D6947_Y), .D(D8378_Y), .B(D1755_Y),     .C(D6406_Y), .A(D8431_Y));
KC_OAI22BB_X1 D6886 ( .Y(D6886_Y), .D(D8378_Y), .B(D64_Y), .C(D9617_Y),     .A(D8431_Y));
KC_OAI22BB_X1 D6885 ( .Y(D6885_Y), .D(D8378_Y), .B(D6937_Y),     .C(D8336_Y), .A(D8431_Y));
KC_OAI22BB_X1 D6807 ( .Y(D6807_Y), .D(D8280_Y), .B(D6804_Y),     .C(D8336_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6806 ( .Y(D6806_Y), .D(D8280_Y), .B(D6789_Y),     .C(D10358_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6803 ( .Y(D6803_Y), .D(D6490_Y), .B(D1758_Y),     .C(D8336_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6802 ( .Y(D6802_Y), .D(D6490_Y), .B(D6785_Y),     .C(D10358_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6799 ( .Y(D6799_Y), .D(D8280_Y), .B(D6801_Y),     .C(D6406_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6796 ( .Y(D6796_Y), .D(D1846_Y), .B(D881_Y),     .C(D8336_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6739 ( .Y(D6739_Y), .D(D8280_Y), .B(D6737_Y),     .C(D6410_Y), .A(D8212_Y));
KC_OAI22BB_X1 D6738 ( .Y(D6738_Y), .D(D8280_Y), .B(D6741_Y),     .C(D1814_Y), .A(D8212_Y));
KC_OAI22BB_X1 D6736 ( .Y(D6736_Y), .D(D8280_Y), .B(D6734_Y),     .C(D1813_Y), .A(D8212_Y));
KC_OAI22BB_X1 D6732 ( .Y(D6732_Y), .D(D6490_Y), .B(D6740_Y),     .C(D813_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6729 ( .Y(D6729_Y), .D(D8280_Y), .B(D6733_Y),     .C(D813_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6728 ( .Y(D6728_Y), .D(D8280_Y), .B(D6730_Y),     .C(D9617_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6727 ( .Y(D6727_Y), .D(D6490_Y), .B(D1690_Y),     .C(D9617_Y), .A(D8227_Y));
KC_OAI22BB_X1 D6650 ( .Y(D6650_Y), .D(D6490_Y), .B(D6651_Y),     .C(D463_Y), .A(D8212_Y));
KC_OAI22BB_X1 D6648 ( .Y(D6648_Y), .D(D6490_Y), .B(D6644_Y),     .C(D1814_Y), .A(D8212_Y));
KC_OAI22BB_X1 D6642 ( .Y(D6642_Y), .D(D6490_Y), .B(D6643_Y),     .C(D6410_Y), .A(D8212_Y));
KC_OAI22BB_X1 D6593 ( .Y(D6593_Y), .D(D6490_Y), .B(D8033_Y),     .C(D1813_Y), .A(D8212_Y));
KC_OAI22BB_X1 D6536 ( .Y(D6536_Y), .D(D6508_Y), .B(D6551_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6535 ( .Y(D6535_Y), .D(D6507_Y), .B(D524_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6533 ( .Y(D6533_Y), .D(D7908_Y), .B(D515_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6532 ( .Y(D6532_Y), .D(D6498_Y), .B(D6550_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6531 ( .Y(D6531_Y), .D(D6499_Y), .B(D519_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6530 ( .Y(D6530_Y), .D(D6504_Y), .B(D6548_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6529 ( .Y(D6529_Y), .D(D6509_Y), .B(D6549_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6528 ( .Y(D6528_Y), .D(D6501_Y), .B(D6546_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6527 ( .Y(D6527_Y), .D(D1692_Y), .B(D6539_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D6526 ( .Y(D6526_Y), .D(D7909_Y), .B(D6540_Q),     .C(D6517_Y), .A(D7911_Y));
KC_OAI22BB_X1 D6523 ( .Y(D6523_Y), .D(D6502_Y), .B(D513_Q),     .C(D6517_Y), .A(D7920_Y));
KC_OAI22BB_X1 D5929 ( .Y(D5929_Y), .D(D6024_Y), .B(D5871_Y),     .C(D5868_Y), .A(D249_Y));
KC_OAI22BB_X1 D5924 ( .Y(D5924_Y), .D(D5888_Y), .B(D7461_Y),     .C(D5857_Y), .A(D247_Y));
KC_OAI22BB_X1 D5796 ( .Y(D5796_Y), .D(D7292_Y), .B(D4378_Y),     .C(D7211_Y), .A(D5698_Y));
KC_OAI22BB_X1 D5074 ( .Y(D5074_Y), .D(D5042_Y), .B(D1415_Y),     .C(D4865_Y), .A(D4877_Y));
KC_OAI22BB_X1 D5072 ( .Y(D5072_Y), .D(D4880_Y), .B(D5029_Y),     .C(D5023_Y), .A(D4897_Y));
KC_OAI22BB_X1 D4710 ( .Y(D4710_Y), .D(D4763_Y), .B(D4798_Y),     .C(D3203_Y), .A(D4660_Y));
KC_OAI22BB_X1 D4079 ( .Y(D4079_Y), .D(D4035_Y), .B(D4035_Y),     .C(D4076_Y), .A(D4038_Y));
KC_OAI22BB_X1 D3557 ( .Y(D3557_Y), .D(D3511_Y), .B(D3514_Y),     .C(D3576_Q), .A(D4887_Y));
KC_OAI22BB_X1 D3555 ( .Y(D3555_Y), .D(D3603_Y), .B(D3633_Y),     .C(D5083_Y), .A(D3603_Y));
KC_OAI22BB_X1 D3474 ( .Y(D3474_Y), .D(D3520_Y), .B(D3414_Y),     .C(D3431_Y), .A(D4911_Y));
KC_OAI22BB_X1 D2875 ( .Y(D2875_Y), .D(D2895_Y), .B(D2802_Y),     .C(D2743_Y), .A(D2743_Y));
KC_OAI22BB_X1 D2872 ( .Y(D2872_Y), .D(D2_Y), .B(D2837_Y), .C(D2804_Y),     .A(D2885_Q));
KC_OAI22BB_X1 D2785 ( .Y(D2785_Y), .D(D2767_Y), .B(D2875_Y),     .C(D2809_Y), .A(D2781_Y));
KC_OAI22BB_X1 D2335 ( .Y(D2335_Y), .D(D12770_Y), .B(D12417_Q),     .C(D2328_Y), .A(D2326_Y));
KC_OAI22BB_X1 D2334 ( .Y(D2334_Y), .D(D12771_Y), .B(D12342_Q),     .C(D2328_Y), .A(D2326_Y));
KC_OAI22BB_X1 D2333 ( .Y(D2333_Y), .D(D12771_Y), .B(D12416_Q),     .C(D2327_Y), .A(D2325_Y));
KC_OAI22BB_X1 D2332 ( .Y(D2332_Y), .D(D12309_Y), .B(D12794_Y),     .C(D12855_Q), .A(D2393_Q));
KC_OAI22BB_X1 D2281 ( .Y(D2281_Y), .D(D8470_Y), .B(D2282_Y),     .C(D10358_Y), .A(D10788_Y));
KC_OAI22BB_X1 D2280 ( .Y(D2280_Y), .D(D8470_Y), .B(D2241_Y),     .C(D9617_Y), .A(D10788_Y));
KC_OAI22BB_X1 D2279 ( .Y(D2279_Y), .D(D8461_Y), .B(D12033_Y),     .C(D10191_Y), .A(D8430_Y));
KC_OAI22BB_X1 D2278 ( .Y(D2278_Y), .D(D8461_Y), .B(D11464_Y),     .C(D10358_Y), .A(D8430_Y));
KC_OAI22BB_X1 D2239 ( .Y(D2239_Y), .D(D8470_Y), .B(D2240_Y),     .C(D464_Y), .A(D10788_Y));
KC_OAI22BB_X1 D2236 ( .Y(D2236_Y), .D(D8461_Y), .B(D11529_Y),     .C(D6407_Y), .A(D8431_Y));
KC_OAI22BB_X1 D2065 ( .Y(D2065_Y), .D(D1907_Y), .B(D8068_Y),     .C(D2027_Y), .A(D7473_Y));
KC_OAI22BB_X1 D2064 ( .Y(D2064_Y), .D(D1907_Y), .B(D9333_Y),     .C(D8877_Y), .A(D9068_Y));
KC_OAI22BB_X1 D1916 ( .Y(D1916_Y), .D(D6490_Y), .B(D1843_Y),     .C(D6406_Y), .A(D8212_Y));
KC_OAI22BB_X1 D1913 ( .Y(D1913_Y), .D(D8378_Y), .B(D8576_Y),     .C(D6405_Y), .A(D8533_Y));
KC_OAI22BB_X1 D1912 ( .Y(D1912_Y), .D(D8378_Y), .B(D8480_Y),     .C(D10192_Y), .A(D8533_Y));
KC_OAI22BB_X1 D1911 ( .Y(D1911_Y), .D(D8370_Y), .B(D8479_Y),     .C(D10192_Y), .A(D8533_Y));
KC_OAI22BB_X1 D1767 ( .Y(D1767_Y), .D(D1769_Y), .B(D6198_Y),     .C(D6637_Y), .A(D6173_Y));
KC_OAI22BB_X1 D1762 ( .Y(D1762_Y), .D(D4747_Y), .B(D1785_Q),     .C(D8018_Y), .A(D8212_Y));
KC_OAI22BB_X1 D1757 ( .Y(D1757_Y), .D(D8378_Y), .B(D6953_Y),     .C(D10358_Y), .A(D8431_Y));
KC_OAI22BB_X1 D1756 ( .Y(D1756_Y), .D(D8378_Y), .B(D6951_Y),     .C(D813_Y), .A(D8431_Y));
KC_OAI22BB_X1 D1466 ( .Y(D1466_Y), .D(D3447_Y), .B(D3489_Y),     .C(D4748_Y), .A(D1570_Y));
KC_OAI22BB_X1 D1114 ( .Y(D1114_Y), .D(D8461_Y), .B(D11533_Y),     .C(D462_Y), .A(D8430_Y));
KC_OAI22BB_X1 D1112 ( .Y(D1112_Y), .D(D8461_Y), .B(D11461_Y),     .C(D6410_Y), .A(D8430_Y));
KC_OAI22BB_X1 D1110 ( .Y(D1110_Y), .D(D813_Y), .B(D1979_Y),     .C(D8370_Y), .A(D8533_Y));
KC_OAI22BB_X1 D1109 ( .Y(D1109_Y), .D(D8370_Y), .B(D1084_Y),     .C(D463_Y), .A(D8533_Y));
KC_OAI22BB_X1 D1001 ( .Y(D1001_Y), .D(D1846_Y), .B(D8439_Y),     .C(D10358_Y), .A(D8431_Y));
KC_OAI22BB_X1 D889 ( .Y(D889_Y), .D(D8464_Y), .B(D11313_Y),     .C(D1813_Y), .A(D10788_Y));
KC_OAI22BB_X1 D887 ( .Y(D887_Y), .D(D8464_Y), .B(D11314_Y),     .C(D9617_Y), .A(D10788_Y));
KC_OAI22BB_X1 D882 ( .Y(D882_Y), .D(D8280_Y), .B(D2209_Y), .C(D6405_Y),     .A(D8431_Y));
KC_OAI22BB_X1 D773 ( .Y(D773_Y), .D(D8470_Y), .B(D11242_Y),     .C(D1814_Y), .A(D10788_Y));
KC_OAI22BB_X1 D771 ( .Y(D771_Y), .D(D15531_Y), .B(D15803_Y),     .C(D16800_Y), .A(D15563_Y));
KC_OAI22BB_X1 D650 ( .Y(D650_Y), .D(D16140_Y), .B(D16140_Y),     .C(D16107_Y), .A(D15441_Y));
KC_OAI22BB_X1 D578 ( .Y(D578_Y), .D(D6490_Y), .B(D8005_Y), .C(D464_Y),     .A(D8212_Y));
KC_OAI22BB_X1 D498 ( .Y(D498_Y), .D(D6503_Y), .B(D5131_Q), .C(D6517_Y),     .A(D7920_Y));
KC_OAI22BB_X1 D497 ( .Y(D497_Y), .D(D392_Y), .B(D5142_Q), .C(D8018_Y),     .A(D8212_Y));
KC_OAI22BB_X1 D348 ( .Y(D348_Y), .D(D1865_Y), .B(D5966_Y), .C(D8908_Y),     .A(D8709_Q));
KC_OAI22BB_X1 D318 ( .Y(D318_Y), .D(D10142_Y), .B(D6271_Y),     .C(D1709_Y), .A(D266_Y));
KC_OAI22BB_X1 D103 ( .Y(D103_Y), .D(D15453_Y), .B(D15395_Y),     .C(D15453_Y), .A(D2630_Y));
KC_AOI22_X4 D172 ( .A1(D9482_Y), .B0(D8748_Y), .B1(D2054_Y),     .Y(D172_Y), .A0(D1975_Y));
KC_NAND2_X3 D7163 ( .Y(D7163_Y), .B(D5804_Y), .A(D7153_Y));
KC_NAND2_X3 D171 ( .Y(D171_Y), .B(D11536_Y), .A(D2229_Y));
KC_OAI21_X3 D13636 ( .A1(D13409_Y), .B(D13504_Y), .A0(D2443_Y),     .Y(D13636_Y));
KC_OAI21_X3 D13635 ( .A1(D13409_Y), .B(D13595_Y), .A0(D13508_Y),     .Y(D13635_Y));
KC_OAI21_X3 D13634 ( .A1(D13409_Y), .B(D13586_Y), .A0(D13585_Y),     .Y(D13634_Y));
KC_OAI21_X3 D13526 ( .A1(D13409_Y), .B(D13502_Y), .A0(D13488_Y),     .Y(D13526_Y));
KC_OAI21_X3 D13525 ( .A1(D13409_Y), .B(D13505_Y), .A0(D13484_Y),     .Y(D13525_Y));
KC_OAI21_X3 D13524 ( .A1(D13409_Y), .B(D13507_Y), .A0(D13493_Y),     .Y(D13524_Y));
KC_OAI21_X3 D7405 ( .A1(D7358_Y), .B(D7377_Y), .A0(D7163_Y),     .Y(D7405_Y));
KC_OAI21_X3 D6408 ( .A1(D6483_Y), .B(D6291_Y), .A0(D6447_Y),     .Y(D6408_Y));
KC_OAI21_X3 D1823 ( .A1(D6281_Y), .B(D1822_Y), .A0(D8018_Y),     .Y(D1823_Y));
KC_OAI21_X3 D1072 ( .A1(D13409_Y), .B(D13580_Y), .A0(D13584_Y),     .Y(D1072_Y));
KC_OAI21_X3 D169 ( .A1(D6287_Y), .B(D1674_Y), .A0(D8018_Y),     .Y(D169_Y));
KC_INV_X1 D16695 ( .Y(D16695_Y), .A(D16694_Y));
KC_INV_X1 D16693 ( .Y(D16693_Y), .A(D16692_Y));
KC_INV_X1 D16691 ( .Y(D16691_Y), .A(D16690_Y));
KC_INV_X1 D16689 ( .Y(D16689_Y), .A(D16688_Y));
KC_INV_X1 D16671 ( .Y(D16671_Y), .A(D16670_Y));
KC_INV_X1 D16669 ( .Y(D16669_Y), .A(D16668_Y));
KC_INV_X1 D16665 ( .Y(D16665_Y), .A(D16666_Y));
KC_INV_X1 D16655 ( .Y(D16655_Y), .A(D16660_Q));
KC_INV_X1 D16646 ( .Y(D16646_Y), .A(D1406_Y));
KC_INV_X1 D16643 ( .Y(D16643_Y), .A(D16642_Y));
KC_INV_X1 D16640 ( .Y(D16640_Y), .A(D2691_Y));
KC_INV_X1 D16595 ( .Y(D16595_Y), .A(D16598_Q));
KC_INV_X1 D16561 ( .Y(D16561_Y), .A(D16564_Q));
KC_INV_X1 D16543 ( .Y(D16543_Y), .A(D16558_Q));
KC_INV_X1 D16541 ( .Y(D16541_Y), .A(D16547_Y));
KC_INV_X1 D16537 ( .Y(D16537_Y), .A(D1385_Q));
KC_INV_X1 D16536 ( .Y(D16536_Y), .A(D16556_Q));
KC_INV_X1 D16533 ( .Y(D16533_Y), .A(D16387_Q));
KC_INV_X1 D16501 ( .Y(D16501_Y), .A(D16497_Y));
KC_INV_X1 D16494 ( .Y(D16494_Y), .A(D1343_Y));
KC_INV_X1 D16492 ( .Y(D16492_Y), .A(D16530_Y));
KC_INV_X1 D16488 ( .Y(D16488_Y), .A(D1381_Q));
KC_INV_X1 D16482 ( .Y(D16482_Y), .A(D16405_Y));
KC_INV_X1 D16481 ( .Y(D16481_Y), .A(D16472_Q));
KC_INV_X1 D16466 ( .Y(D16466_Y), .A(D16478_Y));
KC_INV_X1 D16463 ( .Y(D16463_Y), .A(D16416_Y));
KC_INV_X1 D16444 ( .Y(D16444_Y), .A(D1324_Q));
KC_INV_X1 D16443 ( .Y(D16443_Y), .A(D16459_Q));
KC_INV_X1 D16439 ( .Y(D16439_Y), .A(D1378_Q));
KC_INV_X1 D16438 ( .Y(D16438_Y), .A(D16470_Q));
KC_INV_X1 D16433 ( .Y(D16433_Y), .A(D16471_Q));
KC_INV_X1 D16430 ( .Y(D16430_Y), .A(D16461_Y));
KC_INV_X1 D16429 ( .Y(D16429_Y), .A(D1281_Y));
KC_INV_X1 D16426 ( .Y(D16426_Y), .A(D1322_Q));
KC_INV_X1 D16425 ( .Y(D16425_Y), .A(D16473_Q));
KC_INV_X1 D16422 ( .Y(D16422_Y), .A(D16449_Y));
KC_INV_X1 D16419 ( .Y(D16419_Y), .A(D16424_Y));
KC_INV_X1 D16373 ( .Y(D16373_Y), .A(D16400_Y));
KC_INV_X1 D16347 ( .Y(D16347_Y), .A(D16360_Q));
KC_INV_X1 D16305 ( .Y(D16305_Y), .A(D16362_Q));
KC_INV_X1 D16266 ( .Y(D16266_Y), .A(D16289_Q));
KC_INV_X1 D16265 ( .Y(D16265_Y), .A(D2681_Q));
KC_INV_X1 D16261 ( .Y(D16261_Y), .A(D16291_Q));
KC_INV_X1 D16257 ( .Y(D16257_Y), .A(D2680_Q));
KC_INV_X1 D16256 ( .Y(D16256_Y), .A(D16292_Q));
KC_INV_X1 D16255 ( .Y(D16255_Y), .A(D16260_Y));
KC_INV_X1 D16254 ( .Y(D16254_Y), .A(D16246_Y));
KC_INV_X1 D16192 ( .Y(D16192_Y), .A(D16270_Y));
KC_INV_X1 D16188 ( .Y(D16188_Y), .A(D16187_Y));
KC_INV_X1 D16120 ( .Y(D16120_Y), .A(D16103_Y));
KC_INV_X1 D16119 ( .Y(D16119_Y), .A(D16137_Y));
KC_INV_X1 D16118 ( .Y(D16118_Y), .A(D16127_Y));
KC_INV_X1 D16115 ( .Y(D16115_Y), .A(D16161_Y));
KC_INV_X1 D16114 ( .Y(D16114_Y), .A(D2651_Y));
KC_INV_X1 D16111 ( .Y(D16111_Y), .A(D16108_Y));
KC_INV_X1 D16110 ( .Y(D16110_Y), .A(D16155_Y));
KC_INV_X1 D16107 ( .Y(D16107_Y), .A(D2591_Y));
KC_INV_X1 D16106 ( .Y(D16106_Y), .A(D15329_Y));
KC_INV_X1 D16105 ( .Y(D16105_Y), .A(D16182_Y));
KC_INV_X1 D16104 ( .Y(D16104_Y), .A(D16180_Y));
KC_INV_X1 D16103 ( .Y(D16103_Y), .A(D16148_Y));
KC_INV_X1 D16102 ( .Y(D16102_Y), .A(D16150_Y));
KC_INV_X1 D16101 ( .Y(D16101_Y), .A(D16100_Y));
KC_INV_X1 D16061 ( .Y(D16061_Y), .A(D16033_Y));
KC_INV_X1 D16060 ( .Y(D16060_Y), .A(D15306_Y));
KC_INV_X1 D16059 ( .Y(D16059_Y), .A(D16043_Y));
KC_INV_X1 D16054 ( .Y(D16054_Y), .A(D15335_Y));
KC_INV_X1 D16053 ( .Y(D16053_Y), .A(D16088_Y));
KC_INV_X1 D16049 ( .Y(D16049_Y), .A(D16084_Y));
KC_INV_X1 D15971 ( .Y(D15971_Y), .A(D1326_Q));
KC_INV_X1 D15969 ( .Y(D15969_Y), .A(D1273_Y));
KC_INV_X1 D15964 ( .Y(D15964_Y), .A(D15991_Q));
KC_INV_X1 D15961 ( .Y(D15961_Y), .A(D16013_Q));
KC_INV_X1 D15960 ( .Y(D15960_Y), .A(D15992_Q));
KC_INV_X1 D15958 ( .Y(D15958_Y), .A(D14698_Y));
KC_INV_X1 D15913 ( .Y(D15913_Y), .A(D142_Q));
KC_INV_X1 D15910 ( .Y(D15910_Y), .A(D16392_Q));
KC_INV_X1 D15909 ( .Y(D15909_Y), .A(D2638_Q));
KC_INV_X1 D15899 ( .Y(D15899_Y), .A(D15949_Q));
KC_INV_X1 D15897 ( .Y(D15897_Y), .A(D15995_Q));
KC_INV_X1 D15896 ( .Y(D15896_Y), .A(D1230_Q));
KC_INV_X1 D15895 ( .Y(D15895_Y), .A(D1233_Q));
KC_INV_X1 D15888 ( .Y(D15888_Y), .A(D1228_Q));
KC_INV_X1 D15884 ( .Y(D15884_Y), .A(D1229_Q));
KC_INV_X1 D15883 ( .Y(D15883_Y), .A(D1236_Q));
KC_INV_X1 D15882 ( .Y(D15882_Y), .A(D15998_Q));
KC_INV_X1 D15831 ( .Y(D15831_Y), .A(D16358_Q));
KC_INV_X1 D15829 ( .Y(D15829_Y), .A(D16369_Q));
KC_INV_X1 D15826 ( .Y(D15826_Y), .A(D144_Q));
KC_INV_X1 D15823 ( .Y(D15823_Y), .A(D16354_Q));
KC_INV_X1 D15821 ( .Y(D15821_Y), .A(D1156_Q));
KC_INV_X1 D15820 ( .Y(D15820_Y), .A(D16355_Q));
KC_INV_X1 D15818 ( .Y(D15818_Y), .A(D15872_Q));
KC_INV_X1 D15810 ( .Y(D15810_Y), .A(D1149_Q));
KC_INV_X1 D15745 ( .Y(D15745_Y), .A(D1050_Q));
KC_INV_X1 D15739 ( .Y(D15739_Y), .A(D16319_Q));
KC_INV_X1 D15735 ( .Y(D15735_Y), .A(D2640_Q));
KC_INV_X1 D15734 ( .Y(D15734_Y), .A(D15796_Q));
KC_INV_X1 D15729 ( .Y(D15729_Y), .A(D16318_Q));
KC_INV_X1 D15728 ( .Y(D15728_Y), .A(D16340_Q));
KC_INV_X1 D15720 ( .Y(D15720_Y), .A(D16316_Q));
KC_INV_X1 D15715 ( .Y(D15715_Y), .A(D15873_Q));
KC_INV_X1 D15707 ( .Y(D15707_Y), .A(D14845_Y));
KC_INV_X1 D15706 ( .Y(D15706_Y), .A(D15621_Y));
KC_INV_X1 D15704 ( .Y(D15704_Y), .A(D15615_Y));
KC_INV_X1 D15703 ( .Y(D15703_Y), .A(D15633_Y));
KC_INV_X1 D15647 ( .Y(D15647_Y), .A(D15632_Y));
KC_INV_X1 D15630 ( .Y(D15630_Y), .A(D16293_Q));
KC_INV_X1 D15629 ( .Y(D15629_Y), .A(D15651_Y));
KC_INV_X1 D15628 ( .Y(D15628_Y), .A(D2607_Y));
KC_INV_X1 D15617 ( .Y(D15617_Y), .A(D15634_Y));
KC_INV_X1 D15611 ( .Y(D15611_Y), .A(D16461_Y));
KC_INV_X1 D15610 ( .Y(D15610_Y), .A(D2611_Y));
KC_INV_X1 D15607 ( .Y(D15607_Y), .A(D14564_Y));
KC_INV_X1 D15606 ( .Y(D15606_Y), .A(D15518_Y));
KC_INV_X1 D15605 ( .Y(D15605_Y), .A(D15513_Y));
KC_INV_X1 D15603 ( .Y(D15603_Y), .A(D15527_Y));
KC_INV_X1 D15602 ( .Y(D15602_Y), .A(D15519_Y));
KC_INV_X1 D15531 ( .Y(D15531_Y), .A(D15522_Y));
KC_INV_X1 D15526 ( .Y(D15526_Y), .A(D15385_Y));
KC_INV_X1 D15516 ( .Y(D15516_Y), .A(D755_Y));
KC_INV_X1 D15509 ( .Y(D15509_Y), .A(D3707_Y));
KC_INV_X1 D15508 ( .Y(D15508_Y), .A(D16275_Y));
KC_INV_X1 D15503 ( .Y(D15503_Y), .A(D15502_Y));
KC_INV_X1 D15497 ( .Y(D15497_Y), .A(D15341_Y));
KC_INV_X1 D15489 ( .Y(D15489_Y), .A(D15626_Y));
KC_INV_X1 D15488 ( .Y(D15488_Y), .A(D15657_Y));
KC_INV_X1 D15485 ( .Y(D15485_Y), .A(D15482_Y));
KC_INV_X1 D15484 ( .Y(D15484_Y), .A(D14719_Y));
KC_INV_X1 D15476 ( .Y(D15476_Y), .A(D816_Q));
KC_INV_X1 D15473 ( .Y(D15473_Y), .A(D2604_Y));
KC_INV_X1 D15472 ( .Y(D15472_Y), .A(D15465_Y));
KC_INV_X1 D15471 ( .Y(D15471_Y), .A(D15480_Y));
KC_INV_X1 D15409 ( .Y(D15409_Y), .A(D15270_Y));
KC_INV_X1 D15408 ( .Y(D15408_Y), .A(D564_Y));
KC_INV_X1 D15407 ( .Y(D15407_Y), .A(D16056_Y));
KC_INV_X1 D15404 ( .Y(D15404_Y), .A(D14749_Y));
KC_INV_X1 D15397 ( .Y(D15397_Y), .A(D15271_Y));
KC_INV_X1 D15395 ( .Y(D15395_Y), .A(D13186_Y));
KC_INV_X1 D15390 ( .Y(D15390_Y), .A(D16037_Y));
KC_INV_X1 D15380 ( .Y(D15380_Y), .A(D650_Y));
KC_INV_X1 D15378 ( .Y(D15378_Y), .A(D15373_Y));
KC_INV_X1 D15377 ( .Y(D15377_Y), .A(D14513_Y));
KC_INV_X1 D15367 ( .Y(D15367_Y), .A(D15363_Y));
KC_INV_X1 D15366 ( .Y(D15366_Y), .A(D15359_Y));
KC_INV_X1 D15365 ( .Y(D15365_Y), .A(D15374_Y));
KC_INV_X1 D15357 ( .Y(D15357_Y), .A(D15523_Y));
KC_INV_X1 D15355 ( .Y(D15355_Y), .A(D15521_Y));
KC_INV_X1 D15354 ( .Y(D15354_Y), .A(D636_Y));
KC_INV_X1 D15353 ( .Y(D15353_Y), .A(D15530_Y));
KC_INV_X1 D15352 ( .Y(D15352_Y), .A(D14625_Y));
KC_INV_X1 D15346 ( .Y(D15346_Y), .A(D15551_Y));
KC_INV_X1 D15345 ( .Y(D15345_Y), .A(D15375_Y));
KC_INV_X1 D15344 ( .Y(D15344_Y), .A(D15349_Y));
KC_INV_X1 D15302 ( .Y(D15302_Y), .A(D15305_Y));
KC_INV_X1 D15300 ( .Y(D15300_Y), .A(D15304_Y));
KC_INV_X1 D15291 ( .Y(D15291_Y), .A(D2636_Y));
KC_INV_X1 D15290 ( .Y(D15290_Y), .A(D16090_Y));
KC_INV_X1 D15280 ( .Y(D15280_Y), .A(D16089_Y));
KC_INV_X1 D15244 ( .Y(D15244_Y), .A(D327_Y));
KC_INV_X1 D15243 ( .Y(D15243_Y), .A(D15250_Y));
KC_INV_X1 D15241 ( .Y(D15241_Y), .A(D15240_Y));
KC_INV_X1 D15226 ( .Y(D15226_Y), .A(D15238_Q));
KC_INV_X1 D15224 ( .Y(D15224_Y), .A(D1377_Q));
KC_INV_X1 D15172 ( .Y(D15172_Y), .A(D15237_Q));
KC_INV_X1 D15165 ( .Y(D15165_Y), .A(D1384_Q));
KC_INV_X1 D15164 ( .Y(D15164_Y), .A(D16009_Q));
KC_INV_X1 D15161 ( .Y(D15161_Y), .A(D15229_Q));
KC_INV_X1 D15110 ( .Y(D15110_Y), .A(D1327_Q));
KC_INV_X1 D15107 ( .Y(D15107_Y), .A(D15236_Q));
KC_INV_X1 D15106 ( .Y(D15106_Y), .A(D15231_Q));
KC_INV_X1 D15102 ( .Y(D15102_Y), .A(D1153_Q));
KC_INV_X1 D15101 ( .Y(D15101_Y), .A(D15134_Q));
KC_INV_X1 D15099 ( .Y(D15099_Y), .A(D1231_Q));
KC_INV_X1 D15094 ( .Y(D15094_Y), .A(D16385_Q));
KC_INV_X1 D15048 ( .Y(D15048_Y), .A(D14300_Q));
KC_INV_X1 D15039 ( .Y(D15039_Y), .A(D15874_Q));
KC_INV_X1 D15032 ( .Y(D15032_Y), .A(D1154_Q));
KC_INV_X1 D15025 ( .Y(D15025_Y), .A(D15871_Q));
KC_INV_X1 D15019 ( .Y(D15019_Y), .A(D16356_Q));
KC_INV_X1 D15018 ( .Y(D15018_Y), .A(D1151_Q));
KC_INV_X1 D15009 ( .Y(D15009_Y), .A(D15669_Q));
KC_INV_X1 D15008 ( .Y(D15008_Y), .A(D16393_Q));
KC_INV_X1 D14947 ( .Y(D14947_Y), .A(D1052_Q));
KC_INV_X1 D14946 ( .Y(D14946_Y), .A(D2641_Q));
KC_INV_X1 D14941 ( .Y(D14941_Y), .A(D924_Q));
KC_INV_X1 D14935 ( .Y(D14935_Y), .A(D14872_Q));
KC_INV_X1 D14934 ( .Y(D14934_Y), .A(D16314_Q));
KC_INV_X1 D14933 ( .Y(D14933_Y), .A(D15794_Q));
KC_INV_X1 D14928 ( .Y(D14928_Y), .A(D14995_Q));
KC_INV_X1 D14924 ( .Y(D14924_Y), .A(D16317_Q));
KC_INV_X1 D14922 ( .Y(D14922_Y), .A(D14263_Q));
KC_INV_X1 D14916 ( .Y(D14916_Y), .A(D1048_Q));
KC_INV_X1 D14915 ( .Y(D14915_Y), .A(D143_Q));
KC_INV_X1 D14912 ( .Y(D14912_Y), .A(D14876_Q));
KC_INV_X1 D14911 ( .Y(D14911_Y), .A(D14815_Q));
KC_INV_X1 D14854 ( .Y(D14854_Y), .A(D14813_Y));
KC_INV_X1 D14847 ( .Y(D14847_Y), .A(D14841_Y));
KC_INV_X1 D14830 ( .Y(D14830_Y), .A(D14563_Y));
KC_INV_X1 D14828 ( .Y(D14828_Y), .A(D14081_Y));
KC_INV_X1 D14821 ( .Y(D14821_Y), .A(D15674_Y));
KC_INV_X1 D14809 ( .Y(D14809_Y), .A(D14788_Q));
KC_INV_X1 D14748 ( .Y(D14748_Y), .A(D13935_Y));
KC_INV_X1 D14745 ( .Y(D14745_Y), .A(D14744_Y));
KC_INV_X1 D14735 ( .Y(D14735_Y), .A(D16398_Y));
KC_INV_X1 D14727 ( .Y(D14727_Y), .A(D818_Q));
KC_INV_X1 D14726 ( .Y(D14726_Y), .A(D14808_Q));
KC_INV_X1 D14725 ( .Y(D14725_Y), .A(D856_Q));
KC_INV_X1 D14720 ( .Y(D14720_Y), .A(D14514_Y));
KC_INV_X1 D14718 ( .Y(D14718_Y), .A(D14086_Y));
KC_INV_X1 D14710 ( .Y(D14710_Y), .A(D14705_Y));
KC_INV_X1 D14656 ( .Y(D14656_Y), .A(D15443_Y));
KC_INV_X1 D14655 ( .Y(D14655_Y), .A(D14753_Y));
KC_INV_X1 D14653 ( .Y(D14653_Y), .A(D645_Y));
KC_INV_X1 D14652 ( .Y(D14652_Y), .A(D14664_Y));
KC_INV_X1 D14651 ( .Y(D14651_Y), .A(D13958_Y));
KC_INV_X1 D14650 ( .Y(D14650_Y), .A(D13988_Y));
KC_INV_X1 D14643 ( .Y(D14643_Y), .A(D14688_Q));
KC_INV_X1 D14631 ( .Y(D14631_Y), .A(D14666_Y));
KC_INV_X1 D14630 ( .Y(D14630_Y), .A(D14689_Q));
KC_INV_X1 D14622 ( .Y(D14622_Y), .A(D14685_Q));
KC_INV_X1 D14619 ( .Y(D14619_Y), .A(D14686_Q));
KC_INV_X1 D14615 ( .Y(D14615_Y), .A(D14777_Y));
KC_INV_X1 D16769 ( .Y(D16769_Y), .A(D16770_Y));
KC_INV_X1 D14609 ( .Y(D14609_Y), .A(D14608_Y));
KC_INV_X1 D14607 ( .Y(D14607_Y), .A(D14606_Y));
KC_INV_X1 D14605 ( .Y(D14605_Y), .A(D14604_Y));
KC_INV_X1 D14603 ( .Y(D14603_Y), .A(D14602_Y));
KC_INV_X1 D14557 ( .Y(D14557_Y), .A(D14708_Y));
KC_INV_X1 D14553 ( .Y(D14553_Y), .A(D14518_Q));
KC_INV_X1 D14552 ( .Y(D14552_Y), .A(D608_Q));
KC_INV_X1 D14549 ( .Y(D14549_Y), .A(D14519_Q));
KC_INV_X1 D14548 ( .Y(D14548_Y), .A(D14567_Y));
KC_INV_X1 D14547 ( .Y(D14547_Y), .A(D14520_Q));
KC_INV_X1 D14543 ( .Y(D14543_Y), .A(D14601_Q));
KC_INV_X1 D14542 ( .Y(D14542_Y), .A(D14534_Y));
KC_INV_X1 D14535 ( .Y(D14535_Y), .A(D14519_Q));
KC_INV_X1 D14532 ( .Y(D14532_Y), .A(D14687_Q));
KC_INV_X1 D14531 ( .Y(D14531_Y), .A(D14805_Y));
KC_INV_X1 D14502 ( .Y(D14502_Y), .A(D14516_Y));
KC_INV_X1 D14501 ( .Y(D14501_Y), .A(D12173_Y));
KC_INV_X1 D14497 ( .Y(D14497_Y), .A(D9457_Y));
KC_INV_X1 D14486 ( .Y(D14486_Y), .A(D14495_Q));
KC_INV_X1 D14484 ( .Y(D14484_Y), .A(D14480_Y));
KC_INV_X1 D14481 ( .Y(D14481_Y), .A(D1401_Q));
KC_INV_X1 D14455 ( .Y(D14455_Y), .A(D14491_Q));
KC_INV_X1 D14454 ( .Y(D14454_Y), .A(D14410_Y));
KC_INV_X1 D14453 ( .Y(D14453_Y), .A(D15212_Q));
KC_INV_X1 D14441 ( .Y(D14441_Y), .A(D14446_Y));
KC_INV_X1 D14440 ( .Y(D14440_Y), .A(D1375_Q));
KC_INV_X1 D14439 ( .Y(D14439_Y), .A(D14432_Y));
KC_INV_X1 D14438 ( .Y(D14438_Y), .A(D15215_Q));
KC_INV_X1 D14431 ( .Y(D14431_Y), .A(D14427_Y));
KC_INV_X1 D14430 ( .Y(D14430_Y), .A(D14494_Q));
KC_INV_X1 D14424 ( .Y(D14424_Y), .A(D13808_Q));
KC_INV_X1 D14418 ( .Y(D14418_Y), .A(D1386_Q));
KC_INV_X1 D14417 ( .Y(D14417_Y), .A(D15216_Q));
KC_INV_X1 D14414 ( .Y(D14414_Y), .A(D14492_Q));
KC_INV_X1 D14413 ( .Y(D14413_Y), .A(D13826_Q));
KC_INV_X1 D14408 ( .Y(D14408_Y), .A(D1383_Q));
KC_INV_X1 D14407 ( .Y(D14407_Y), .A(D14406_Y));
KC_INV_X1 D14356 ( .Y(D14356_Y), .A(D1382_Q));
KC_INV_X1 D14350 ( .Y(D14350_Y), .A(D2523_Q));
KC_INV_X1 D14349 ( .Y(D14349_Y), .A(D14351_Y));
KC_INV_X1 D14348 ( .Y(D14348_Y), .A(D15234_Q));
KC_INV_X1 D14343 ( .Y(D14343_Y), .A(D15230_Q));
KC_INV_X1 D14336 ( .Y(D14336_Y), .A(D1182_Y));
KC_INV_X1 D14335 ( .Y(D14335_Y), .A(D14374_Q));
KC_INV_X1 D14222 ( .Y(D14222_Y), .A(D2515_Q));
KC_INV_X1 D14212 ( .Y(D14212_Y), .A(D14196_Q));
KC_INV_X1 D14204 ( .Y(D14204_Y), .A(D2626_Y));
KC_INV_X1 D14200 ( .Y(D14200_Y), .A(D14237_Q));
KC_INV_X1 D14138 ( .Y(D14138_Y), .A(D2502_Y));
KC_INV_X1 D14127 ( .Y(D14127_Y), .A(D14166_Q));
KC_INV_X1 D14108 ( .Y(D14108_Y), .A(D13986_Y));
KC_INV_X1 D14107 ( .Y(D14107_Y), .A(D16765_Y));
KC_INV_X1 D14106 ( .Y(D14106_Y), .A(D2514_Y));
KC_INV_X1 D14105 ( .Y(D14105_Y), .A(D13983_Y));
KC_INV_X1 D14104 ( .Y(D14104_Y), .A(D13984_Y));
KC_INV_X1 D14103 ( .Y(D14103_Y), .A(D13982_Y));
KC_INV_X1 D14047 ( .Y(D14047_Y), .A(D14046_Y));
KC_INV_X1 D14044 ( .Y(D14044_Y), .A(D13953_Y));
KC_INV_X1 D14030 ( .Y(D14030_Y), .A(D14002_Y));
KC_INV_X1 D14026 ( .Y(D14026_Y), .A(D13253_Y));
KC_INV_X1 D14025 ( .Y(D14025_Y), .A(D13330_Y));
KC_INV_X1 D14022 ( .Y(D14022_Y), .A(D14050_Y));
KC_INV_X1 D14021 ( .Y(D14021_Y), .A(D13985_Y));
KC_INV_X1 D14020 ( .Y(D14020_Y), .A(D16226_Q));
KC_INV_X1 D14019 ( .Y(D14019_Y), .A(D13321_Y));
KC_INV_X1 D14018 ( .Y(D14018_Y), .A(D14029_Y));
KC_INV_X1 D14017 ( .Y(D14017_Y), .A(D13977_Y));
KC_INV_X1 D14016 ( .Y(D14016_Y), .A(D14093_Q));
KC_INV_X1 D14011 ( .Y(D14011_Y), .A(D817_Q));
KC_INV_X1 D14010 ( .Y(D14010_Y), .A(D14116_Y));
KC_INV_X1 D13941 ( .Y(D13941_Y), .A(D573_Y));
KC_INV_X1 D13930 ( .Y(D13930_Y), .A(D13970_Y));
KC_INV_X1 D13925 ( .Y(D13925_Y), .A(D13924_Y));
KC_INV_X1 D13923 ( .Y(D13923_Y), .A(D13922_Y));
KC_INV_X1 D13874 ( .Y(D13874_Y), .A(D13873_Y));
KC_INV_X1 D13870 ( .Y(D13870_Y), .A(D13871_Y));
KC_INV_X1 D13869 ( .Y(D13869_Y), .A(D13868_Y));
KC_INV_X1 D13847 ( .Y(D13847_Y), .A(D13858_Y));
KC_INV_X1 D13846 ( .Y(D13846_Y), .A(D13846_A));
KC_INV_X1 D13779 ( .Y(D13779_Y), .A(D13806_Q));
KC_INV_X1 D13775 ( .Y(D13775_Y), .A(D13816_Q));
KC_INV_X1 D13774 ( .Y(D13774_Y), .A(D13827_Q));
KC_INV_X1 D13730 ( .Y(D13730_Y), .A(D14424_Y));
KC_INV_X1 D13729 ( .Y(D13729_Y), .A(D13812_Q));
KC_INV_X1 D13727 ( .Y(D13727_Y), .A(D14299_Q));
KC_INV_X1 D13719 ( .Y(D13719_Y), .A(D13759_Q));
KC_INV_X1 D13717 ( .Y(D13717_Y), .A(D13805_Q));
KC_INV_X1 D13716 ( .Y(D13716_Y), .A(D13813_Q));
KC_INV_X1 D13673 ( .Y(D13673_Y), .A(D14298_Q));
KC_INV_X1 D13672 ( .Y(D13672_Y), .A(D164_Q));
KC_INV_X1 D13671 ( .Y(D13671_Y), .A(D2474_Q));
KC_INV_X1 D13670 ( .Y(D13670_Y), .A(D13770_Q));
KC_INV_X1 D13666 ( .Y(D13666_Y), .A(D14240_Q));
KC_INV_X1 D13665 ( .Y(D13665_Y), .A(D14306_Q));
KC_INV_X1 D13664 ( .Y(D13664_Y), .A(D14303_Q));
KC_INV_X1 D13656 ( .Y(D13656_Y), .A(D14302_Q));
KC_INV_X1 D13655 ( .Y(D13655_Y), .A(D14307_Q));
KC_INV_X1 D13649 ( .Y(D13649_Y), .A(D13539_Y));
KC_INV_X1 D13646 ( .Y(D13646_Y), .A(D14316_Q));
KC_INV_X1 D13645 ( .Y(D13645_Y), .A(D14297_Q));
KC_INV_X1 D13579 ( .Y(D13579_Y), .A(D13552_Y));
KC_INV_X1 D13578 ( .Y(D13578_Y), .A(D13409_Y));
KC_INV_X1 D13572 ( .Y(D13572_Y), .A(D14220_Y));
KC_INV_X1 D13571 ( .Y(D13571_Y), .A(D13595_Y));
KC_INV_X1 D13570 ( .Y(D13570_Y), .A(D14247_Y));
KC_INV_X1 D13569 ( .Y(D13569_Y), .A(D13417_Y));
KC_INV_X1 D13567 ( .Y(D13567_Y), .A(D2430_Y));
KC_INV_X1 D13561 ( .Y(D13561_Y), .A(D13546_Y));
KC_INV_X1 D13560 ( .Y(D13560_Y), .A(D13580_Y));
KC_INV_X1 D13559 ( .Y(D13559_Y), .A(D13553_Y));
KC_INV_X1 D13558 ( .Y(D13558_Y), .A(D13586_Y));
KC_INV_X1 D13557 ( .Y(D13557_Y), .A(D13610_Y));
KC_INV_X1 D13556 ( .Y(D13556_Y), .A(D13554_Y));
KC_INV_X1 D13550 ( .Y(D13550_Y), .A(D13547_Y));
KC_INV_X1 D13549 ( .Y(D13549_Y), .A(D2436_Y));
KC_INV_X1 D13548 ( .Y(D13548_Y), .A(D13297_Y));
KC_INV_X1 D13544 ( .Y(D13544_Y), .A(D13538_Y));
KC_INV_X1 D13543 ( .Y(D13543_Y), .A(D13295_Y));
KC_INV_X1 D13534 ( .Y(D13534_Y), .A(D13447_Y));
KC_INV_X1 D13479 ( .Y(D13479_Y), .A(D984_Y));
KC_INV_X1 D13478 ( .Y(D13478_Y), .A(D13322_Y));
KC_INV_X1 D13477 ( .Y(D13477_Y), .A(D13410_Y));
KC_INV_X1 D13476 ( .Y(D13476_Y), .A(D13314_Y));
KC_INV_X1 D13475 ( .Y(D13475_Y), .A(D13316_Y));
KC_INV_X1 D13474 ( .Y(D13474_Y), .A(D13329_Y));
KC_INV_X1 D13473 ( .Y(D13473_Y), .A(D13317_Y));
KC_INV_X1 D13472 ( .Y(D13472_Y), .A(D13312_Y));
KC_INV_X1 D13469 ( .Y(D13469_Y), .A(D13515_Q));
KC_INV_X1 D13468 ( .Y(D13468_Y), .A(D2394_Y));
KC_INV_X1 D13467 ( .Y(D13467_Y), .A(D13513_Y));
KC_INV_X1 D13466 ( .Y(D13466_Y), .A(D2433_Y));
KC_INV_X1 D13461 ( .Y(D13461_Y), .A(D13456_Y));
KC_INV_X1 D13460 ( .Y(D13460_Y), .A(D13448_Y));
KC_INV_X1 D13459 ( .Y(D13459_Y), .A(D13507_Y));
KC_INV_X1 D13458 ( .Y(D13458_Y), .A(D2429_Y));
KC_INV_X1 D13457 ( .Y(D13457_Y), .A(D13502_Y));
KC_INV_X1 D13451 ( .Y(D13451_Y), .A(D13505_Y));
KC_INV_X1 D13450 ( .Y(D13450_Y), .A(D13428_Y));
KC_INV_X1 D13449 ( .Y(D13449_Y), .A(D13445_Y));
KC_INV_X1 D13437 ( .Y(D13437_Y), .A(D15694_Y));
KC_INV_X1 D13436 ( .Y(D13436_Y), .A(D15583_Y));
KC_INV_X1 D13430 ( .Y(D13430_Y), .A(D886_Y));
KC_INV_X1 D13423 ( .Y(D13423_Y), .A(D13540_Y));
KC_INV_X1 D13422 ( .Y(D13422_Y), .A(D13429_Y));
KC_INV_X1 D13421 ( .Y(D13421_Y), .A(D13393_Y));
KC_INV_X1 D13359 ( .Y(D13359_Y), .A(D13221_Y));
KC_INV_X1 D13358 ( .Y(D13358_Y), .A(D13269_Q));
KC_INV_X1 D13357 ( .Y(D13357_Y), .A(D13397_Q));
KC_INV_X1 D13349 ( .Y(D13349_Y), .A(D13343_Y));
KC_INV_X1 D13348 ( .Y(D13348_Y), .A(D14024_Y));
KC_INV_X1 D13347 ( .Y(D13347_Y), .A(D13398_Q));
KC_INV_X1 D13346 ( .Y(D13346_Y), .A(D13396_Q));
KC_INV_X1 D13333 ( .Y(D13333_Y), .A(D13339_Y));
KC_INV_X1 D13332 ( .Y(D13332_Y), .A(D12822_Y));
KC_INV_X1 D13323 ( .Y(D13323_Y), .A(D13338_Y));
KC_INV_X1 D13309 ( .Y(D13309_Y), .A(D13318_Y));
KC_INV_X1 D13302 ( .Y(D13302_Y), .A(D12277_Q));
KC_INV_X1 D13236 ( .Y(D13236_Y), .A(D7609_Y));
KC_INV_X1 D13234 ( .Y(D13234_Y), .A(D7609_Y));
KC_INV_X1 D13231 ( .Y(D13231_Y), .A(D13241_Y));
KC_INV_X1 D13228 ( .Y(D13228_Y), .A(D12296_Y));
KC_INV_X1 D13227 ( .Y(D13227_Y), .A(D12739_Y));
KC_INV_X1 D13226 ( .Y(D13226_Y), .A(D12298_Y));
KC_INV_X1 D13225 ( .Y(D13225_Y), .A(D12254_Y));
KC_INV_X1 D13220 ( .Y(D13220_Y), .A(D13252_Y));
KC_INV_X1 D13179 ( .Y(D13179_Y), .A(D13235_Y));
KC_INV_X1 D13178 ( .Y(D13178_Y), .A(D13213_Q));
KC_INV_X1 D16764 ( .Y(D16764_Y), .A(D16763_Y));
KC_INV_X1 D13015 ( .Y(D13015_Y), .A(D956_Q));
KC_INV_X1 D13010 ( .Y(D13010_Y), .A(D13442_Y));
KC_INV_X1 D12960 ( .Y(D12960_Y), .A(D2372_Y));
KC_INV_X1 D12952 ( .Y(D12952_Y), .A(D12930_Y));
KC_INV_X1 D12951 ( .Y(D12951_Y), .A(D13536_Y));
KC_INV_X1 D12947 ( .Y(D12947_Y), .A(D13454_Y));
KC_INV_X1 D12942 ( .Y(D12942_Y), .A(D12889_Y));
KC_INV_X1 D12941 ( .Y(D12941_Y), .A(D12872_Y));
KC_INV_X1 D12893 ( .Y(D12893_Y), .A(D2401_Y));
KC_INV_X1 D12890 ( .Y(D12890_Y), .A(D12888_Y));
KC_INV_X1 D12879 ( .Y(D12879_Y), .A(D961_Y));
KC_INV_X1 D12878 ( .Y(D12878_Y), .A(D12926_Q));
KC_INV_X1 D12876 ( .Y(D12876_Y), .A(D929_Q));
KC_INV_X1 D12870 ( .Y(D12870_Y), .A(D12932_Y));
KC_INV_X1 D12868 ( .Y(D12868_Y), .A(D12770_Y));
KC_INV_X1 D12865 ( .Y(D12865_Y), .A(D12823_Y));
KC_INV_X1 D12815 ( .Y(D12815_Y), .A(D13370_Y));
KC_INV_X1 D12814 ( .Y(D12814_Y), .A(D12753_Q));
KC_INV_X1 D12813 ( .Y(D12813_Y), .A(D12754_Q));
KC_INV_X1 D12810 ( .Y(D12810_Y), .A(D15491_Y));
KC_INV_X1 D12809 ( .Y(D12809_Y), .A(D12749_Q));
KC_INV_X1 D12806 ( .Y(D12806_Y), .A(D12808_Y));
KC_INV_X1 D12805 ( .Y(D12805_Y), .A(D12804_Y));
KC_INV_X1 D12800 ( .Y(D12800_Y), .A(D843_Q));
KC_INV_X1 D12799 ( .Y(D12799_Y), .A(D12854_Q));
KC_INV_X1 D12798 ( .Y(D12798_Y), .A(D12857_Q));
KC_INV_X1 D12795 ( .Y(D12795_Y), .A(D15474_Y));
KC_INV_X1 D12794 ( .Y(D12794_Y), .A(D12858_Q));
KC_INV_X1 D12788 ( .Y(D12788_Y), .A(D14730_Y));
KC_INV_X1 D12787 ( .Y(D12787_Y), .A(D15498_Y));
KC_INV_X1 D12786 ( .Y(D12786_Y), .A(D12866_Y));
KC_INV_X1 D12773 ( .Y(D12773_Y), .A(D12855_Q));
KC_INV_X1 D12772 ( .Y(D12772_Y), .A(D146_Q));
KC_INV_X1 D12769 ( .Y(D12769_Y), .A(D12748_Q));
KC_INV_X1 D12767 ( .Y(D12767_Y), .A(D12719_Y));
KC_INV_X1 D12757 ( .Y(D12757_Y), .A(D2363_Y));
KC_INV_X1 D12718 ( .Y(D12718_Y), .A(D12250_Y));
KC_INV_X1 D12716 ( .Y(D12716_Y), .A(D12755_Q));
KC_INV_X1 D12715 ( .Y(D12715_Y), .A(D12752_Q));
KC_INV_X1 D12714 ( .Y(D12714_Y), .A(D12204_Y));
KC_INV_X1 D12712 ( .Y(D12712_Y), .A(D12713_Y));
KC_INV_X1 D12704 ( .Y(D12704_Y), .A(D12725_Y));
KC_INV_X1 D12703 ( .Y(D12703_Y), .A(D12753_Q));
KC_INV_X1 D12658 ( .Y(D12658_Y), .A(D2360_Y));
KC_INV_X1 D12326 ( .Y(D12326_Y), .A(D12699_Y));
KC_INV_X1 D12325 ( .Y(D12325_Y), .A(D716_Q));
KC_INV_X1 D12322 ( .Y(D12322_Y), .A(D12869_Y));
KC_INV_X1 D12321 ( .Y(D12321_Y), .A(D12351_Q));
KC_INV_X1 D12320 ( .Y(D12320_Y), .A(D1814_Y));
KC_INV_X1 D12319 ( .Y(D12319_Y), .A(D6410_Y));
KC_INV_X1 D12318 ( .Y(D12318_Y), .A(D12782_Y));
KC_INV_X1 D12317 ( .Y(D12317_Y), .A(D12771_Y));
KC_INV_X1 D12316 ( .Y(D12316_Y), .A(D14057_Y));
KC_INV_X1 D12315 ( .Y(D12315_Y), .A(D12779_Y));
KC_INV_X1 D12314 ( .Y(D12314_Y), .A(D12344_Q));
KC_INV_X1 D12309 ( .Y(D12309_Y), .A(D12341_Q));
KC_INV_X1 D12299 ( .Y(D12299_Y), .A(D12211_Y));
KC_INV_X1 D12248 ( .Y(D12248_Y), .A(D717_Q));
KC_INV_X1 D12243 ( .Y(D12243_Y), .A(D13400_Y));
KC_INV_X1 D12201 ( .Y(D12201_Y), .A(D558_Y));
KC_INV_X1 D12200 ( .Y(D12200_Y), .A(D10134_Y));
KC_INV_X1 D12197 ( .Y(D12197_Y), .A(D12141_Y));
KC_INV_X1 D12192 ( .Y(D12192_Y), .A(D12193_Y));
KC_INV_X1 D12191 ( .Y(D12191_Y), .A(D12198_Y));
KC_INV_X1 D12132 ( .Y(D12132_Y), .A(D12178_Q));
KC_INV_X1 D12131 ( .Y(D12131_Y), .A(D548_Q));
KC_INV_X1 D12059 ( .Y(D12059_Y), .A(D13074_Y));
KC_INV_X1 D12028 ( .Y(D12028_Y), .A(D11990_Y));
KC_INV_X1 D12017 ( .Y(D12017_Y), .A(D11957_Y));
KC_INV_X1 D12013 ( .Y(D12013_Y), .A(D12027_Y));
KC_INV_X1 D12006 ( .Y(D12006_Y), .A(D13058_Y));
KC_INV_X1 D12000 ( .Y(D12000_Y), .A(D13072_Y));
KC_INV_X1 D11955 ( .Y(D11955_Y), .A(D11945_Y));
KC_INV_X1 D11954 ( .Y(D11954_Y), .A(D11969_Y));
KC_INV_X1 D11946 ( .Y(D11946_Y), .A(D11941_Y));
KC_INV_X1 D11842 ( .Y(D11842_Y), .A(D12375_Y));
KC_INV_X1 D11738 ( .Y(D11738_Y), .A(D11753_Y));
KC_INV_X1 D11737 ( .Y(D11737_Y), .A(D11770_Y));
KC_INV_X1 D11678 ( .Y(D11678_Y), .A(D11670_Y));
KC_INV_X1 D11646 ( .Y(D11646_Y), .A(D11648_Y));
KC_INV_X1 D11614 ( .Y(D11614_Y), .A(D8_Y));
KC_INV_X1 D11505 ( .Y(D11505_Y), .A(D10861_Y));
KC_INV_X1 D11504 ( .Y(D11504_Y), .A(D12022_Y));
KC_INV_X1 D11499 ( .Y(D11499_Y), .A(D12538_Y));
KC_INV_X1 D11494 ( .Y(D11494_Y), .A(D13103_Y));
KC_INV_X1 D11493 ( .Y(D11493_Y), .A(D12570_Y));
KC_INV_X1 D11492 ( .Y(D11492_Y), .A(D12004_Y));
KC_INV_X1 D11491 ( .Y(D11491_Y), .A(D12537_Y));
KC_INV_X1 D11490 ( .Y(D11490_Y), .A(D12517_Y));
KC_INV_X1 D11488 ( .Y(D11488_Y), .A(D12568_Y));
KC_INV_X1 D11484 ( .Y(D11484_Y), .A(D13057_Y));
KC_INV_X1 D11483 ( .Y(D11483_Y), .A(D1264_Y));
KC_INV_X1 D11481 ( .Y(D11481_Y), .A(D12061_Y));
KC_INV_X1 D11479 ( .Y(D11479_Y), .A(D12070_Y));
KC_INV_X1 D11432 ( .Y(D11432_Y), .A(D12492_Y));
KC_INV_X1 D11431 ( .Y(D11431_Y), .A(D2269_Y));
KC_INV_X1 D11426 ( .Y(D11426_Y), .A(D12489_Y));
KC_INV_X1 D11425 ( .Y(D11425_Y), .A(D12484_Y));
KC_INV_X1 D11421 ( .Y(D11421_Y), .A(D11438_Y));
KC_INV_X1 D11419 ( .Y(D11419_Y), .A(D12436_Y));
KC_INV_X1 D11372 ( .Y(D11372_Y), .A(D11947_Y));
KC_INV_X1 D11366 ( .Y(D11366_Y), .A(D12439_Y));
KC_INV_X1 D11354 ( .Y(D11354_Y), .A(D12491_Y));
KC_INV_X1 D11302 ( .Y(D11302_Y), .A(D11834_Y));
KC_INV_X1 D11297 ( .Y(D11297_Y), .A(D11878_Y));
KC_INV_X1 D11296 ( .Y(D11296_Y), .A(D12391_Y));
KC_INV_X1 D11295 ( .Y(D11295_Y), .A(D2276_Y));
KC_INV_X1 D11288 ( .Y(D11288_Y), .A(D11837_Y));
KC_INV_X1 D11287 ( .Y(D11287_Y), .A(D12423_Y));
KC_INV_X1 D11228 ( .Y(D11228_Y), .A(D1813_Y));
KC_INV_X1 D11212 ( .Y(D11212_Y), .A(D463_Y));
KC_INV_X1 D11210 ( .Y(D11210_Y), .A(D11697_Y));
KC_INV_X1 D11209 ( .Y(D11209_Y), .A(D11699_Y));
KC_INV_X1 D11205 ( .Y(D11205_Y), .A(D11222_Y));
KC_INV_X1 D11204 ( .Y(D11204_Y), .A(D10675_Y));
KC_INV_X1 D11200 ( .Y(D11200_Y), .A(D10754_Y));
KC_INV_X1 D11194 ( .Y(D11194_Y), .A(D11214_Y));
KC_INV_X1 D11192 ( .Y(D11192_Y), .A(D11754_Y));
KC_INV_X1 D11146 ( .Y(D11146_Y), .A(D10192_Y));
KC_INV_X1 D11091 ( .Y(D11091_Y), .A(D11101_Y));
KC_INV_X1 D10980 ( .Y(D10980_Y), .A(D11428_Y));
KC_INV_X1 D10964 ( .Y(D10964_Y), .A(D10963_Y));
KC_INV_X1 D10936 ( .Y(D10936_Y), .A(D10972_Y));
KC_INV_X1 D10905 ( .Y(D10905_Y), .A(D10967_Y));
KC_INV_X1 D10858 ( .Y(D10858_Y), .A(D5339_Y));
KC_INV_X1 D10849 ( .Y(D10849_Y), .A(D10856_Y));
KC_INV_X1 D10751 ( .Y(D10751_Y), .A(D7824_Y));
KC_INV_X1 D10748 ( .Y(D10748_Y), .A(D7974_Y));
KC_INV_X1 D10747 ( .Y(D10747_Y), .A(D10729_Y));
KC_INV_X1 D10746 ( .Y(D10746_Y), .A(D10306_Q));
KC_INV_X1 D10744 ( .Y(D10744_Y), .A(D10699_Y));
KC_INV_X1 D10741 ( .Y(D10741_Y), .A(D10760_Y));
KC_INV_X1 D10735 ( .Y(D10735_Y), .A(D10295_Q));
KC_INV_X1 D10732 ( .Y(D10732_Y), .A(D10308_Q));
KC_INV_X1 D10701 ( .Y(D10701_Y), .A(D1964_Y));
KC_INV_X1 D10681 ( .Y(D10681_Y), .A(D6406_Y));
KC_INV_X1 D10664 ( .Y(D10664_Y), .A(D10734_Y));
KC_INV_X1 D10536 ( .Y(D10536_Y), .A(D10965_Y));
KC_INV_X1 D10466 ( .Y(D10466_Y), .A(D10513_Q));
KC_INV_X1 D10464 ( .Y(D10464_Y), .A(D10515_Q));
KC_INV_X1 D10460 ( .Y(D10460_Y), .A(D10509_Q));
KC_INV_X1 D10459 ( .Y(D10459_Y), .A(D1127_Q));
KC_INV_X1 D10458 ( .Y(D10458_Y), .A(D10508_Q));
KC_INV_X1 D10455 ( .Y(D10455_Y), .A(D2131_Y));
KC_INV_X1 D10454 ( .Y(D10454_Y), .A(D10470_Y));
KC_INV_X1 D10453 ( .Y(D10453_Y), .A(D10531_Y));
KC_INV_X1 D10452 ( .Y(D10452_Y), .A(D2157_Q));
KC_INV_X1 D10451 ( .Y(D10451_Y), .A(D1123_Q));
KC_INV_X1 D10447 ( .Y(D10447_Y), .A(D116_Q));
KC_INV_X1 D10446 ( .Y(D10446_Y), .A(D10579_Y));
KC_INV_X1 D10408 ( .Y(D10408_Y), .A(D10908_Y));
KC_INV_X1 D10407 ( .Y(D10407_Y), .A(D10901_Y));
KC_INV_X1 D10389 ( .Y(D10389_Y), .A(D2200_Y));
KC_INV_X1 D10388 ( .Y(D10388_Y), .A(D10962_Y));
KC_INV_X1 D10321 ( .Y(D10321_Y), .A(D10366_Q));
KC_INV_X1 D10320 ( .Y(D10320_Y), .A(D8295_Y));
KC_INV_X1 D10319 ( .Y(D10319_Y), .A(D10360_Q));
KC_INV_X1 D10248 ( .Y(D10248_Y), .A(D2155_Y));
KC_INV_X1 D10247 ( .Y(D10247_Y), .A(D10302_Q));
KC_INV_X1 D10246 ( .Y(D10246_Y), .A(D10301_Q));
KC_INV_X1 D10244 ( .Y(D10244_Y), .A(D10299_Q));
KC_INV_X1 D10243 ( .Y(D10243_Y), .A(D10294_Q));
KC_INV_X1 D10241 ( .Y(D10241_Y), .A(D10305_Q));
KC_INV_X1 D10201 ( .Y(D10201_Y), .A(D462_Y));
KC_INV_X1 D10197 ( .Y(D10197_Y), .A(D9472_Q));
KC_INV_X1 D10196 ( .Y(D10196_Y), .A(D702_Q));
KC_INV_X1 D10179 ( .Y(D10179_Y), .A(D6285_Y));
KC_INV_X1 D10178 ( .Y(D10178_Y), .A(D6407_Y));
KC_INV_X1 D10177 ( .Y(D10177_Y), .A(D6287_Y));
KC_INV_X1 D10152 ( .Y(D10152_Y), .A(D9983_Q));
KC_INV_X1 D10137 ( .Y(D10137_Y), .A(D11114_Y));
KC_INV_X1 D10134 ( .Y(D10134_Y), .A(D7527_Y));
KC_INV_X1 D10130 ( .Y(D10130_Y), .A(D10086_Y));
KC_INV_X1 D10128 ( .Y(D10128_Y), .A(D10047_Q));
KC_INV_X1 D10125 ( .Y(D10125_Y), .A(D10051_Q));
KC_INV_X1 D10123 ( .Y(D10123_Y), .A(D10032_Q));
KC_INV_X1 D10120 ( .Y(D10120_Y), .A(D10009_Q));
KC_INV_X1 D10118 ( .Y(D10118_Y), .A(D2166_Q));
KC_INV_X1 D10102 ( .Y(D10102_Y), .A(D10072_Y));
KC_INV_X1 D10096 ( .Y(D10096_Y), .A(D10116_Y));
KC_INV_X1 D10082 ( .Y(D10082_Y), .A(D9104_Y));
KC_INV_X1 D10081 ( .Y(D10081_Y), .A(D10087_Y));
KC_INV_X1 D10076 ( .Y(D10076_Y), .A(D419_Q));
KC_INV_X1 D10071 ( .Y(D10071_Y), .A(D9218_Q));
KC_INV_X1 D10066 ( .Y(D10066_Y), .A(D11623_Y));
KC_INV_X1 D10052 ( .Y(D10052_Y), .A(D10062_Q));
KC_INV_X1 D10039 ( .Y(D10039_Y), .A(D10031_Q));
KC_INV_X1 D10000 ( .Y(D10000_Y), .A(D10007_Q));
KC_INV_X1 D9996 ( .Y(D9996_Y), .A(D8901_Y));
KC_INV_X1 D9990 ( .Y(D9990_Y), .A(D7407_Y));
KC_INV_X1 D9968 ( .Y(D9968_Y), .A(D9959_Y));
KC_INV_X1 D9961 ( .Y(D9961_Y), .A(D7882_Y));
KC_INV_X1 D9960 ( .Y(D9960_Y), .A(D8702_Y));
KC_INV_X1 D9928 ( .Y(D9928_Y), .A(D9967_Y));
KC_INV_X1 D9927 ( .Y(D9927_Y), .A(D8697_Y));
KC_INV_X1 D9926 ( .Y(D9926_Y), .A(D9940_Y));
KC_INV_X1 D9924 ( .Y(D9924_Y), .A(D9941_Q));
KC_INV_X1 D9923 ( .Y(D9923_Y), .A(D9950_Q));
KC_INV_X1 D9830 ( .Y(D9830_Y), .A(D10569_Y));
KC_INV_X1 D9752 ( .Y(D9752_Y), .A(D9784_Q));
KC_INV_X1 D9750 ( .Y(D9750_Y), .A(D2079_Q));
KC_INV_X1 D9746 ( .Y(D9746_Y), .A(D2032_Y));
KC_INV_X1 D9744 ( .Y(D9744_Y), .A(D9785_Q));
KC_INV_X1 D9743 ( .Y(D9743_Y), .A(D10585_Y));
KC_INV_X1 D9742 ( .Y(D9742_Y), .A(D1131_Q));
KC_INV_X1 D9741 ( .Y(D9741_Y), .A(D9791_Q));
KC_INV_X1 D9740 ( .Y(D9740_Y), .A(D9792_Q));
KC_INV_X1 D9739 ( .Y(D9739_Y), .A(D10521_Y));
KC_INV_X1 D9738 ( .Y(D9738_Y), .A(D10591_Y));
KC_INV_X1 D9737 ( .Y(D9737_Y), .A(D9820_Y));
KC_INV_X1 D9736 ( .Y(D9736_Y), .A(D9793_Q));
KC_INV_X1 D9735 ( .Y(D9735_Y), .A(D9823_Y));
KC_INV_X1 D9733 ( .Y(D9733_Y), .A(D9790_Q));
KC_INV_X1 D9728 ( .Y(D9728_Y), .A(D9874_Y));
KC_INV_X1 D9727 ( .Y(D9727_Y), .A(D9839_Q));
KC_INV_X1 D9726 ( .Y(D9726_Y), .A(D9789_Q));
KC_INV_X1 D9683 ( .Y(D9683_Y), .A(D9661_Y));
KC_INV_X1 D9682 ( .Y(D9682_Y), .A(D9787_Q));
KC_INV_X1 D9681 ( .Y(D9681_Y), .A(D9788_Q));
KC_INV_X1 D9672 ( .Y(D9672_Y), .A(D1895_Y));
KC_INV_X1 D9648 ( .Y(D9648_Y), .A(D10935_Y));
KC_INV_X1 D9647 ( .Y(D9647_Y), .A(D10376_Y));
KC_INV_X1 D9646 ( .Y(D9646_Y), .A(D10384_Y));
KC_INV_X1 D9645 ( .Y(D9645_Y), .A(D9704_Q));
KC_INV_X1 D9644 ( .Y(D9644_Y), .A(D10391_Y));
KC_INV_X1 D9643 ( .Y(D9643_Y), .A(D9786_Q));
KC_INV_X1 D9642 ( .Y(D9642_Y), .A(D10400_Y));
KC_INV_X1 D9641 ( .Y(D9641_Y), .A(D9667_Y));
KC_INV_X1 D9640 ( .Y(D9640_Y), .A(D9671_Y));
KC_INV_X1 D9597 ( .Y(D9597_Y), .A(D9574_Q));
KC_INV_X1 D9536 ( .Y(D9536_Y), .A(D643_Y));
KC_INV_X1 D9535 ( .Y(D9535_Y), .A(D826_Q));
KC_INV_X1 D9528 ( .Y(D9528_Y), .A(D9576_Q));
KC_INV_X1 D9524 ( .Y(D9524_Y), .A(D9542_Y));
KC_INV_X1 D9522 ( .Y(D9522_Y), .A(D9578_Q));
KC_INV_X1 D9521 ( .Y(D9521_Y), .A(D9575_Q));
KC_INV_X1 D9516 ( .Y(D9516_Y), .A(D9583_Y));
KC_INV_X1 D9514 ( .Y(D9514_Y), .A(D9579_Q));
KC_INV_X1 D9513 ( .Y(D9513_Y), .A(D9577_Q));
KC_INV_X1 D9512 ( .Y(D9512_Y), .A(D9506_Y));
KC_INV_X1 D9511 ( .Y(D9511_Y), .A(D9532_Y));
KC_INV_X1 D9504 ( .Y(D9504_Y), .A(D2108_Y));
KC_INV_X1 D9503 ( .Y(D9503_Y), .A(D9584_Y));
KC_INV_X1 D9499 ( .Y(D9499_Y), .A(D2039_Y));
KC_INV_X1 D9494 ( .Y(D9494_Y), .A(D933_Q));
KC_INV_X1 D9425 ( .Y(D9425_Y), .A(D704_Q));
KC_INV_X1 D9424 ( .Y(D9424_Y), .A(D10225_Q));
KC_INV_X1 D9423 ( .Y(D9423_Y), .A(D9581_Q));
KC_INV_X1 D9422 ( .Y(D9422_Y), .A(D10226_Q));
KC_INV_X1 D9421 ( .Y(D9421_Y), .A(D9473_Y));
KC_INV_X1 D9419 ( .Y(D9419_Y), .A(D9488_Q));
KC_INV_X1 D9415 ( .Y(D9415_Y), .A(D9580_Q));
KC_INV_X1 D9414 ( .Y(D9414_Y), .A(D701_Q));
KC_INV_X1 D9413 ( .Y(D9413_Y), .A(D703_Q));
KC_INV_X1 D9407 ( .Y(D9407_Y), .A(D8221_Y));
KC_INV_X1 D9406 ( .Y(D9406_Y), .A(D9470_Q));
KC_INV_X1 D9400 ( .Y(D9400_Y), .A(D7402_Y));
KC_INV_X1 D9399 ( .Y(D9399_Y), .A(D8220_Y));
KC_INV_X1 D9395 ( .Y(D9395_Y), .A(D10211_Y));
KC_INV_X1 D9394 ( .Y(D9394_Y), .A(D9398_Y));
KC_INV_X1 D9371 ( .Y(D9371_Y), .A(D6288_Y));
KC_INV_X1 D9366 ( .Y(D9366_Y), .A(D9370_Y));
KC_INV_X1 D9342 ( .Y(D9342_Y), .A(D155_Q));
KC_INV_X1 D9341 ( .Y(D9341_Y), .A(D1924_Y));
KC_INV_X1 D9306 ( .Y(D9306_Y), .A(D490_Y));
KC_INV_X1 D9300 ( .Y(D9300_Y), .A(D9299_Y));
KC_INV_X1 D9243 ( .Y(D9243_Y), .A(D2003_Y));
KC_INV_X1 D9236 ( .Y(D9236_Y), .A(D465_Y));
KC_INV_X1 D9235 ( .Y(D9235_Y), .A(D9275_Q));
KC_INV_X1 D9234 ( .Y(D9234_Y), .A(D9285_Y));
KC_INV_X1 D9186 ( .Y(D9186_Y), .A(D7638_Y));
KC_INV_X1 D9181 ( .Y(D9181_Y), .A(D7643_Y));
KC_INV_X1 D9168 ( .Y(D9168_Y), .A(D7136_Y));
KC_INV_X1 D9166 ( .Y(D9166_Y), .A(D7497_Y));
KC_INV_X1 D9122 ( .Y(D9122_Y), .A(D36_Y));
KC_INV_X1 D9120 ( .Y(D9120_Y), .A(D15450_Y));
KC_INV_X1 D9118 ( .Y(D9118_Y), .A(D273_Y));
KC_INV_X1 D9115 ( .Y(D9115_Y), .A(D7631_Y));
KC_INV_X1 D9114 ( .Y(D9114_Y), .A(D7644_Y));
KC_INV_X1 D9109 ( .Y(D9109_Y), .A(D9099_Y));
KC_INV_X1 D9108 ( .Y(D9108_Y), .A(D385_Q));
KC_INV_X1 D9102 ( .Y(D9102_Y), .A(D1904_Y));
KC_INV_X1 D9059 ( .Y(D9059_Y), .A(D8970_Y));
KC_INV_X1 D9057 ( .Y(D9057_Y), .A(D40_Q));
KC_INV_X1 D9056 ( .Y(D9056_Y), .A(D41_Y));
KC_INV_X1 D9041 ( .Y(D9041_Y), .A(D7510_Y));
KC_INV_X1 D9033 ( .Y(D9033_Y), .A(D8951_Q));
KC_INV_X1 D8986 ( .Y(D8986_Y), .A(D1880_Y));
KC_INV_X1 D8985 ( .Y(D8985_Y), .A(D57_Y));
KC_INV_X1 D8980 ( .Y(D8980_Y), .A(D7315_Y));
KC_INV_X1 D8976 ( .Y(D8976_Y), .A(D9025_Y));
KC_INV_X1 D8973 ( .Y(D8973_Y), .A(D8899_Q));
KC_INV_X1 D8972 ( .Y(D8972_Y), .A(D8824_Q));
KC_INV_X1 D8971 ( .Y(D8971_Y), .A(D9019_Q));
KC_INV_X1 D8917 ( .Y(D8917_Y), .A(D1907_Y));
KC_INV_X1 D8908 ( .Y(D8908_Y), .A(D334_Q));
KC_INV_X1 D8904 ( .Y(D8904_Y), .A(D8954_Q));
KC_INV_X1 D8877 ( .Y(D8877_Y), .A(D9482_Y));
KC_INV_X1 D8865 ( .Y(D8865_Y), .A(D5710_Y));
KC_INV_X1 D8861 ( .Y(D8861_Y), .A(D12176_Y));
KC_INV_X1 D8851 ( .Y(D8851_Y), .A(D2070_Y));
KC_INV_X1 D8844 ( .Y(D8844_Y), .A(D2029_Y));
KC_INV_X1 D8840 ( .Y(D8840_Y), .A(D8811_Y));
KC_INV_X1 D8839 ( .Y(D8839_Y), .A(D8822_Q));
KC_INV_X1 D8769 ( .Y(D8769_Y), .A(D227_Q));
KC_INV_X1 D8767 ( .Y(D8767_Y), .A(D233_Q));
KC_INV_X1 D8760 ( .Y(D8760_Y), .A(D8781_Y));
KC_INV_X1 D8759 ( .Y(D8759_Y), .A(D8737_Y));
KC_INV_X1 D8757 ( .Y(D8757_Y), .A(D8782_Y));
KC_INV_X1 D8756 ( .Y(D8756_Y), .A(D2095_Y));
KC_INV_X1 D8751 ( .Y(D8751_Y), .A(D8876_Y));
KC_INV_X1 D8749 ( .Y(D8749_Y), .A(D9479_Y));
KC_INV_X1 D8748 ( .Y(D8748_Y), .A(D9477_Y));
KC_INV_X1 D8744 ( .Y(D8744_Y), .A(D2026_Y));
KC_INV_X1 D8743 ( .Y(D8743_Y), .A(D204_Y));
KC_INV_X1 D8738 ( .Y(D8738_Y), .A(D201_Y));
KC_INV_X1 D8676 ( .Y(D8676_Y), .A(D8768_Y));
KC_INV_X1 D8675 ( .Y(D8675_Y), .A(D8688_Y));
KC_INV_X1 D8671 ( .Y(D8671_Y), .A(D8685_Y));
KC_INV_X1 D8669 ( .Y(D8669_Y), .A(D8712_Q));
KC_INV_X1 D8666 ( .Y(D8666_Y), .A(D8665_Y));
KC_INV_X1 D8665 ( .Y(D8665_Y), .A(D2055_Y));
KC_INV_X1 D8564 ( .Y(D8564_Y), .A(D8595_Q));
KC_INV_X1 D8561 ( .Y(D8561_Y), .A(D7039_Y));
KC_INV_X1 D8559 ( .Y(D8559_Y), .A(D10565_Y));
KC_INV_X1 D8558 ( .Y(D8558_Y), .A(D5547_Y));
KC_INV_X1 D8504 ( .Y(D8504_Y), .A(D8545_Q));
KC_INV_X1 D8503 ( .Y(D8503_Y), .A(D1929_Q));
KC_INV_X1 D8502 ( .Y(D8502_Y), .A(D8534_Y));
KC_INV_X1 D8501 ( .Y(D8501_Y), .A(D8544_Q));
KC_INV_X1 D8499 ( .Y(D8499_Y), .A(D8500_Y));
KC_INV_X1 D8498 ( .Y(D8498_Y), .A(D8500_Y));
KC_INV_X1 D8497 ( .Y(D8497_Y), .A(D8546_Q));
KC_INV_X1 D8494 ( .Y(D8494_Y), .A(D8547_Q));
KC_INV_X1 D8493 ( .Y(D8493_Y), .A(D8548_Q));
KC_INV_X1 D8492 ( .Y(D8492_Y), .A(D8549_Q));
KC_INV_X1 D8488 ( .Y(D8488_Y), .A(D8541_Q));
KC_INV_X1 D8487 ( .Y(D8487_Y), .A(D9871_Y));
KC_INV_X1 D8485 ( .Y(D8485_Y), .A(D1255_Y));
KC_INV_X1 D8484 ( .Y(D8484_Y), .A(D9822_Y));
KC_INV_X1 D8482 ( .Y(D8482_Y), .A(D8539_Q));
KC_INV_X1 D8481 ( .Y(D8481_Y), .A(D115_Q));
KC_INV_X1 D8477 ( .Y(D8477_Y), .A(D5420_Y));
KC_INV_X1 D8424 ( .Y(D8424_Y), .A(D8543_Q));
KC_INV_X1 D8423 ( .Y(D8423_Y), .A(D9660_Y));
KC_INV_X1 D8422 ( .Y(D8422_Y), .A(D545_Y));
KC_INV_X1 D8421 ( .Y(D8421_Y), .A(D6847_Y));
KC_INV_X1 D8420 ( .Y(D8420_Y), .A(D6859_Y));
KC_INV_X1 D8414 ( .Y(D8414_Y), .A(D8419_Y));
KC_INV_X1 D8405 ( .Y(D8405_Y), .A(D1837_Y));
KC_INV_X1 D8404 ( .Y(D8404_Y), .A(D3916_Y));
KC_INV_X1 D8395 ( .Y(D8395_Y), .A(D545_Y));
KC_INV_X1 D8394 ( .Y(D8394_Y), .A(D8392_Y));
KC_INV_X1 D8388 ( .Y(D8388_Y), .A(D8368_Y));
KC_INV_X1 D8387 ( .Y(D8387_Y), .A(D8369_Y));
KC_INV_X1 D8366 ( .Y(D8366_Y), .A(D8458_Q));
KC_INV_X1 D8365 ( .Y(D8365_Y), .A(D545_Y));
KC_INV_X1 D8364 ( .Y(D8364_Y), .A(D11024_Y));
KC_INV_X1 D8363 ( .Y(D8363_Y), .A(D8466_Y));
KC_INV_X1 D8362 ( .Y(D8362_Y), .A(D11887_Y));
KC_INV_X1 D8358 ( .Y(D8358_Y), .A(D8357_Y));
KC_INV_X1 D8296 ( .Y(D8296_Y), .A(D8342_Q));
KC_INV_X1 D8292 ( .Y(D8292_Y), .A(D1920_Y));
KC_INV_X1 D8290 ( .Y(D8290_Y), .A(D8048_Y));
KC_INV_X1 D8282 ( .Y(D8282_Y), .A(D8310_Y));
KC_INV_X1 D8261 ( .Y(D8261_Y), .A(D8262_Y));
KC_INV_X1 D8193 ( .Y(D8193_Y), .A(D740_Y));
KC_INV_X1 D8192 ( .Y(D8192_Y), .A(D8261_Y));
KC_INV_X1 D8191 ( .Y(D8191_Y), .A(D8244_Q));
KC_INV_X1 D8187 ( .Y(D8187_Y), .A(D5293_Y));
KC_INV_X1 D8186 ( .Y(D8186_Y), .A(D8240_Y));
KC_INV_X1 D8175 ( .Y(D8175_Y), .A(D8174_Y));
KC_INV_X1 D8172 ( .Y(D8172_Y), .A(D8207_Y));
KC_INV_X1 D8171 ( .Y(D8171_Y), .A(D5331_Y));
KC_INV_X1 D8170 ( .Y(D8170_Y), .A(D5268_Y));
KC_INV_X1 D8121 ( .Y(D8121_Y), .A(D8145_Q));
KC_INV_X1 D8120 ( .Y(D8120_Y), .A(D8242_Y));
KC_INV_X1 D8117 ( .Y(D8117_Y), .A(D8151_Q));
KC_INV_X1 D8110 ( .Y(D8110_Y), .A(D6633_Y));
KC_INV_X1 D8102 ( .Y(D8102_Y), .A(D674_Q));
KC_INV_X1 D8095 ( .Y(D8095_Y), .A(D8149_Q));
KC_INV_X1 D8088 ( .Y(D8088_Y), .A(D8156_Y));
KC_INV_X1 D8084 ( .Y(D8084_Y), .A(D9444_Y));
KC_INV_X1 D8083 ( .Y(D8083_Y), .A(D1839_Y));
KC_INV_X1 D8082 ( .Y(D8082_Y), .A(D3792_Y));
KC_INV_X1 D8079 ( .Y(D8079_Y), .A(D8254_Y));
KC_INV_X1 D8016 ( .Y(D8016_Y), .A(D1849_Y));
KC_INV_X1 D8015 ( .Y(D8015_Y), .A(D8073_Q));
KC_INV_X1 D8011 ( .Y(D8011_Y), .A(D7974_Y));
KC_INV_X1 D8009 ( .Y(D8009_Y), .A(D5172_Y));
KC_INV_X1 D8008 ( .Y(D8008_Y), .A(D6589_Y));
KC_INV_X1 D8007 ( .Y(D8007_Y), .A(D545_Y));
KC_INV_X1 D8006 ( .Y(D8006_Y), .A(D5154_Y));
KC_INV_X1 D8003 ( .Y(D8003_Y), .A(D9374_Y));
KC_INV_X1 D8002 ( .Y(D8002_Y), .A(D9368_Y));
KC_INV_X1 D8000 ( .Y(D8000_Y), .A(D5160_Y));
KC_INV_X1 D7999 ( .Y(D7999_Y), .A(D6585_Y));
KC_INV_X1 D7994 ( .Y(D7994_Y), .A(D5180_Y));
KC_INV_X1 D7988 ( .Y(D7988_Y), .A(D7937_Y));
KC_INV_X1 D7949 ( .Y(D7949_Y), .A(D152_Q));
KC_INV_X1 D7947 ( .Y(D7947_Y), .A(D7924_Y));
KC_INV_X1 D7941 ( .Y(D7941_Y), .A(D531_Q));
KC_INV_X1 D7940 ( .Y(D7940_Y), .A(D7986_Y));
KC_INV_X1 D7939 ( .Y(D7939_Y), .A(D7933_Y));
KC_INV_X1 D7927 ( .Y(D7927_Y), .A(D7922_Y));
KC_INV_X1 D7926 ( .Y(D7926_Y), .A(D533_Q));
KC_INV_X1 D7917 ( .Y(D7917_Y), .A(D532_Q));
KC_INV_X1 D7913 ( .Y(D7913_Y), .A(D6431_Y));
KC_INV_X1 D7910 ( .Y(D7910_Y), .A(D8375_Y));
KC_INV_X1 D7909 ( .Y(D7909_Y), .A(D8380_Y));
KC_INV_X1 D7908 ( .Y(D7908_Y), .A(D8398_Y));
KC_INV_X1 D7907 ( .Y(D7907_Y), .A(D8466_Y));
KC_INV_X1 D7905 ( .Y(D7905_Y), .A(D7827_Y));
KC_INV_X1 D7861 ( .Y(D7861_Y), .A(D7857_Y));
KC_INV_X1 D7860 ( .Y(D7860_Y), .A(D3379_Y));
KC_INV_X1 D7858 ( .Y(D7858_Y), .A(D7884_Q));
KC_INV_X1 D7856 ( .Y(D7856_Y), .A(D7846_Y));
KC_INV_X1 D7854 ( .Y(D7854_Y), .A(D7851_Y));
KC_INV_X1 D7850 ( .Y(D7850_Y), .A(D7886_Q));
KC_INV_X1 D7849 ( .Y(D7849_Y), .A(D7841_Y));
KC_INV_X1 D7843 ( .Y(D7843_Y), .A(D7828_Y));
KC_INV_X1 D7839 ( .Y(D7839_Y), .A(D7888_Q));
KC_INV_X1 D7835 ( .Y(D7835_Y), .A(D7955_Y));
KC_INV_X1 D7834 ( .Y(D7834_Y), .A(D7932_Y));
KC_INV_X1 D7833 ( .Y(D7833_Y), .A(D7862_Y));
KC_INV_X1 D7771 ( .Y(D7771_Y), .A(D4614_Y));
KC_INV_X1 D7767 ( .Y(D7767_Y), .A(D4770_Y));
KC_INV_X1 D7763 ( .Y(D7763_Y), .A(D7792_Y));
KC_INV_X1 D7759 ( .Y(D7759_Y), .A(D7823_Y));
KC_INV_X1 D7758 ( .Y(D7758_Y), .A(D7822_Y));
KC_INV_X1 D7752 ( .Y(D7752_Y), .A(D7753_Y));
KC_INV_X1 D7684 ( .Y(D7684_Y), .A(D6077_Y));
KC_INV_X1 D7680 ( .Y(D7680_Y), .A(D7737_Q));
KC_INV_X1 D7672 ( .Y(D7672_Y), .A(D7678_Y));
KC_INV_X1 D7639 ( .Y(D7639_Y), .A(D7727_Y));
KC_INV_X1 D7635 ( .Y(D7635_Y), .A(D7136_Y));
KC_INV_X1 D7633 ( .Y(D7633_Y), .A(D7667_Q));
KC_INV_X1 D7629 ( .Y(D7629_Y), .A(D7499_Y));
KC_INV_X1 D7621 ( .Y(D7621_Y), .A(D7620_Y));
KC_INV_X1 D7618 ( .Y(D7618_Y), .A(D6215_Y));
KC_INV_X1 D7567 ( .Y(D7567_Y), .A(D7519_Y));
KC_INV_X1 D7555 ( .Y(D7555_Y), .A(D7617_Y));
KC_INV_X1 D7545 ( .Y(D7545_Y), .A(D7564_Y));
KC_INV_X1 D7544 ( .Y(D7544_Y), .A(D1938_Y));
KC_INV_X1 D7506 ( .Y(D7506_Y), .A(D5641_Y));
KC_INV_X1 D7505 ( .Y(D7505_Y), .A(D7619_Y));
KC_INV_X1 D7501 ( .Y(D7501_Y), .A(D1711_Y));
KC_INV_X1 D7496 ( .Y(D7496_Y), .A(D7739_Y));
KC_INV_X1 D7490 ( .Y(D7490_Y), .A(D7573_Y));
KC_INV_X1 D7443 ( .Y(D7443_Y), .A(D7500_Y));
KC_INV_X1 D7442 ( .Y(D7442_Y), .A(D4116_Y));
KC_INV_X1 D7441 ( .Y(D7441_Y), .A(D7634_Y));
KC_INV_X1 D7436 ( .Y(D7436_Y), .A(D6021_Y));
KC_INV_X1 D7435 ( .Y(D7435_Y), .A(D179_Y));
KC_INV_X1 D7430 ( .Y(D7430_Y), .A(D7361_Y));
KC_INV_X1 D7429 ( .Y(D7429_Y), .A(D5984_Y));
KC_INV_X1 D7428 ( .Y(D7428_Y), .A(D7472_Y));
KC_INV_X1 D7421 ( .Y(D7421_Y), .A(D7476_Q));
KC_INV_X1 D7419 ( .Y(D7419_Y), .A(D5684_Y));
KC_INV_X1 D7411 ( .Y(D7411_Y), .A(D244_Y));
KC_INV_X1 D7360 ( .Y(D7360_Y), .A(D7201_Y));
KC_INV_X1 D7353 ( .Y(D7353_Y), .A(D7267_Y));
KC_INV_X1 D7344 ( .Y(D7344_Y), .A(D5705_Y));
KC_INV_X1 D7338 ( .Y(D7338_Y), .A(D1581_Y));
KC_INV_X1 D7337 ( .Y(D7337_Y), .A(D7352_Y));
KC_INV_X1 D7335 ( .Y(D7335_Y), .A(D7382_Y));
KC_INV_X1 D7334 ( .Y(D7334_Y), .A(D9478_Y));
KC_INV_X1 D7331 ( .Y(D7331_Y), .A(D7381_Y));
KC_INV_X1 D7329 ( .Y(D7329_Y), .A(D7210_Y));
KC_INV_X1 D7328 ( .Y(D7328_Y), .A(D7233_Y));
KC_INV_X1 D7327 ( .Y(D7327_Y), .A(D7232_Y));
KC_INV_X1 D7324 ( .Y(D7324_Y), .A(D7393_Y));
KC_INV_X1 D7323 ( .Y(D7323_Y), .A(D177_Y));
KC_INV_X1 D7318 ( .Y(D7318_Y), .A(D5864_Y));
KC_INV_X1 D7317 ( .Y(D7317_Y), .A(D7409_Q));
KC_INV_X1 D7308 ( .Y(D7308_Y), .A(D1740_Y));
KC_INV_X1 D7260 ( .Y(D7260_Y), .A(D6470_Y));
KC_INV_X1 D7250 ( .Y(D7250_Y), .A(D7241_Y));
KC_INV_X1 D7249 ( .Y(D7249_Y), .A(D5769_Y));
KC_INV_X1 D7248 ( .Y(D7248_Y), .A(D7152_Q));
KC_INV_X1 D7247 ( .Y(D7247_Y), .A(D7254_Y));
KC_INV_X1 D7239 ( .Y(D7239_Y), .A(D8742_Y));
KC_INV_X1 D7226 ( .Y(D7226_Y), .A(D7237_Y));
KC_INV_X1 D7225 ( .Y(D7225_Y), .A(D7266_Y));
KC_INV_X1 D7218 ( .Y(D7218_Y), .A(D7216_Y));
KC_INV_X1 D7217 ( .Y(D7217_Y), .A(D8747_Y));
KC_INV_X1 D7214 ( .Y(D7214_Y), .A(D220_Y));
KC_INV_X1 D7213 ( .Y(D7213_Y), .A(D7271_Y));
KC_INV_X1 D7212 ( .Y(D7212_Y), .A(D7234_Y));
KC_INV_X1 D7204 ( .Y(D7204_Y), .A(D7193_Y));
KC_INV_X1 D7203 ( .Y(D7203_Y), .A(D7304_Y));
KC_INV_X1 D7199 ( .Y(D7199_Y), .A(D7194_Y));
KC_INV_X1 D7188 ( .Y(D7188_Y), .A(D7268_Y));
KC_INV_X1 D7186 ( .Y(D7186_Y), .A(D7178_Y));
KC_INV_X1 D7185 ( .Y(D7185_Y), .A(D1956_Y));
KC_INV_X1 D7184 ( .Y(D7184_Y), .A(D5703_Y));
KC_INV_X1 D7183 ( .Y(D7183_Y), .A(D9476_Y));
KC_INV_X1 D7182 ( .Y(D7182_Y), .A(D7187_Y));
KC_INV_X1 D7172 ( .Y(D7172_Y), .A(D9475_Y));
KC_INV_X1 D7171 ( .Y(D7171_Y), .A(D7240_Y));
KC_INV_X1 D7170 ( .Y(D7170_Y), .A(D7303_Y));
KC_INV_X1 D7117 ( .Y(D7117_Y), .A(D7146_Q));
KC_INV_X1 D7112 ( .Y(D7112_Y), .A(D192_Q));
KC_INV_X1 D7109 ( .Y(D7109_Y), .A(D5672_Y));
KC_INV_X1 D7107 ( .Y(D7107_Y), .A(D6333_Y));
KC_INV_X1 D7106 ( .Y(D7106_Y), .A(D189_Y));
KC_INV_X1 D7101 ( .Y(D7101_Y), .A(D7141_Y));
KC_INV_X1 D7100 ( .Y(D7100_Y), .A(D7108_Y));
KC_INV_X1 D7099 ( .Y(D7099_Y), .A(D7137_Y));
KC_INV_X1 D7098 ( .Y(D7098_Y), .A(D7163_Y));
KC_INV_X1 D6992 ( .Y(D6992_Y), .A(D7026_Y));
KC_INV_X1 D6989 ( .Y(D6989_Y), .A(D5579_Y));
KC_INV_X1 D6986 ( .Y(D6986_Y), .A(D6985_Y));
KC_INV_X1 D6936 ( .Y(D6936_Y), .A(D6965_Q));
KC_INV_X1 D6931 ( .Y(D6931_Y), .A(D5502_Y));
KC_INV_X1 D6929 ( .Y(D6929_Y), .A(D5587_Y));
KC_INV_X1 D6927 ( .Y(D6927_Y), .A(D7074_Y));
KC_INV_X1 D6925 ( .Y(D6925_Y), .A(D6963_Q));
KC_INV_X1 D6924 ( .Y(D6924_Y), .A(D7021_Y));
KC_INV_X1 D6923 ( .Y(D6923_Y), .A(D6935_Y));
KC_INV_X1 D6922 ( .Y(D6922_Y), .A(D6962_Q));
KC_INV_X1 D6916 ( .Y(D6916_Y), .A(D5623_Y));
KC_INV_X1 D6877 ( .Y(D6877_Y), .A(D8393_Y));
KC_INV_X1 D6873 ( .Y(D6873_Y), .A(D976_Y));
KC_INV_X1 D6864 ( .Y(D6864_Y), .A(D6848_Y));
KC_INV_X1 D6855 ( .Y(D6855_Y), .A(D6854_Y));
KC_INV_X1 D6843 ( .Y(D6843_Y), .A(D970_Y));
KC_INV_X1 D6788 ( .Y(D6788_Y), .A(D5366_Y));
KC_INV_X1 D6787 ( .Y(D6787_Y), .A(D7928_Y));
KC_INV_X1 D6786 ( .Y(D6786_Y), .A(D8352_Y));
KC_INV_X1 D6783 ( .Y(D6783_Y), .A(D8330_Q));
KC_INV_X1 D6781 ( .Y(D6781_Y), .A(D1552_Y));
KC_INV_X1 D6777 ( .Y(D6777_Y), .A(D5387_Y));
KC_INV_X1 D6773 ( .Y(D6773_Y), .A(D8343_Q));
KC_INV_X1 D6772 ( .Y(D6772_Y), .A(D7974_Y));
KC_INV_X1 D6768 ( .Y(D6768_Y), .A(D3923_Y));
KC_INV_X1 D6767 ( .Y(D6767_Y), .A(D3903_Y));
KC_INV_X1 D6766 ( .Y(D6766_Y), .A(D8328_Q));
KC_INV_X1 D6765 ( .Y(D6765_Y), .A(D5429_Y));
KC_INV_X1 D6720 ( .Y(D6720_Y), .A(D6625_Y));
KC_INV_X1 D6711 ( .Y(D6711_Y), .A(D3829_Y));
KC_INV_X1 D6710 ( .Y(D6710_Y), .A(D6725_Y));
KC_INV_X1 D6702 ( .Y(D6702_Y), .A(D9365_Y));
KC_INV_X1 D6517 ( .Y(D6517_Y), .A(D7919_Y));
KC_INV_X1 D6512 ( .Y(D6512_Y), .A(D7920_Y));
KC_INV_X1 D6509 ( .Y(D6509_Y), .A(D8270_Y));
KC_INV_X1 D6508 ( .Y(D6508_Y), .A(D8277_Y));
KC_INV_X1 D6507 ( .Y(D6507_Y), .A(D8272_Y));
KC_INV_X1 D6506 ( .Y(D6506_Y), .A(D8409_Y));
KC_INV_X1 D6505 ( .Y(D6505_Y), .A(D8417_Y));
KC_INV_X1 D6504 ( .Y(D6504_Y), .A(D8273_Y));
KC_INV_X1 D6503 ( .Y(D6503_Y), .A(D8275_Y));
KC_INV_X1 D6502 ( .Y(D6502_Y), .A(D8391_Y));
KC_INV_X1 D6501 ( .Y(D6501_Y), .A(D8274_Y));
KC_INV_X1 D6499 ( .Y(D6499_Y), .A(D8269_Y));
KC_INV_X1 D6498 ( .Y(D6498_Y), .A(D1834_Y));
KC_INV_X1 D6449 ( .Y(D6449_Y), .A(D4865_Y));
KC_INV_X1 D6448 ( .Y(D6448_Y), .A(D6476_Q));
KC_INV_X1 D6438 ( .Y(D6438_Y), .A(D4885_Y));
KC_INV_X1 D6427 ( .Y(D6427_Y), .A(D7935_Y));
KC_INV_X1 D6423 ( .Y(D6423_Y), .A(D6472_Q));
KC_INV_X1 D6422 ( .Y(D6422_Y), .A(D6482_Y));
KC_INV_X1 D6418 ( .Y(D6418_Y), .A(D6516_Y));
KC_INV_X1 D6417 ( .Y(D6417_Y), .A(D6474_Q));
KC_INV_X1 D6416 ( .Y(D6416_Y), .A(D4995_Y));
KC_INV_X1 D6361 ( .Y(D6361_Y), .A(D1745_Y));
KC_INV_X1 D6298 ( .Y(D6298_Y), .A(D6348_Y));
KC_INV_X1 D6291 ( .Y(D6291_Y), .A(D1945_Y));
KC_INV_X1 D14498 ( .Y(D14498_Y), .A(D14139_Y));
KC_INV_X1 D13173 ( .Y(D13173_Y), .A(D12130_Y));
KC_INV_X1 D6231 ( .Y(D6231_Y), .A(D6229_Y));
KC_INV_X1 D6229 ( .Y(D6229_Y), .A(D6137_Y));
KC_INV_X1 D6228 ( .Y(D6228_Y), .A(D6337_Y));
KC_INV_X1 D6221 ( .Y(D6221_Y), .A(D6280_Y));
KC_INV_X1 D6218 ( .Y(D6218_Y), .A(D6238_Y));
KC_INV_X1 D6217 ( .Y(D6217_Y), .A(D6304_Y));
KC_INV_X1 D6212 ( .Y(D6212_Y), .A(D1419_Y));
KC_INV_X1 D6211 ( .Y(D6211_Y), .A(D430_Q));
KC_INV_X1 D6637 ( .Y(D6637_Y), .A(D9105_Y));
KC_INV_X1 D6149 ( .Y(D6149_Y), .A(D6196_Y));
KC_INV_X1 D6147 ( .Y(D6147_Y), .A(D6151_Y));
KC_INV_X1 D6146 ( .Y(D6146_Y), .A(D6202_Y));
KC_INV_X1 D6500 ( .Y(D6500_Y), .A(D6368_Y));
KC_INV_X1 D6098 ( .Y(D6098_Y), .A(D7512_Y));
KC_INV_X1 D6093 ( .Y(D6093_Y), .A(D1709_Y));
KC_INV_X1 D6091 ( .Y(D6091_Y), .A(D12305_Y));
KC_INV_X1 D6089 ( .Y(D6089_Y), .A(D335_Co));
KC_INV_X1 D6086 ( .Y(D6086_Y), .A(D6136_Y));
KC_INV_X1 D6039 ( .Y(D6039_Y), .A(D5685_Y));
KC_INV_X1 D6038 ( .Y(D6038_Y), .A(D6033_Y));
KC_INV_X1 D6037 ( .Y(D6037_Y), .A(D5792_Y));
KC_INV_X1 D6026 ( .Y(D6026_Y), .A(D4437_Y));
KC_INV_X1 D6025 ( .Y(D6025_Y), .A(D6113_Y));
KC_INV_X1 D6024 ( .Y(D6024_Y), .A(D5872_Y));
KC_INV_X1 D6023 ( .Y(D6023_Y), .A(D6020_Y));
KC_INV_X1 D6022 ( .Y(D6022_Y), .A(D7094_Y));
KC_INV_X1 D6013 ( .Y(D6013_Y), .A(D7480_Q));
KC_INV_X1 D6012 ( .Y(D6012_Y), .A(D6073_Q));
KC_INV_X1 D6002 ( .Y(D6002_Y), .A(D7177_Y));
KC_INV_X1 D6001 ( .Y(D6001_Y), .A(D266_Y));
KC_INV_X1 D5992 ( .Y(D5992_Y), .A(D5978_Y));
KC_INV_X1 D5990 ( .Y(D5990_Y), .A(D5971_Y));
KC_INV_X1 D5989 ( .Y(D5989_Y), .A(D6097_Y));
KC_INV_X1 D5988 ( .Y(D5988_Y), .A(D6044_Y));
KC_INV_X1 D5987 ( .Y(D5987_Y), .A(D5869_Y));
KC_INV_X1 D5986 ( .Y(D5986_Y), .A(D4415_Y));
KC_INV_X1 D5977 ( .Y(D5977_Y), .A(D6008_Y));
KC_INV_X1 D5976 ( .Y(D5976_Y), .A(D6099_Y));
KC_INV_X1 D5965 ( .Y(D5965_Y), .A(D6080_Y));
KC_INV_X1 D5964 ( .Y(D5964_Y), .A(D6046_Y));
KC_INV_X1 D5958 ( .Y(D5958_Y), .A(D275_Y));
KC_INV_X1 D5947 ( .Y(D5947_Y), .A(D4454_Y));
KC_INV_X1 D5890 ( .Y(D5890_Y), .A(D5771_Y));
KC_INV_X1 D5889 ( .Y(D5889_Y), .A(D5651_Y));
KC_INV_X1 D5877 ( .Y(D5877_Y), .A(D5876_Y));
KC_INV_X1 D5867 ( .Y(D5867_Y), .A(D5698_Y));
KC_INV_X1 D5866 ( .Y(D5866_Y), .A(D7164_Y));
KC_INV_X1 D5852 ( .Y(D5852_Y), .A(D5857_Y));
KC_INV_X1 D5851 ( .Y(D5851_Y), .A(D1735_Y));
KC_INV_X1 D5850 ( .Y(D5850_Y), .A(D5888_Y));
KC_INV_X1 D5841 ( .Y(D5841_Y), .A(D5973_Y));
KC_INV_X1 D5831 ( .Y(D5831_Y), .A(D7103_Y));
KC_INV_X1 D5830 ( .Y(D5830_Y), .A(D5677_Y));
KC_INV_X1 D5768 ( .Y(D5768_Y), .A(D5647_Y));
KC_INV_X1 D5763 ( .Y(D5763_Y), .A(D7263_Y));
KC_INV_X1 D5756 ( .Y(D5756_Y), .A(D7242_Y));
KC_INV_X1 D5755 ( .Y(D5755_Y), .A(D213_Y));
KC_INV_X1 D5754 ( .Y(D5754_Y), .A(D5745_Y));
KC_INV_X1 D5738 ( .Y(D5738_Y), .A(D5656_Y));
KC_INV_X1 D5730 ( .Y(D5730_Y), .A(D5715_Y));
KC_INV_X1 D5729 ( .Y(D5729_Y), .A(D5882_Y));
KC_INV_X1 D5723 ( .Y(D5723_Y), .A(D5714_Y));
KC_INV_X1 D5722 ( .Y(D5722_Y), .A(D5693_Q));
KC_INV_X1 D5670 ( .Y(D5670_Y), .A(D5690_Q));
KC_INV_X1 D5669 ( .Y(D5669_Y), .A(D5687_Q));
KC_INV_X1 D5665 ( .Y(D5665_Y), .A(D5691_Q));
KC_INV_X1 D5664 ( .Y(D5664_Y), .A(D5688_Q));
KC_INV_X1 D5655 ( .Y(D5655_Y), .A(D5666_Y));
KC_INV_X1 D5649 ( .Y(D5649_Y), .A(D4119_Q));
KC_INV_X1 D5648 ( .Y(D5648_Y), .A(D4129_Y));
KC_INV_X1 D5642 ( .Y(D5642_Y), .A(D6334_Y));
KC_INV_X1 D5510 ( .Y(D5510_Y), .A(D5520_Y));
KC_INV_X1 D5441 ( .Y(D5441_Y), .A(D5442_Y));
KC_INV_X1 D5432 ( .Y(D5432_Y), .A(D1628_Y));
KC_INV_X1 D5361 ( .Y(D5361_Y), .A(D5358_Y));
KC_INV_X1 D5360 ( .Y(D5360_Y), .A(D5369_Y));
KC_INV_X1 D5341 ( .Y(D5341_Y), .A(D5357_Y));
KC_INV_X1 D5260 ( .Y(D5260_Y), .A(D5267_Y));
KC_INV_X1 D5259 ( .Y(D5259_Y), .A(D6782_Y));
KC_INV_X1 D5098 ( .Y(D5098_Y), .A(D8399_Y));
KC_INV_X1 D5096 ( .Y(D5096_Y), .A(D5097_Y));
KC_INV_X1 D5095 ( .Y(D5095_Y), .A(D5017_Y));
KC_INV_X1 D5091 ( .Y(D5091_Y), .A(D4886_Y));
KC_INV_X1 D5044 ( .Y(D5044_Y), .A(D1567_Y));
KC_INV_X1 D5043 ( .Y(D5043_Y), .A(D1563_Y));
KC_INV_X1 D5033 ( .Y(D5033_Y), .A(D5019_Y));
KC_INV_X1 D5032 ( .Y(D5032_Y), .A(D5038_Y));
KC_INV_X1 D5023 ( .Y(D5023_Y), .A(D4877_Y));
KC_INV_X1 D5022 ( .Y(D5022_Y), .A(D4999_Y));
KC_INV_X1 D5012 ( .Y(D5012_Y), .A(D5020_Y));
KC_INV_X1 D5011 ( .Y(D5011_Y), .A(D3413_Y));
KC_INV_X1 D5004 ( .Y(D5004_Y), .A(D5009_Y));
KC_INV_X1 D5003 ( .Y(D5003_Y), .A(D4996_Y));
KC_INV_X1 D5002 ( .Y(D5002_Y), .A(D4881_Y));
KC_INV_X1 D4985 ( .Y(D4985_Y), .A(D1564_Y));
KC_INV_X1 D4977 ( .Y(D4977_Y), .A(D4976_Y));
KC_INV_X1 D4926 ( .Y(D4926_Y), .A(D3484_Q));
KC_INV_X1 D4925 ( .Y(D4925_Y), .A(D3388_Q));
KC_INV_X1 D4924 ( .Y(D4924_Y), .A(D454_Y));
KC_INV_X1 D4918 ( .Y(D4918_Y), .A(D4959_Y));
KC_INV_X1 D4917 ( .Y(D4917_Y), .A(D4965_Y));
KC_INV_X1 D4912 ( .Y(D4912_Y), .A(D4908_Y));
KC_INV_X1 D4911 ( .Y(D4911_Y), .A(D1537_Y));
KC_INV_X1 D4910 ( .Y(D4910_Y), .A(D4920_Y));
KC_INV_X1 D4903 ( .Y(D4903_Y), .A(D4914_Y));
KC_INV_X1 D4898 ( .Y(D4898_Y), .A(D3421_Y));
KC_INV_X1 D4897 ( .Y(D4897_Y), .A(D4916_Y));
KC_INV_X1 D4889 ( .Y(D4889_Y), .A(D3446_Y));
KC_INV_X1 D4883 ( .Y(D4883_Y), .A(D4922_Y));
KC_INV_X1 D4882 ( .Y(D4882_Y), .A(D4906_Y));
KC_INV_X1 D4869 ( .Y(D4869_Y), .A(D4907_Y));
KC_INV_X1 D4868 ( .Y(D4868_Y), .A(D4913_Y));
KC_INV_X1 D4867 ( .Y(D4867_Y), .A(D4900_Y));
KC_INV_X1 D4866 ( .Y(D4866_Y), .A(D3408_Y));
KC_INV_X1 D4857 ( .Y(D4857_Y), .A(D4858_Y));
KC_INV_X1 D4856 ( .Y(D4856_Y), .A(D4855_Y));
KC_INV_X1 D4853 ( .Y(D4853_Y), .A(D4854_Y));
KC_INV_X1 D4852 ( .Y(D4852_Y), .A(D4851_Y));
KC_INV_X1 D4849 ( .Y(D4849_Y), .A(D4850_Y));
KC_INV_X1 D4848 ( .Y(D4848_Y), .A(D4847_Y));
KC_INV_X1 D4846 ( .Y(D4846_Y), .A(D4845_Y));
KC_INV_X1 D4844 ( .Y(D4844_Y), .A(D4843_Y));
KC_INV_X1 D4779 ( .Y(D4779_Y), .A(D4785_Y));
KC_INV_X1 D4778 ( .Y(D4778_Y), .A(D4844_Y));
KC_INV_X1 D4771 ( .Y(D4771_Y), .A(D3383_Q));
KC_INV_X1 D4768 ( .Y(D4768_Y), .A(D4821_Q));
KC_INV_X1 D4767 ( .Y(D4767_Y), .A(D4822_Q));
KC_INV_X1 D4762 ( .Y(D4762_Y), .A(D4820_Q));
KC_INV_X1 D4756 ( .Y(D4756_Y), .A(D4823_Q));
KC_INV_X1 D4753 ( .Y(D4753_Y), .A(D9352_Y));
KC_INV_X1 D4745 ( .Y(D4745_Y), .A(D3380_Y));
KC_INV_X1 D4741 ( .Y(D4741_Y), .A(D371_Y));
KC_INV_X1 D4739 ( .Y(D4739_Y), .A(D92_Y));
KC_INV_X1 D4691 ( .Y(D4691_Y), .A(D4737_Y));
KC_INV_X1 D4683 ( .Y(D4683_Y), .A(D4724_Y));
KC_INV_X1 D4682 ( .Y(D4682_Y), .A(D4728_Q));
KC_INV_X1 D4681 ( .Y(D4681_Y), .A(D371_Y));
KC_INV_X1 D4667 ( .Y(D4667_Y), .A(D3319_Y));
KC_INV_X1 D4666 ( .Y(D4666_Y), .A(D4727_Q));
KC_INV_X1 D4664 ( .Y(D4664_Y), .A(D4702_Y));
KC_INV_X1 D4661 ( .Y(D4661_Y), .A(D4803_Y));
KC_INV_X1 D4660 ( .Y(D4660_Y), .A(D3298_Y));
KC_INV_X1 D4659 ( .Y(D4659_Y), .A(D3097_Y));
KC_INV_X1 D4606 ( .Y(D4606_Y), .A(D4568_Q));
KC_INV_X1 D4604 ( .Y(D4604_Y), .A(D4504_Y));
KC_INV_X1 D4603 ( .Y(D4603_Y), .A(D4612_Y));
KC_INV_X1 D4602 ( .Y(D4602_Y), .A(D7984_Y));
KC_INV_X1 D4598 ( .Y(D4598_Y), .A(D4601_Y));
KC_INV_X1 D4591 ( .Y(D4591_Y), .A(D3243_Y));
KC_INV_X1 D4589 ( .Y(D4589_Y), .A(D4637_Q));
KC_INV_X1 D4588 ( .Y(D4588_Y), .A(D4586_Y));
KC_INV_X1 D4587 ( .Y(D4587_Y), .A(D4639_Q));
KC_INV_X1 D4582 ( .Y(D4582_Y), .A(D4636_Q));
KC_INV_X1 D4581 ( .Y(D4581_Y), .A(D4638_Q));
KC_INV_X1 D4576 ( .Y(D4576_Y), .A(D3118_Y));
KC_INV_X1 D4575 ( .Y(D4575_Y), .A(D3112_Y));
KC_INV_X1 D4572 ( .Y(D4572_Y), .A(D3126_Y));
KC_INV_X1 D46 ( .Y(D46_Y), .A(D3037_Y));
KC_INV_X1 D4518 ( .Y(D4518_Y), .A(D4514_Y));
KC_INV_X1 D4517 ( .Y(D4517_Y), .A(D1593_Y));
KC_INV_X1 D4516 ( .Y(D4516_Y), .A(D4729_Q));
KC_INV_X1 D4515 ( .Y(D4515_Y), .A(D4495_Q));
KC_INV_X1 D4513 ( .Y(D4513_Y), .A(D6191_Y));
KC_INV_X1 D4506 ( .Y(D4506_Y), .A(D4587_Y));
KC_INV_X1 D4505 ( .Y(D4505_Y), .A(D328_Q));
KC_INV_X1 D4500 ( .Y(D4500_Y), .A(D47_Y));
KC_INV_X1 D4449 ( .Y(D4449_Y), .A(D4470_Y));
KC_INV_X1 D4441 ( .Y(D4441_Y), .A(D3038_Y));
KC_INV_X1 D4440 ( .Y(D4440_Y), .A(D8313_Q));
KC_INV_X1 D4439 ( .Y(D4439_Y), .A(D5969_Y));
KC_INV_X1 D4435 ( .Y(D4435_Y), .A(D302_Q));
KC_INV_X1 D4434 ( .Y(D4434_Y), .A(D2878_Y));
KC_INV_X1 D4428 ( .Y(D4428_Y), .A(D4488_Q));
KC_INV_X1 D4427 ( .Y(D4427_Y), .A(D4420_Y));
KC_INV_X1 D4421 ( .Y(D4421_Y), .A(D4149_Q));
KC_INV_X1 D4417 ( .Y(D4417_Y), .A(D165_Y));
KC_INV_X1 D4416 ( .Y(D4416_Y), .A(D239_Q));
KC_INV_X1 D4412 ( .Y(D4412_Y), .A(D228_Q));
KC_INV_X1 D4411 ( .Y(D4411_Y), .A(D4245_Y));
KC_INV_X1 D4405 ( .Y(D4405_Y), .A(D4438_Y));
KC_INV_X1 D4404 ( .Y(D4404_Y), .A(D1661_Y));
KC_INV_X1 D4401 ( .Y(D4401_Y), .A(D4400_Y));
KC_INV_X1 D4361 ( .Y(D4361_Y), .A(D4349_Y));
KC_INV_X1 D4350 ( .Y(D4350_Y), .A(D4301_Y));
KC_INV_X1 D4340 ( .Y(D4340_Y), .A(D5793_Y));
KC_INV_X1 D4339 ( .Y(D4339_Y), .A(D6007_Y));
KC_INV_X1 D4338 ( .Y(D4338_Y), .A(D249_Y));
KC_INV_X1 D4330 ( .Y(D4330_Y), .A(D4377_Y));
KC_INV_X1 D4328 ( .Y(D4328_Y), .A(D4368_Y));
KC_INV_X1 D4327 ( .Y(D4327_Y), .A(D4291_Y));
KC_INV_X1 D4320 ( .Y(D4320_Y), .A(D4422_Y));
KC_INV_X1 D4319 ( .Y(D4319_Y), .A(D262_Y));
KC_INV_X1 D4318 ( .Y(D4318_Y), .A(D4322_Y));
KC_INV_X1 D4310 ( .Y(D4310_Y), .A(D255_Y));
KC_INV_X1 D4306 ( .Y(D4306_Y), .A(D1629_Y));
KC_INV_X1 D4305 ( .Y(D4305_Y), .A(D4136_Q));
KC_INV_X1 D4304 ( .Y(D4304_Y), .A(D5863_Y));
KC_INV_X1 D4294 ( .Y(D4294_Y), .A(D4235_Q));
KC_INV_X1 D4293 ( .Y(D4293_Y), .A(D4296_Y));
KC_INV_X1 D4284 ( .Y(D4284_Y), .A(D5936_Y));
KC_INV_X1 D4270 ( .Y(D4270_Y), .A(D148_Q));
KC_INV_X1 D4267 ( .Y(D4267_Y), .A(D4268_Y));
KC_INV_X1 D4266 ( .Y(D4266_Y), .A(D4265_Y));
KC_INV_X1 D4261 ( .Y(D4261_Y), .A(D4260_Y));
KC_INV_X1 D4258 ( .Y(D4258_Y), .A(D4259_Y));
KC_INV_X1 D4256 ( .Y(D4256_Y), .A(D4255_Y));
KC_INV_X1 D4253 ( .Y(D4253_Y), .A(D4254_Y));
KC_INV_X1 D4252 ( .Y(D4252_Y), .A(D4251_Y));
KC_INV_X1 D4205 ( .Y(D4205_Y), .A(D3572_Y));
KC_INV_X1 D4188 ( .Y(D4188_Y), .A(D5847_Y));
KC_INV_X1 D4187 ( .Y(D4187_Y), .A(D232_Q));
KC_INV_X1 D4173 ( .Y(D4173_Y), .A(D4121_Q));
KC_INV_X1 D4172 ( .Y(D4172_Y), .A(D4347_Y));
KC_INV_X1 D4168 ( .Y(D4168_Y), .A(D229_Q));
KC_INV_X1 D4167 ( .Y(D4167_Y), .A(D4186_Y));
KC_INV_X1 D4159 ( .Y(D4159_Y), .A(D5825_Y));
KC_INV_X1 D4158 ( .Y(D4158_Y), .A(D5721_Y));
KC_INV_X1 D4151 ( .Y(D4151_Y), .A(D4152_Y));
KC_INV_X1 D4148 ( .Y(D4148_Y), .A(D4147_Y));
KC_INV_X1 D4146 ( .Y(D4146_Y), .A(D4208_Y));
KC_INV_X1 D4144 ( .Y(D4144_Y), .A(D4143_Y));
KC_INV_X1 D4141 ( .Y(D4141_Y), .A(D4142_Y));
KC_INV_X1 D4139 ( .Y(D4139_Y), .A(D4140_Y));
KC_INV_X1 D4097 ( .Y(D4097_Y), .A(D4120_Q));
KC_INV_X1 D4096 ( .Y(D4096_Y), .A(D4118_Q));
KC_INV_X1 D4094 ( .Y(D4094_Y), .A(D4122_Q));
KC_INV_X1 D4076 ( .Y(D4076_Y), .A(D7073_Y));
KC_INV_X1 D4032 ( .Y(D4032_Y), .A(D3881_Y));
KC_INV_X1 D3603 ( .Y(D3603_Y), .A(D4981_Y));
KC_INV_X1 D3602 ( .Y(D3602_Y), .A(D3500_Y));
KC_INV_X1 D3540 ( .Y(D3540_Y), .A(D3538_Y));
KC_INV_X1 D3539 ( .Y(D3539_Y), .A(D3409_Y));
KC_INV_X1 D3528 ( .Y(D3528_Y), .A(D3575_Q));
KC_INV_X1 D3522 ( .Y(D3522_Y), .A(D3533_Y));
KC_INV_X1 D3521 ( .Y(D3521_Y), .A(D4874_Y));
KC_INV_X1 D3517 ( .Y(D3517_Y), .A(D3545_Y));
KC_INV_X1 D3510 ( .Y(D3510_Y), .A(D3516_Y));
KC_INV_X1 D3509 ( .Y(D3509_Y), .A(D3516_Y));
KC_INV_X1 D3504 ( .Y(D3504_Y), .A(D3505_Y));
KC_INV_X1 D3503 ( .Y(D3503_Y), .A(D3542_Y));
KC_INV_X1 D3502 ( .Y(D3502_Y), .A(D3576_Q));
KC_INV_X1 D3497 ( .Y(D3497_Y), .A(D3470_Y));
KC_INV_X1 D3492 ( .Y(D3492_Y), .A(D4939_Y));
KC_INV_X1 D3448 ( .Y(D3448_Y), .A(D3479_Y));
KC_INV_X1 D3443 ( .Y(D3443_Y), .A(D3475_Y));
KC_INV_X1 D3432 ( .Y(D3432_Y), .A(D3415_Y));
KC_INV_X1 D3431 ( .Y(D3431_Y), .A(D3438_Y));
KC_INV_X1 D3430 ( .Y(D3430_Y), .A(D3428_Y));
KC_INV_X1 D3423 ( .Y(D3423_Y), .A(D4891_Y));
KC_INV_X1 D3416 ( .Y(D3416_Y), .A(D3477_Y));
KC_INV_X1 D3407 ( .Y(D3407_Y), .A(D3451_Y));
KC_INV_X1 D3406 ( .Y(D3406_Y), .A(D4923_Y));
KC_INV_X1 D3993 ( .Y(D3993_Y), .A(D3391_Y));
KC_INV_X1 D3398 ( .Y(D3398_Y), .A(D6344_Q));
KC_INV_X1 D3333 ( .Y(D3333_Y), .A(D3330_Y));
KC_INV_X1 D3332 ( .Y(D3332_Y), .A(D3205_Y));
KC_INV_X1 D3326 ( .Y(D3326_Y), .A(D3387_Q));
KC_INV_X1 D3318 ( .Y(D3318_Y), .A(D3369_Y));
KC_INV_X1 D3317 ( .Y(D3317_Y), .A(D3384_Q));
KC_INV_X1 D3315 ( .Y(D3315_Y), .A(D3389_Y));
KC_INV_X1 D3312 ( .Y(D3312_Y), .A(D3390_Y));
KC_INV_X1 D3309 ( .Y(D3309_Y), .A(D4749_Y));
KC_INV_X1 D3307 ( .Y(D3307_Y), .A(D6369_Y));
KC_INV_X1 D3306 ( .Y(D3306_Y), .A(D3374_Q));
KC_INV_X1 D3305 ( .Y(D3305_Y), .A(D3375_Q));
KC_INV_X1 D3303 ( .Y(D3303_Y), .A(D3373_Q));
KC_INV_X1 D3301 ( .Y(D3301_Y), .A(D12653_Y));
KC_INV_X1 D3299 ( .Y(D3299_Y), .A(D3322_Y));
KC_INV_X1 D3296 ( .Y(D3296_Y), .A(D3295_Y));
KC_INV_X1 D3234 ( .Y(D3234_Y), .A(D3349_Y));
KC_INV_X1 D3230 ( .Y(D3230_Y), .A(D3282_Q));
KC_INV_X1 D3226 ( .Y(D3226_Y), .A(D3296_Y));
KC_INV_X1 D3224 ( .Y(D3224_Y), .A(D3222_Y));
KC_INV_X1 D3223 ( .Y(D3223_Y), .A(D1469_Y));
KC_INV_X1 D3222 ( .Y(D3222_Y), .A(D3362_Y));
KC_INV_X1 D3219 ( .Y(D3219_Y), .A(D3261_Y));
KC_INV_X1 D3215 ( .Y(D3215_Y), .A(D3270_Y));
KC_INV_X1 D3209 ( .Y(D3209_Y), .A(D4815_Y));
KC_INV_X1 D3208 ( .Y(D3208_Y), .A(D3273_Y));
KC_INV_X1 D3207 ( .Y(D3207_Y), .A(D3291_Y));
KC_INV_X1 D3200 ( .Y(D3200_Y), .A(D4773_Y));
KC_INV_X1 D3198 ( .Y(D3198_Y), .A(D4592_Y));
KC_INV_X1 D3146 ( .Y(D3146_Y), .A(D3189_Q));
KC_INV_X1 D3145 ( .Y(D3145_Y), .A(D3139_Y));
KC_INV_X1 D3144 ( .Y(D3144_Y), .A(D3185_Q));
KC_INV_X1 D3143 ( .Y(D3143_Y), .A(D7641_Y));
KC_INV_X1 D3135 ( .Y(D3135_Y), .A(D3183_Y));
KC_INV_X1 D3134 ( .Y(D3134_Y), .A(D3186_Q));
KC_INV_X1 D3133 ( .Y(D3133_Y), .A(D3130_Y));
KC_INV_X1 D3120 ( .Y(D3120_Y), .A(D3137_Y));
KC_INV_X1 D3114 ( .Y(D3114_Y), .A(D3165_Y));
KC_INV_X1 D3113 ( .Y(D3113_Y), .A(D3116_Y));
KC_INV_X1 D3108 ( .Y(D3108_Y), .A(D1429_Y));
KC_INV_X1 D3094 ( .Y(D3094_Y), .A(D3195_Y));
KC_INV_X1 D45 ( .Y(D45_Y), .A(D3079_Q));
KC_INV_X1 D3031 ( .Y(D3031_Y), .A(D3073_Y));
KC_INV_X1 D3029 ( .Y(D3029_Y), .A(D3046_Y));
KC_INV_X1 D3028 ( .Y(D3028_Y), .A(D1516_Q));
KC_INV_X1 D3027 ( .Y(D3027_Y), .A(D3071_Y));
KC_INV_X1 D3023 ( .Y(D3023_Y), .A(D1515_Q));
KC_INV_X1 D3022 ( .Y(D3022_Y), .A(D3044_Y));
KC_INV_X1 D3021 ( .Y(D3021_Y), .A(D3062_Y));
KC_INV_X1 D3020 ( .Y(D3020_Y), .A(D3025_Y));
KC_INV_X1 D3016 ( .Y(D3016_Y), .A(D3084_Q));
KC_INV_X1 D3015 ( .Y(D3015_Y), .A(D3078_Q));
KC_INV_X1 D3011 ( .Y(D3011_Y), .A(D3036_Y));
KC_INV_X1 D2947 ( .Y(D2947_Y), .A(D3004_Q));
KC_INV_X1 D2946 ( .Y(D2946_Y), .A(D2857_Y));
KC_INV_X1 D2936 ( .Y(D2936_Y), .A(D301_Q));
KC_INV_X1 D2933 ( .Y(D2933_Y), .A(D2819_Y));
KC_INV_X1 D2916 ( .Y(D2916_Y), .A(D1438_Y));
KC_INV_X1 D2910 ( .Y(D2910_Y), .A(D5930_Y));
KC_INV_X1 D2908 ( .Y(D2908_Y), .A(D1435_Y));
KC_INV_X1 D2 ( .Y(D2_Y), .A(D1_Y));
KC_INV_X1 D2901 ( .Y(D2901_Y), .A(D2900_Y));
KC_INV_X1 D2852 ( .Y(D2852_Y), .A(D2766_Y));
KC_INV_X1 D2851 ( .Y(D2851_Y), .A(D2891_Q));
KC_INV_X1 D2848 ( .Y(D2848_Y), .A(D2816_Q));
KC_INV_X1 D2847 ( .Y(D2847_Y), .A(D2890_Q));
KC_INV_X1 D2844 ( .Y(D2844_Y), .A(D2792_Y));
KC_INV_X1 D2839 ( .Y(D2839_Y), .A(D2822_Y));
KC_INV_X1 D2835 ( .Y(D2835_Y), .A(D2886_Q));
KC_INV_X1 D2829 ( .Y(D2829_Y), .A(D2881_Y));
KC_INV_X1 D2826 ( .Y(D2826_Y), .A(D2887_Q));
KC_INV_X1 D2821 ( .Y(D2821_Y), .A(D2884_Q));
KC_INV_X1 D2820 ( .Y(D2820_Y), .A(D2836_Y));
KC_INV_X1 D2740 ( .Y(D2740_Y), .A(D2795_Q));
KC_INV_X1 D2815 ( .Y(D2815_Y), .A(D238_Y));
KC_INV_X1 D2810 ( .Y(D2810_Y), .A(D237_Y));
KC_INV_X1 D2770 ( .Y(D2770_Y), .A(D2799_Q));
KC_INV_X1 D2768 ( .Y(D2768_Y), .A(D2797_Q));
KC_INV_X1 D2767 ( .Y(D2767_Y), .A(D2783_Y));
KC_INV_X1 D2764 ( .Y(D2764_Y), .A(D2793_Y));
KC_INV_X1 D2758 ( .Y(D2758_Y), .A(D2813_Y));
KC_INV_X1 D2757 ( .Y(D2757_Y), .A(D2765_Y));
KC_INV_X1 D2750 ( .Y(D2750_Y), .A(D2845_Y));
KC_INV_X1 D2747 ( .Y(D2747_Y), .A(D2796_Q));
KC_INV_X1 D2741 ( .Y(D2741_Y), .A(D2798_Q));
KC_INV_X1 D2739 ( .Y(D2739_Y), .A(D2794_Q));
KC_INV_X1 D2663 ( .Y(D2663_Y), .A(D16189_Y));
KC_INV_X1 D2662 ( .Y(D2662_Y), .A(D16252_Y));
KC_INV_X1 D2654 ( .Y(D2654_Y), .A(D16047_Y));
KC_INV_X1 D2653 ( .Y(D2653_Y), .A(D16083_Y));
KC_INV_X1 D2652 ( .Y(D2652_Y), .A(D16085_Y));
KC_INV_X1 D2617 ( .Y(D2617_Y), .A(D16263_Y));
KC_INV_X1 D2616 ( .Y(D2616_Y), .A(D749_Y));
KC_INV_X1 D2610 ( .Y(D2610_Y), .A(D752_Y));
KC_INV_X1 D2609 ( .Y(D2609_Y), .A(D15469_Y));
KC_INV_X1 D2608 ( .Y(D2608_Y), .A(D14728_Y));
KC_INV_X1 D2603 ( .Y(D2603_Y), .A(D15668_Q));
KC_INV_X1 D2596 ( .Y(D2596_Y), .A(D15869_Q));
KC_INV_X1 D2591 ( .Y(D2591_Y), .A(D2587_Y));
KC_INV_X1 D2590 ( .Y(D2590_Y), .A(D15394_Y));
KC_INV_X1 D2548 ( .Y(D2548_Y), .A(D14499_Y));
KC_INV_X1 D2543 ( .Y(D2543_Y), .A(D14863_Y));
KC_INV_X1 D2539 ( .Y(D2539_Y), .A(D14875_Q));
KC_INV_X1 D2538 ( .Y(D2538_Y), .A(D953_Q));
KC_INV_X1 D2537 ( .Y(D2537_Y), .A(D14870_Q));
KC_INV_X1 D2529 ( .Y(D2529_Y), .A(D15996_Q));
KC_INV_X1 D2498 ( .Y(D2498_Y), .A(D13872_Q));
KC_INV_X1 D2428 ( .Y(D2428_Y), .A(D2426_Y));
KC_INV_X1 D2427 ( .Y(D2427_Y), .A(D13504_Y));
KC_INV_X1 D2414 ( .Y(D2414_Y), .A(D14301_Q));
KC_INV_X1 D2413 ( .Y(D2413_Y), .A(D14308_Q));
KC_INV_X1 D2375 ( .Y(D2375_Y), .A(D12928_Y));
KC_INV_X1 D2374 ( .Y(D2374_Y), .A(D12929_Y));
KC_INV_X1 D2373 ( .Y(D2373_Y), .A(D2371_Y));
KC_INV_X1 D2365 ( .Y(D2365_Y), .A(D13224_Y));
KC_INV_X1 D2328 ( .Y(D2328_Y), .A(D12780_Y));
KC_INV_X1 D2327 ( .Y(D2327_Y), .A(D12783_Y));
KC_INV_X1 D2312 ( .Y(D2312_Y), .A(D7670_Y));
KC_INV_X1 D2311 ( .Y(D2311_Y), .A(D12241_Y));
KC_INV_X1 D2230 ( .Y(D2230_Y), .A(D12071_Y));
KC_INV_X1 D2206 ( .Y(D2206_Y), .A(D10765_Y));
KC_INV_X1 D2205 ( .Y(D2205_Y), .A(D10692_Y));
KC_INV_X1 D2204 ( .Y(D2204_Y), .A(D10680_Y));
KC_INV_X1 D2202 ( .Y(D2202_Y), .A(D545_Y));
KC_INV_X1 D2123 ( .Y(D2123_Y), .A(D10629_Y));
KC_INV_X1 D2122 ( .Y(D2122_Y), .A(D5966_Y));
KC_INV_X1 D2119 ( .Y(D2119_Y), .A(D10191_Y));
KC_INV_X1 D2118 ( .Y(D2118_Y), .A(D10296_Q));
KC_INV_X1 D2110 ( .Y(D2110_Y), .A(D2109_Y));
KC_INV_X1 D2029 ( .Y(D2029_Y), .A(D2028_Y));
KC_INV_X1 D2028 ( .Y(D2028_Y), .A(D8854_Y));
KC_INV_X1 D2027 ( .Y(D2027_Y), .A(D9481_Y));
KC_INV_X1 D2016 ( .Y(D2016_Y), .A(D7522_Y));
KC_INV_X1 D2008 ( .Y(D2008_Y), .A(D9068_Y));
KC_INV_X1 D1998 ( .Y(D1998_Y), .A(D7896_Q));
KC_INV_X1 D1997 ( .Y(D1997_Y), .A(D154_Q));
KC_INV_X1 D1995 ( .Y(D1995_Y), .A(D9382_Y));
KC_INV_X1 D1994 ( .Y(D1994_Y), .A(D700_Q));
KC_INV_X1 D1991 ( .Y(D1991_Y), .A(D622_Y));
KC_INV_X1 D1990 ( .Y(D1990_Y), .A(D1983_Y));
KC_INV_X1 D1989 ( .Y(D1989_Y), .A(D1984_Y));
KC_INV_X1 D1988 ( .Y(D1988_Y), .A(D9582_Q));
KC_INV_X1 D1987 ( .Y(D1987_Y), .A(D1897_Y));
KC_INV_X1 D1978 ( .Y(D1978_Y), .A(D9870_Y));
KC_INV_X1 D1975 ( .Y(D1975_Y), .A(D2053_Y));
KC_INV_X1 D1971 ( .Y(D1971_Y), .A(D7227_Y));
KC_INV_X1 D1872 ( .Y(D1872_Y), .A(D726_Y));
KC_INV_X1 D1871 ( .Y(D1871_Y), .A(D6062_Y));
KC_INV_X1 D1859 ( .Y(D1859_Y), .A(D7923_Y));
KC_INV_X1 D1848 ( .Y(D1848_Y), .A(D1937_Y));
KC_INV_X1 D1845 ( .Y(D1845_Y), .A(D8018_Y));
KC_INV_X1 D1841 ( .Y(D1841_Y), .A(D8086_Y));
KC_INV_X1 D1840 ( .Y(D1840_Y), .A(D8246_Q));
KC_INV_X1 D1838 ( .Y(D1838_Y), .A(D8381_Y));
KC_INV_X1 D1832 ( .Y(D1832_Y), .A(D1212_Q));
KC_INV_X1 D1831 ( .Y(D1831_Y), .A(D1681_Y));
KC_INV_X1 D1828 ( .Y(D1828_Y), .A(D1935_Y));
KC_INV_X1 D1824 ( .Y(D1824_Y), .A(D1931_Q));
KC_INV_X1 D1821 ( .Y(D1821_Y), .A(D6426_Y));
KC_INV_X1 D1739 ( .Y(D1739_Y), .A(D5646_Y));
KC_INV_X1 D1738 ( .Y(D1738_Y), .A(D5737_Y));
KC_INV_X1 D1737 ( .Y(D1737_Y), .A(D1726_Y));
KC_INV_X1 D1736 ( .Y(D1736_Y), .A(D5644_Y));
KC_INV_X1 D1723 ( .Y(D1723_Y), .A(D7438_Y));
KC_INV_X1 D1713 ( .Y(D1713_Y), .A(D8838_Y));
KC_INV_X1 D1712 ( .Y(D1712_Y), .A(D6047_Y));
KC_INV_X1 D1706 ( .Y(D1706_Y), .A(D6239_Y));
KC_INV_X1 D1700 ( .Y(D1700_Y), .A(D6375_Q));
KC_INV_X1 D1699 ( .Y(D1699_Y), .A(D6376_Q));
KC_INV_X1 D1692 ( .Y(D1692_Y), .A(D8390_Y));
KC_INV_X1 D1592 ( .Y(D1592_Y), .A(D7243_Y));
KC_INV_X1 D1591 ( .Y(D1591_Y), .A(D5919_Y));
KC_INV_X1 D1586 ( .Y(D1586_Y), .A(D1627_Y));
KC_INV_X1 D1585 ( .Y(D1585_Y), .A(D4279_Y));
KC_INV_X1 D1584 ( .Y(D1584_Y), .A(D4448_Y));
KC_INV_X1 D1577 ( .Y(D1577_Y), .A(D4503_Y));
KC_INV_X1 D1576 ( .Y(D1576_Y), .A(D309_Y));
KC_INV_X1 D1574 ( .Y(D1574_Y), .A(D4640_Q));
KC_INV_X1 D1570 ( .Y(D1570_Y), .A(D3599_Y));
KC_INV_X1 D1565 ( .Y(D1565_Y), .A(D4902_Y));
KC_INV_X1 D1533 ( .Y(D1533_Y), .A(D3405_Y));
KC_INV_X1 D1442 ( .Y(D1442_Y), .A(D2737_Y));
KC_INV_X1 D1441 ( .Y(D1441_Y), .A(D2738_Y));
KC_INV_X1 D1432 ( .Y(D1432_Y), .A(D3190_Q));
KC_INV_X1 D1431 ( .Y(D1431_Y), .A(D3009_Y));
KC_INV_X1 D1428 ( .Y(D1428_Y), .A(D4687_Y));
KC_INV_X1 D1427 ( .Y(D1427_Y), .A(D1453_Y));
KC_INV_X1 D1426 ( .Y(D1426_Y), .A(D3184_Q));
KC_INV_X1 D1425 ( .Y(D1425_Y), .A(D3237_Y));
KC_INV_X1 D1424 ( .Y(D1424_Y), .A(D3128_Y));
KC_INV_X1 D1269 ( .Y(D1269_Y), .A(D15233_Q));
KC_INV_X1 D1268 ( .Y(D1268_Y), .A(D15232_Q));
KC_INV_X1 D1185 ( .Y(D1185_Y), .A(D13810_Q));
KC_INV_X1 D988 ( .Y(D988_Y), .A(D12950_Y));
KC_INV_X1 D966 ( .Y(D966_Y), .A(D13420_Y));
KC_INV_X1 D870 ( .Y(D870_Y), .A(D14305_Q));
KC_INV_X1 D866 ( .Y(D866_Y), .A(D13452_Y));
KC_INV_X1 D757 ( .Y(D757_Y), .A(D15425_Y));
KC_INV_X1 D754 ( .Y(D754_Y), .A(D13328_Y));
KC_INV_X1 D746 ( .Y(D746_Y), .A(D11218_Y));
KC_INV_X1 D744 ( .Y(D744_Y), .A(D11683_Y));
KC_INV_X1 D637 ( .Y(D637_Y), .A(D13995_Q));
KC_INV_X1 D569 ( .Y(D569_Y), .A(D2668_Y));
KC_INV_X1 D493 ( .Y(D493_Y), .A(D610_Y));
KC_INV_X1 D492 ( .Y(D492_Y), .A(D8057_Y));
KC_INV_X1 D432 ( .Y(D432_Y), .A(D3447_Y));
KC_INV_X1 D404 ( .Y(D404_Y), .A(D7749_Y));
KC_INV_X1 D402 ( .Y(D402_Y), .A(D3372_Q));
KC_INV_X1 D397 ( .Y(D397_Y), .A(D4763_Y));
KC_INV_X1 D370 ( .Y(D370_Y), .A(D7625_Y));
KC_INV_X1 D338 ( .Y(D338_Y), .A(D6248_Q));
KC_INV_X1 D336 ( .Y(D336_Y), .A(D3127_Y));
KC_INV_X1 D308 ( .Y(D308_Y), .A(D7447_Y));
KC_INV_X1 D287 ( .Y(D287_Y), .A(D5671_Y));
KC_INV_X1 D285 ( .Y(D285_Y), .A(D11_Y));
KC_INV_X1 D282 ( .Y(D282_Y), .A(D7479_Q));
KC_INV_X1 D247 ( .Y(D247_Y), .A(D214_Y));
KC_INV_X1 D243 ( .Y(D243_Y), .A(D7295_Y));
KC_INV_X1 D242 ( .Y(D242_Y), .A(D8900_Y));
KC_INV_X1 D240 ( .Y(D240_Y), .A(D1721_Y));
KC_INV_X1 D212 ( .Y(D212_Y), .A(D9980_Q));
KC_INV_X1 D209 ( .Y(D209_Y), .A(D9480_Y));
KC_INV_X1 D208 ( .Y(D208_Y), .A(D9982_Q));
KC_INV_X1 D203 ( .Y(D203_Y), .A(D7119_Y));
KC_INV_X1 D199 ( .Y(D199_Y), .A(D7211_Y));
KC_INV_X1 D175 ( .Y(D175_Y), .A(D8746_Y));
KC_INV_X1 D168 ( .Y(D168_Y), .A(D7918_Y));
KC_DFFSNHQ_X2 D16483 ( .Q(D16483_Q), .D(D16477_Y), .SN(D16377_Y),     .CK(D16455_Y));
KC_DFFSNHQ_X2 D16399 ( .Q(D16399_Q), .D(D16378_Y), .SN(D16376_Y),     .CK(D16455_Y));
KC_DFFSNHQ_X2 D16226 ( .Q(D16226_Q), .D(D2663_Y), .SN(D16383_Y),     .CK(D2568_Y));
KC_DFFSNHQ_X2 D13207 ( .Q(D13207_Q), .D(D2410_Y), .SN(D13192_Y),     .CK(D2460_Y));
KC_DFFSNHQ_X2 D12759 ( .Q(D12759_Q), .D(D12241_Y), .SN(D12258_Y),     .CK(D12740_Y));
KC_DFFSNHQ_X2 D12185 ( .Q(D12185_Q), .D(D12166_Y), .SN(D11636_SN),     .CK(D10707_Y));
KC_DFFSNHQ_X2 D12181 ( .Q(D12181_Q), .D(D11615_Y), .SN(D11636_SN),     .CK(D11635_Y));
KC_DFFSNHQ_X2 D12178 ( .Q(D12178_Q), .D(D12132_Y), .SN(D11636_SN),     .CK(D10707_Y));
KC_DFFSNHQ_X2 D11637 ( .Q(D11637_Q), .D(D509_Y), .SN(D11636_SN),     .CK(D540_Q));
KC_DFFSNHQ_X2 D11636 ( .Q(D11636_Q), .D(D11626_Y), .SN(D11636_SN),     .CK(D11133_Y));
KC_DFFSNHQ_X2 D10374 ( .Q(D10374_Q), .D(D951_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D10371 ( .Q(D10371_Q), .D(D945_Q), .SN(D9538_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D10370 ( .Q(D10370_Q), .D(D10366_Q), .SN(D9538_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D10366 ( .Q(D10366_Q), .D(D10368_Q), .SN(D9538_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D10316 ( .Q(D10316_Q), .D(D10309_Y), .SN(D10726_Y),     .CK(D11631_Y));
KC_DFFSNHQ_X2 D9639 ( .Q(D9639_Q), .D(D9630_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9638 ( .Q(D9638_Q), .D(D9628_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9637 ( .Q(D9637_Q), .D(D9638_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9635 ( .Q(D9635_Q), .D(D9634_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9634 ( .Q(D9634_Q), .D(D9625_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9630 ( .Q(D9630_Q), .D(D9637_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9629 ( .Q(D9629_Q), .D(D9623_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9628 ( .Q(D9628_Q), .D(D9620_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D9488 ( .Q(D9488_Q), .D(D714_Q), .SN(D9381_Y),     .CK(D10176_Y));
KC_DFFSNHQ_X2 D9385 ( .Q(D9385_Q), .D(D9384_Q), .SN(D9374_Y),     .CK(D9447_Y));
KC_DFFSNHQ_X2 D9384 ( .Q(D9384_Q), .D(D614_Q), .SN(D9374_Y),     .CK(D9447_Y));
KC_DFFSNHQ_X2 D9361 ( .Q(D9361_Q), .D(D9252_Y), .SN(D7893_Y),     .CK(D10107_QN));
KC_DFFSNHQ_X2 D9227 ( .Q(D9227_Q), .D(D9203_Y), .SN(D9214_Y),     .CK(D9212_QN));
KC_DFFSNHQ_X2 D9163 ( .Q(D9163_Q), .D(D9132_Y), .SN(D9214_Y),     .CK(D9143_QN));
KC_DFFSNHQ_X2 D9160 ( .Q(D9160_Q), .D(D9131_Y), .SN(D9214_Y),     .CK(D9143_QN));
KC_DFFSNHQ_X2 D9159 ( .Q(D9159_Q), .D(D9107_Y), .SN(D9214_Y),     .CK(D7530_QN));
KC_DFFSNHQ_X2 D7751 ( .Q(D7751_Q), .D(D7711_Y), .SN(D7788_Y),     .CK(D9211_QN));
KC_DFFSNHQ_X2 D7742 ( .Q(D7742_Q), .D(D7707_Y), .SN(D7788_Y),     .CK(D9211_QN));
KC_DFFSNHQ_X2 D7741 ( .Q(D7741_Q), .D(D1861_Y), .SN(D7893_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D7667 ( .Q(D7667_Q), .D(D376_Y), .SN(D9214_Y),     .CK(D9211_QN));
KC_DFFSNHQ_X2 D7615 ( .Q(D7615_Q), .D(D7543_Y), .SN(D7583_QN),     .CK(D7575_Y));
KC_DFFSNHQ_X2 D7614 ( .Q(D7614_Q), .D(D7615_Q), .SN(D7583_QN),     .CK(D7575_Y));
KC_DFFSNHQ_X2 D60 ( .Q(D60_Q), .D(D7535_Y), .SN(D9128_Y),     .CK(D9143_QN));
KC_DFFSNHQ_X2 D6491 ( .Q(D6491_Q), .D(D6439_Y), .SN(D6463_Y),     .CK(D4957_QN));
KC_DFFSNHQ_X2 D6486 ( .Q(D6486_Q), .D(D6489_Y), .SN(D6463_Y),     .CK(D6462_Y));
KC_DFFSNHQ_X2 D6359 ( .Q(D6359_Q), .D(D401_Y), .SN(D7893_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D6357 ( .Q(D6357_Q), .D(D6292_Y), .SN(D7795_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D6350 ( .Q(D6350_Q), .D(D6293_Y), .SN(D7893_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D6284 ( .Q(D6284_Q), .D(D6230_Y), .SN(D7660_Y),     .CK(D7575_Y));
KC_DFFSNHQ_X2 D4743 ( .Q(D4743_Q), .D(D3319_Y), .SN(D4827_Y),     .CK(D4799_Y));
KC_DFFSNHQ_X2 D4649 ( .Q(D4649_Q), .D(D6150_Y), .SN(D1934_Y),     .CK(D4527_Y));
KC_DFFSNHQ_X2 D4569 ( .Q(D4569_Q), .D(D4510_Y), .SN(D1652_Y),     .CK(D4527_Y));
KC_DFFSNHQ_X2 D4563 ( .Q(D4563_Q), .D(D4564_Y), .SN(D1652_Y),     .CK(D4462_Y));
KC_DFFSNHQ_X2 D4562 ( .Q(D4562_Q), .D(D4512_Y), .SN(D1652_Y),     .CK(D4527_Y));
KC_DFFSNHQ_X2 D4561 ( .Q(D4561_Q), .D(D4507_Y), .SN(D1652_Y),     .CK(D4527_Y));
KC_DFFSNHQ_X2 D4560 ( .Q(D4560_Q), .D(D4511_Y), .SN(D1652_Y),     .CK(D4527_Y));
KC_DFFSNHQ_X2 D2902 ( .Q(D2902_Q), .D(D2899_Y), .SN(D2882_Y),     .CK(D7712_Y));
KC_DFFSNHQ_X2 D2896 ( .Q(D2896_Q), .D(D13098_Y), .SN(D2882_Y),     .CK(D7712_Y));
KC_DFFSNHQ_X2 D2814 ( .Q(D2814_Q), .D(D2803_Y), .SN(D2882_Y),     .CK(D2864_Y));
KC_DFFSNHQ_X2 D2304 ( .Q(D2304_Q), .D(D12181_Q), .SN(D11636_SN),     .CK(D11635_Y));
KC_DFFSNHQ_X2 D2103 ( .Q(D2103_Q), .D(D9382_Y), .SN(D9375_Y),     .CK(D9346_Y));
KC_DFFSNHQ_X2 D1524 ( .Q(D1524_Q), .D(D1528_Y), .SN(D2882_Y),     .CK(D2864_Y));
KC_DFFSNHQ_X2 D947 ( .Q(D947_Q), .D(D9622_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D946 ( .Q(D946_Q), .D(D10374_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D945 ( .Q(D945_Q), .D(D10364_Q), .SN(D10357_Y),     .CK(D2176_Y));
KC_DFFSNHQ_X2 D837 ( .Q(D837_Q), .D(D9556_Y), .SN(D8229_Y),     .CK(D7962_Y));
KC_DFFSNHQ_X2 D835 ( .Q(D835_Q), .D(D10328_Y), .SN(D9538_Y),     .CK(D11631_Y));
KC_DFFSNHQ_X2 D714 ( .Q(D714_Q), .D(D9450_Y), .SN(D9381_Y),     .CK(D10176_Y));
KC_DFFSNHQ_X2 D614 ( .Q(D614_Q), .D(D538_Q), .SN(D9374_Y),     .CK(D9447_Y));
KC_DFFSNHQ_X2 D613 ( .Q(D613_Q), .D(D9385_Q), .SN(D9374_Y),     .CK(D9447_Y));
KC_DFFSNHQ_X2 D548 ( .Q(D548_Q), .D(D12150_Y), .SN(D11636_SN),     .CK(D10707_Y));
KC_DFFSNHQ_X2 D538 ( .Q(D538_Q), .D(D6483_Y), .SN(D9374_Y),     .CK(D9447_Y));
KC_DFFSNHQ_X2 D486 ( .Q(D486_Q), .D(D7860_Y), .SN(D7880_Y),     .CK(D4799_Y));
KC_DFFSNHQ_X2 D430 ( .Q(D430_Q), .D(D6299_Y), .SN(D7893_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D429 ( .Q(D429_Q), .D(D6214_Y), .SN(D7893_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D427 ( .Q(D427_Q), .D(D6213_Y), .SN(D7893_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D395 ( .Q(D395_Q), .D(D6222_Y), .SN(D1934_Y),     .CK(D6321_Y));
KC_DFFSNHQ_X2 D365 ( .Q(D365_Q), .D(D7583_QN), .SN(D10157_Y),     .CK(D7575_Y));
KC_DFFSNHQ_X2 D364 ( .Q(D364_Q), .D(D339_Y), .SN(D1934_Y),     .CK(D4527_Y));
KC_DFFSNHQ_X2 D363 ( .Q(D363_Q), .D(D348_Y), .SN(D9128_Y),     .CK(D9143_QN));
KC_DFFSNHQ_X2 D267 ( .Q(D267_Q), .D(D7380_Y), .SN(D8894_Y),     .CK(D9211_QN));
KC_DFFSNHQ_X2 D167 ( .Q(D167_Q), .D(D7772_Y), .SN(D7893_Y),     .CK(D6321_Y));
KC_MX2_X3 D16241 ( .Y(D16241_Y), .A(D16231_Y), .B(D16209_Y),     .S0(D16208_Y));
KC_MX2_X3 D16240 ( .Y(D16240_Y), .A(D16201_Y), .B(D14573_Y),     .S0(D15430_Y));
KC_MX2_X3 D16239 ( .Y(D16239_Y), .A(D16162_Y), .B(D16218_Y),     .S0(D16212_Y));
KC_MX2_X3 D16238 ( .Y(D16238_Y), .A(D16163_Y), .B(D15319_Y),     .S0(D15431_Y));
KC_MX2_X3 D16237 ( .Y(D16237_Y), .A(D16144_Y), .B(D16158_Y),     .S0(D16217_Y));
KC_MX2_X3 D16236 ( .Y(D16236_Y), .A(D16221_Y), .B(D16211_Y),     .S0(D16205_Y));
KC_MX2_X3 D16235 ( .Y(D16235_Y), .A(D16180_Y), .B(D16216_Y),     .S0(D16220_Y));
KC_MX2_X3 D16234 ( .Y(D16234_Y), .A(D16238_Y), .B(D15324_Y),     .S0(D14575_Y));
KC_MX2_X3 D16233 ( .Y(D16233_Y), .A(D16184_Y), .B(D15325_Y),     .S0(D15432_Y));
KC_MX2_X3 D16232 ( .Y(D16232_Y), .A(D16202_Y), .B(D15325_Y),     .S0(D15330_Y));
KC_MX2_X3 D16231 ( .Y(D16231_Y), .A(D16179_Y), .B(D15431_Y),     .S0(D15432_Y));
KC_MX2_X3 D16230 ( .Y(D16230_Y), .A(D16232_Y), .B(D15324_Y),     .S0(D16141_Y));
KC_MX2_X3 D16229 ( .Y(D16229_Y), .A(D16206_Y), .B(D16210_Y),     .S0(D16207_Y));
KC_MX2_X3 D16228 ( .Y(D16228_Y), .A(D16233_Y), .B(D16217_Y),     .S0(D16213_Y));
KC_MX2_X3 D16183 ( .Y(D16183_Y), .A(D16149_Y), .B(D16151_Y),     .S0(D16153_Y));
KC_MX2_X3 D16184 ( .Y(D16184_Y), .A(D16142_Y), .B(D15430_Y),     .S0(D15315_Y));
KC_MX2_X3 D16182 ( .Y(D16182_Y), .A(D16146_Y), .B(D16144_Y),     .S0(D15317_Y));
KC_MX2_X3 D16181 ( .Y(D16181_Y), .A(D16222_Y), .B(D16150_Y),     .S0(D16145_Y));
KC_MX2_X3 D16180 ( .Y(D16180_Y), .A(D16177_Y), .B(D14575_Y),     .S0(D15315_Y));
KC_MX2_X3 D16179 ( .Y(D16179_Y), .A(D14574_Y), .B(D15318_Y),     .S0(D15317_Y));
KC_MX2_X3 D16178 ( .Y(D16178_Y), .A(D16239_Y), .B(D16181_Y),     .S0(D16161_Y));
KC_MX2_X3 D16177 ( .Y(D16177_Y), .A(D719_Y), .B(D15330_Y),     .S0(D16222_Y));
KC_MX2_X3 D16176 ( .Y(D16176_Y), .A(D16178_Y), .B(D15319_Y),     .S0(D15434_Y));
KC_MX2_X3 D16098 ( .Y(D16098_Y), .A(D15254_Y), .B(D584_Y),     .S0(D13857_Y));
KC_MX2_X3 D16095 ( .Y(D16095_Y), .A(D16029_Y), .B(D16030_Y),     .S0(D16074_Y));
KC_MX2_X3 D16094 ( .Y(D16094_Y), .A(D16042_Y), .B(D15256_Y),     .S0(D15253_Y));
KC_MX2_X3 D16093 ( .Y(D16093_Y), .A(D15256_Y), .B(D16028_Y),     .S0(D16099_Y));
KC_MX2_X3 D16092 ( .Y(D16092_Y), .A(D16095_Y), .B(D15334_Y),     .S0(D16081_Y));
KC_MX2_X3 D16091 ( .Y(D16091_Y), .A(D16099_Y), .B(D16018_Y),     .S0(D16025_Y));
KC_MX2_X3 D16090 ( .Y(D16090_Y), .A(D16093_Y), .B(D16071_Y),     .S0(D15257_Y));
KC_MX2_X3 D16089 ( .Y(D16089_Y), .A(D16092_Y), .B(D15255_Y),     .S0(D13381_Y));
KC_MX2_X3 D16088 ( .Y(D16088_Y), .A(D2673_Y), .B(D15255_Y),     .S0(D15316_Y));
KC_MX2_X3 D16045 ( .Y(D16045_Y), .A(D16024_Y), .B(D16038_Y),     .S0(D16036_Y));
KC_MX2_X3 D16044 ( .Y(D16044_Y), .A(D15253_Y), .B(D16037_Y),     .S0(D16026_Y));
KC_MX2_X3 D16043 ( .Y(D16043_Y), .A(D542_Y), .B(D15254_Y),     .S0(D2667_Y));
KC_MX2_X3 D16042 ( .Y(D16042_Y), .A(D15261_Y), .B(D16025_Y),     .S0(D16041_Y));
KC_MX2_X3 D16041 ( .Y(D16041_Y), .A(D16022_Y), .B(D16035_Y),     .S0(D16029_Y));
KC_MX2_X3 D16040 ( .Y(D16040_Y), .A(D16045_Y), .B(D16034_Y),     .S0(D16044_Y));
KC_MX2_X3 D15600 ( .Y(D15600_Y), .A(D756_Y), .B(D15568_Y),     .S0(D9326_Y));
KC_MX2_X3 D15336 ( .Y(D15336_Y), .A(D617_Y), .B(D16075_Y),     .S0(D15328_Y));
KC_MX2_X3 D15335 ( .Y(D15335_Y), .A(D15263_Y), .B(D12637_Y),     .S0(D13857_Y));
KC_MX2_X3 D15334 ( .Y(D15334_Y), .A(D14373_Y), .B(D16020_Y),     .S0(D16046_Y));
KC_MX2_X3 D15266 ( .Y(D15266_Y), .A(D13170_Y), .B(D13411_Y),     .S0(D12238_Y));
KC_MX2_X3 D15264 ( .Y(D15264_Y), .A(D505_Y), .B(D16019_Y),     .S0(D16039_Y));
KC_MX2_X3 D15263 ( .Y(D15263_Y), .A(D15336_Y), .B(D13170_Y),     .S0(D13754_Y));
KC_MX2_X3 D15262 ( .Y(D15262_Y), .A(D15260_Y), .B(D12637_Y),     .S0(D12238_Y));
KC_MX2_X3 D15261 ( .Y(D15261_Y), .A(D15264_Y), .B(D15252_Y),     .S0(D110_Y));
KC_MX2_X3 D15260 ( .Y(D15260_Y), .A(D544_Y), .B(D16018_Y),     .S0(D2649_Y));
KC_MX2_X3 D14526 ( .Y(D14526_Y), .A(D14518_Q), .B(D14519_Q),     .S0(D490_Y));
KC_MX2_X3 D14525 ( .Y(D14525_Y), .A(D14518_Q), .B(D14519_Q),     .S0(D490_Y));
KC_MX2_X3 D13866 ( .Y(D13866_Y), .A(D14687_Q), .B(D465_Y),     .S0(D7823_Y));
KC_MX2_X3 D12180 ( .Y(D12180_Y), .A(D465_Y), .B(D9275_Q),     .S0(D7823_Y));
KC_MX2_X3 D10310 ( .Y(D10310_Y), .A(D10289_Y), .B(D10288_Y),     .S0(D10287_Y));
KC_MX2_X3 D10309 ( .Y(D10309_Y), .A(D540_Q), .B(D836_Q), .S0(D9566_Y));
KC_MX2_X3 D10233 ( .Y(D10233_Y), .A(D15440_Y), .B(D2119_Y),     .S0(D11146_Y));
KC_MX2_X3 D10232 ( .Y(D10232_Y), .A(D10233_Y), .B(D10178_Y),     .S0(D10201_Y));
KC_MX2_X3 D9633 ( .Y(D9633_Y), .A(D9631_Y), .B(D934_Q), .S0(D9623_Q));
KC_MX2_X3 D9632 ( .Y(D9632_Y), .A(D9625_Q), .B(D9637_Q), .S0(D946_Q));
KC_MX2_X3 D9631 ( .Y(D9631_Y), .A(D9632_Y), .B(D10370_Q),     .S0(D9638_Q));
KC_MX2_X3 D9484 ( .Y(D9484_Y), .A(D9459_Y), .B(D9460_Y),     .S0(D10215_Y));
KC_MX2_X3 D9297 ( .Y(D9297_Y), .A(D8893_Y), .B(D9258_Y), .S0(D9242_Y));
KC_MX2_X3 D9226 ( .Y(D9226_Y), .A(D9200_Y), .B(D7626_Y), .S0(D9241_Y));
KC_MX2_X3 D58 ( .Y(D58_Y), .A(D8990_Y), .B(D8976_Y), .S0(D2016_Y));
KC_MX2_X3 D8842 ( .Y(D8842_Y), .A(D8789_Y), .B(D8789_Y), .S0(D8773_Y));
KC_MX2_X3 D8733 ( .Y(D8733_Y), .A(D8674_Y), .B(D8728_Y), .S0(D8672_Y));
KC_MX2_X3 D8355 ( .Y(D8355_Y), .A(D8329_Q), .B(D8381_Y), .S0(D8176_Y));
KC_MX2_X3 D8354 ( .Y(D8354_Y), .A(D8283_Y), .B(D942_Y), .S0(D8310_Y));
KC_MX2_X3 D8259 ( .Y(D8259_Y), .A(D6719_Y), .B(D1894_Y), .S0(D6758_Q));
KC_MX2_X3 D8161 ( .Y(D8161_Y), .A(D1844_Y), .B(D8051_Q), .S0(D8437_Y));
KC_MX2_X3 D8160 ( .Y(D8160_Y), .A(D8081_Y), .B(D664_Q), .S0(D8438_Y));
KC_MX2_X3 D6352 ( .Y(D6352_Y), .A(D6349_Y), .B(D6327_Y), .S0(D6311_Y));
KC_MX2_X3 D6203 ( .Y(D6203_Y), .A(D6152_Y), .B(D6233_Y), .S0(D1703_Y));
KC_MX2_X3 D56 ( .Y(D56_Y), .A(D6160_Y), .B(D6205_Y), .S0(D6166_Y));
KC_MX2_X3 D48 ( .Y(D48_Y), .A(D6118_Y), .B(D6103_Y), .S0(D322_Y));
KC_MX2_X3 D34 ( .Y(D34_Y), .A(D7515_Y), .B(D6105_Y), .S0(D6089_Y));
KC_MX2_X3 D5417 ( .Y(D5417_Y), .A(D5342_Y), .B(D5412_Y), .S0(D5384_S));
KC_MX2_X3 D4840 ( .Y(D4840_Y), .A(D4698_Y), .B(D6329_Y), .S0(D4802_Y));
KC_MX2_X3 D4839 ( .Y(D4839_Y), .A(D9352_Y), .B(D4753_Y), .S0(D4752_Y));
KC_MX2_X3 D4735 ( .Y(D4735_Y), .A(D4714_Y), .B(D4714_Y), .S0(D4664_Y));
KC_MX2_X3 D55 ( .Y(D55_Y), .A(D377_Y), .B(D4468_Y), .S0(D395_Q));
KC_MX2_X3 D3588 ( .Y(D3588_Y), .A(D3555_Y), .B(D3587_Y), .S0(D5068_S));
KC_MX2_X3 D3587 ( .Y(D3587_Y), .A(D5083_Y), .B(D4981_Y), .S0(D3603_Y));
KC_MX2_X3 D3586 ( .Y(D3586_Y), .A(D1530_Y), .B(D1479_Y), .S0(D1505_Y));
KC_MX2_X3 D28 ( .Y(D28_Y), .A(D3070_Y), .B(D3070_Y), .S0(D2954_Y));
KC_MX2_X3 D5 ( .Y(D5_Y), .A(D2938_Y), .B(D2910_Y), .S0(D2983_Y));
KC_MX2_X3 D2649 ( .Y(D2649_Y), .A(D16021_Y), .B(D16031_Y),     .S0(D16029_Y));
KC_MX2_X3 D2261 ( .Y(D2261_Y), .A(D11191_Y), .B(D11328_Q),     .S0(D8434_Y));
KC_MX2_X3 D2108 ( .Y(D2108_Y), .A(D1895_Y), .B(D1895_Y), .S0(D9633_Y));
KC_MX2_X3 D2107 ( .Y(D2107_Y), .A(D2060_S), .B(D883_Y), .S0(D9598_Y));
KC_MX2_X3 D2106 ( .Y(D2106_Y), .A(D7896_Q), .B(D7819_Y), .S0(D154_Q));
KC_MX2_X3 D1968 ( .Y(D1968_Y), .A(D1960_Y), .B(D1827_Y), .S0(D1935_Y));
KC_MX2_X3 D1815 ( .Y(D1815_Y), .A(D1808_Y), .B(D1812_Y), .S0(D1968_Y));
KC_MX2_X3 D1531 ( .Y(D1531_Y), .A(D3407_Y), .B(D3454_Y), .S0(D3476_Y));
KC_MX2_X3 D1530 ( .Y(D1530_Y), .A(D3510_Y), .B(D3634_Y), .S0(D3602_Y));
KC_MX2_X3 D1245 ( .Y(D1245_Y), .A(D13724_Y), .B(D13736_Y),     .S0(D13768_Y));
KC_MX2_X3 D848 ( .Y(D848_Y), .A(D847_Y), .B(D12319_Y), .S0(D12320_Y));
KC_MX2_X3 D847 ( .Y(D847_Y), .A(D16070_Y), .B(D10291_Y),     .S0(D10751_Y));
KC_MX2_X3 D846 ( .Y(D846_Y), .A(D16240_Y), .B(D16160_Y),     .S0(D16182_Y));
KC_MX2_X3 D720 ( .Y(D720_Y), .A(D16176_Y), .B(D16148_Y),     .S0(D16159_Y));
KC_MX2_X3 D719 ( .Y(D719_Y), .A(D15318_Y), .B(D659_Y), .S0(D16158_Y));
KC_MX2_X3 D617 ( .Y(D617_Y), .A(D15251_Y), .B(D2670_Y), .S0(D16032_Y));
KC_MX2_X3 D546 ( .Y(D546_Y), .A(D16027_Y), .B(D16033_Y),     .S0(D16023_Y));
KC_MX2_X3 D544 ( .Y(D544_Y), .A(D546_Y), .B(D16028_Y), .S0(D1473_Y));
KC_MX2_X3 D542 ( .Y(D542_Y), .A(D16040_Y), .B(D13411_Y),     .S0(D13754_Y));
KC_MX2_X3 D541 ( .Y(D541_Y), .A(D14687_Q), .B(D465_Y), .S0(D7823_Y));
KC_MX2_X3 D428 ( .Y(D428_Y), .A(D10161_Y), .B(D6294_Y), .S0(D6356_Y));
KC_MX2_X3 D271 ( .Y(D271_Y), .A(D274_Co), .B(D4372_Y), .S0(D4369_Y));
KC_MX2_X3 D166 ( .Y(D166_Y), .A(D55_Y), .B(D5076_Y), .S0(D6494_Y));
KC_CELL_X2 D16405 ( .Y(D16405_Y), .A(D1405_Y), .B(D16455_Y),     .C(D16377_Y));
KC_CELL_X2 D16404 ( .Y(D16404_Y), .A(D16466_Y), .B(D16455_Y),     .C(D16377_Y));
KC_CELL_X2 D16402 ( .Y(D16402_Y), .A(D15699_Y), .B(D16455_Y),     .C(D16384_Y));
KC_CELL_X2 D16401 ( .Y(D16401_Y), .A(D15691_Y), .B(D16455_Y),     .C(D16384_Y));
KC_CELL_X2 D16371 ( .Y(D16371_Y), .A(D15608_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16370 ( .Y(D16370_Y), .A(D15688_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16368 ( .Y(D16368_Y), .A(D15586_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16367 ( .Y(D16367_Y), .A(D15649_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16366 ( .Y(D16366_Y), .A(D15678_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16344 ( .Y(D16344_Y), .A(D15700_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16343 ( .Y(D16343_Y), .A(D14904_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16339 ( .Y(D16339_Y), .A(D15774_Y), .B(D2586_Y),     .C(D16267_Y));
KC_CELL_X2 D16338 ( .Y(D16338_Y), .A(D15765_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D16335 ( .Y(D16335_Y), .A(D15587_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D16304 ( .Y(D16304_Y), .A(D14859_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D16303 ( .Y(D16303_Y), .A(D15684_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D16302 ( .Y(D16302_Y), .A(D15683_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D16301 ( .Y(D16301_Y), .A(D15694_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D16300 ( .Y(D16300_Y), .A(D15595_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D16244 ( .Y(D16244_Y), .A(D14786_Y), .B(D2568_Y),     .C(D15652_Y));
KC_CELL_X2 D16243 ( .Y(D16243_Y), .A(D15583_Y), .B(D2568_Y),     .C(D15652_Y));
KC_CELL_X2 D15957 ( .Y(D15957_Y), .A(D14760_Y), .B(D16455_Y),     .C(D16377_Y));
KC_CELL_X2 D15956 ( .Y(D15956_Y), .A(D15648_Y), .B(D16455_Y),     .C(D16376_Y));
KC_CELL_X2 D15710 ( .Y(D15710_Y), .A(D15597_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D14711 ( .Y(D14711_Y), .A(D14558_Y), .B(D14579_Y),     .C(D13265_Y));
KC_CELL_X2 D13287 ( .Y(D13287_Y), .A(D13913_Y), .B(D13251_Y),     .C(D13194_Y));
KC_CELL_X2 D13289 ( .Y(D13289_Y), .A(D13258_Y), .B(D13251_Y),     .C(D13194_Y));
KC_CELL_X2 D13288 ( .Y(D13288_Y), .A(D13894_Y), .B(D13251_Y),     .C(D13194_Y));
KC_CELL_X2 D13285 ( .Y(D13285_Y), .A(D13956_Y), .B(D13251_Y),     .C(D13194_Y));
KC_CELL_X2 D12863 ( .Y(D12863_Y), .A(D13183_Y), .B(D12740_Y),     .C(D12662_Y));
KC_CELL_X2 D12764 ( .Y(D12764_Y), .A(D13957_Y), .B(D13251_Y),     .C(D12679_Y));
KC_CELL_X2 D12763 ( .Y(D12763_Y), .A(D13915_Y), .B(D12740_Y),     .C(D12662_Y));
KC_CELL_X2 D12762 ( .Y(D12762_Y), .A(D13916_Y), .B(D12740_Y),     .C(D12662_Y));
KC_CELL_X2 D12761 ( .Y(D12761_Y), .A(D13917_Y), .B(D12740_Y),     .C(D12662_Y));
KC_CELL_X2 D12302 ( .Y(D12302_Y), .A(D12177_Q), .B(D10176_Y),     .C(D12177_RN));
KC_CELL_X2 D12301 ( .Y(D12301_Y), .A(D13230_Y), .B(D12740_Y),     .C(D12734_Y));
KC_CELL_X2 D12300 ( .Y(D12300_Y), .A(D2472_Y), .B(D12740_Y),     .C(D12662_Y));
KC_CELL_X2 D9340 ( .Y(D9340_Y), .A(D9252_Y), .B(D9212_QN),     .C(D7892_Y));
KC_CELL_X2 D9099 ( .Y(D9099_Y), .A(D9070_Y), .B(D7466_QN), .C(D324_Y));
KC_CELL_X2 D57 ( .Y(D57_Y), .A(D9073_Y), .B(D7468_QN), .C(D324_Y));
KC_CELL_X2 D51 ( .Y(D51_Y), .A(D311_Y), .B(D7468_QN), .C(D324_Y));
KC_CELL_X2 D41 ( .Y(D41_Y), .A(D8999_Y), .B(D7468_QN), .C(D324_Y));
KC_CELL_X2 D8903 ( .Y(D8903_Y), .A(D7387_Y), .B(D5931_QN),     .C(D8894_Y));
KC_CELL_X2 D8838 ( .Y(D8838_Y), .A(D7272_Y), .B(D5931_QN),     .C(D8818_Y));
KC_CELL_X2 D7823 ( .Y(D7823_Y), .A(D7773_Y), .B(D416_QN), .C(D7892_Y));
KC_CELL_X2 D7822 ( .Y(D7822_Y), .A(D7774_Y), .B(D416_QN), .C(D7788_Y));
KC_CELL_X2 D7819 ( .Y(D7819_Y), .A(D7777_Y), .B(D416_QN), .C(D7788_Y));
KC_CELL_X2 D7613 ( .Y(D7613_Y), .A(D9047_Y), .B(D7468_QN),     .C(D9128_Y));
KC_CELL_X2 D36 ( .Y(D36_Y), .A(D333_Y), .B(D7466_QN), .C(D4483_Y));
KC_CELL_X2 D8 ( .Y(D8_Y), .A(D7434_Y), .B(D4462_Y), .C(D9358_Y));
KC_CELL_X2 D4150 ( .Y(D4150_Y), .A(D4207_Y), .B(D5931_QN),     .C(D4461_Y));
KC_CELL_X2 D2687 ( .Y(D2687_Y), .A(D15680_Y), .B(D16349_Y),     .C(D16384_Y));
KC_CELL_X2 D2686 ( .Y(D2686_Y), .A(D15592_Y), .B(D16349_Y),     .C(D16267_Y));
KC_CELL_X2 D2685 ( .Y(D2685_Y), .A(D15548_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D2684 ( .Y(D2684_Y), .A(D14799_Y), .B(D2586_Y),     .C(D15652_Y));
KC_CELL_X2 D1249 ( .Y(D1249_Y), .A(D15944_Y), .B(D16455_Y),     .C(D16376_Y));
KC_CELL_X2 D1248 ( .Y(D1248_Y), .A(D2500_Y), .B(D16455_Y),     .C(D16377_Y));
KC_CELL_X2 D964 ( .Y(D964_Y), .A(D15701_Y), .B(D2586_Y), .C(D15652_Y));
KC_CELL_X2 D963 ( .Y(D963_Y), .A(D15575_Y), .B(D2586_Y), .C(D15652_Y));
KC_CELL_X2 D959 ( .Y(D959_Y), .A(D762_Y), .B(D2586_Y), .C(D15652_Y));
KC_CELL_X2 D727 ( .Y(D727_Y), .A(D10297_Q), .B(D9447_Y), .C(D10726_Y));
KC_CELL_X2 D726 ( .Y(D726_Y), .A(D12242_Y), .B(D12740_Y),     .C(D12734_Y));
KC_CELL_X2 D725 ( .Y(D725_Y), .A(D13919_Y), .B(D12740_Y),     .C(D12662_Y));
KC_CELL_X2 D724 ( .Y(D724_Y), .A(D13914_Y), .B(D12740_Y),     .C(D12662_Y));
KC_CELL_X2 D545 ( .Y(D545_Y), .A(D7983_Y), .B(D503_QN), .C(D9375_Y));
KC_CELL_X2 D490 ( .Y(D490_Y), .A(D9308_Y), .B(D416_QN), .C(D7892_Y));
KC_CELL_X2 D465 ( .Y(D465_Y), .A(D9248_Y), .B(D416_QN), .C(D7788_Y));
KC_CELL_X2 D7 ( .Y(D7_Y), .A(D8922_Y), .B(D296_QN), .C(D8894_Y));
KC_CELL_X2 D273 ( .Y(D273_Y), .A(D2020_Y), .B(D296_QN), .C(D8894_Y));
KC_CELL_X2 D272 ( .Y(D272_Y), .A(D2022_Y), .B(D296_QN), .C(D8894_Y));
KC_CELL_X2 D235 ( .Y(D235_Y), .A(D4209_Y), .B(D5931_QN), .C(D4461_Y));
KC_CELL_X2 D165 ( .Y(D165_Y), .A(D1811_Y), .B(D5931_QN), .C(D4461_Y));
KC_AOI32_X1 D16172 ( .B1(D16113_Y), .A2(D16137_Y), .Y(D16172_Y),     .A1(D2653_Y), .B0(D16083_Y), .A0(D2590_Y));
KC_AOI32_X1 D16087 ( .B1(D15311_Y), .A2(D16088_Y), .Y(D16087_Y),     .A1(D15311_Y), .B0(D16063_Y), .A0(D16090_Y));
KC_AOI32_X1 D15701 ( .B1(D15614_Y), .A2(D15495_Y), .Y(D15701_Y),     .A1(D15614_Y), .B0(D14830_Y), .A0(D15619_Y));
KC_AOI32_X1 D15700 ( .B1(D15613_Y), .A2(D14826_Y), .Y(D15700_Y),     .A1(D15613_Y), .B0(D14830_Y), .A0(D15467_Y));
KC_AOI32_X1 D15699 ( .B1(D15624_Y), .A2(D15618_Y), .Y(D15699_Y),     .A1(D15624_Y), .B0(D14830_Y), .A0(D15496_Y));
KC_AOI32_X1 D15597 ( .B1(D15515_Y), .A2(D15386_Y), .Y(D15597_Y),     .A1(D15515_Y), .B0(D15607_Y), .A0(D15524_Y));
KC_AOI32_X1 D15596 ( .B1(D14057_Y), .A2(D15509_Y), .Y(D15596_Y),     .A1(D14057_Y), .B0(D14745_Y), .A0(D14747_Y));
KC_AOI32_X1 D15595 ( .B1(D15541_Y), .A2(D15493_Y), .Y(D15595_Y),     .A1(D15541_Y), .B0(D15607_Y), .A0(D15388_Y));
KC_AOI32_X1 D15594 ( .B1(D15510_Y), .A2(D15507_Y), .Y(D15594_Y),     .A1(D15510_Y), .B0(D15607_Y), .A0(D15385_Y));
KC_AOI32_X1 D15593 ( .B1(D15486_Y), .A2(D15471_Y), .Y(D15593_Y),     .A1(D15486_Y), .B0(D15620_Y), .A0(D15465_Y));
KC_AOI32_X1 D15459 ( .B1(D15340_Y), .A2(D15530_Y), .Y(D15459_Y),     .A1(D15340_Y), .B0(D15512_Y), .A0(D15402_Y));
KC_AOI32_X1 D15458 ( .B1(D15370_Y), .A2(D15366_Y), .Y(D15458_Y),     .A1(D15370_Y), .B0(D15514_Y), .A0(D15374_Y));
KC_AOI32_X1 D15333 ( .B1(D15272_Y), .A2(D16052_Y), .Y(D15333_Y),     .A1(D15272_Y), .B0(D15338_Y), .A0(D15282_Y));
KC_AOI32_X1 D15332 ( .B1(D15293_Y), .A2(D2590_Y), .Y(D15332_Y),     .A1(D15291_Y), .B0(D2636_Y), .A0(D15301_Y));
KC_AOI32_X1 D15331 ( .B1(D15294_Y), .A2(D2590_Y), .Y(D15331_Y),     .A1(D569_Y), .B0(D2668_Y), .A0(D15303_Y));
KC_AOI32_X1 D14907 ( .B1(D888_Y), .A2(D2573_Q), .Y(D14907_Y),     .A1(D888_Y), .B0(D14081_Y), .A0(D815_Q));
KC_AOI32_X1 D14906 ( .B1(D14136_Y), .A2(D14790_Q), .Y(D14906_Y),     .A1(D14136_Y), .B0(D16765_Y), .A0(D820_Q));
KC_AOI32_X1 D14905 ( .B1(D15612_Y), .A2(D14827_Y), .Y(D14905_Y),     .A1(D15612_Y), .B0(D14830_Y), .A0(D752_Y));
KC_AOI32_X1 D14802 ( .B1(D14731_Y), .A2(D14025_Y), .Y(D14802_Y),     .A1(D14731_Y), .B0(D12856_Q), .A0(D2617_Y));
KC_AOI32_X1 D14704 ( .B1(D13947_Y), .A2(D13952_Y), .Y(D14704_Y),     .A1(D13947_Y), .B0(D14635_Y), .A0(D13997_Q));
KC_AOI32_X1 D14706 ( .B1(D14677_Y), .A2(D14708_Y), .Y(D14706_Y),     .A1(D14643_Y), .B0(D14688_Q), .A0(D14687_Q));
KC_AOI32_X1 D14705 ( .B1(D14637_Y), .A2(D14753_Y), .Y(D14705_Y),     .A1(D14532_Y), .B0(D14687_Q), .A0(D14557_Y));
KC_AOI32_X1 D14598 ( .B1(D14597_Y), .A2(D14576_Y), .Y(D14598_Y),     .A1(D14535_Y), .B0(D14519_Q), .A0(D14708_Y));
KC_AOI32_X1 D14597 ( .B1(D14805_Y), .A2(D14544_Y), .Y(D14597_Y),     .A1(D14805_Y), .B0(D14557_Y), .A0(D14518_Q));
KC_AOI32_X1 D14596 ( .B1(D14805_Y), .A2(D14542_Y), .Y(D14596_Y),     .A1(D14805_Y), .B0(D14557_Y), .A0(D14601_Q));
KC_AOI32_X1 D14595 ( .B1(D14596_Y), .A2(D14539_Y), .Y(D14595_Y),     .A1(D14552_Y), .B0(D608_Q), .A0(D14708_Y));
KC_AOI32_X1 D14594 ( .B1(D14567_Y), .A2(D14522_Y), .Y(D14594_Y),     .A1(D14548_Y), .B0(D14549_Y), .A0(D2564_Y));
KC_AOI32_X1 D14593 ( .B1(D14577_Y), .A2(D14542_Y), .Y(D14593_Y),     .A1(D14543_Y), .B0(D14601_Q), .A0(D14708_Y));
KC_AOI32_X1 D14524 ( .B1(D14688_Q), .A2(D14521_Y), .Y(D14524_Y),     .A1(D14643_Y), .B0(D2544_Y), .A0(D9457_Y));
KC_AOI32_X1 D14523 ( .B1(D14524_Y), .A2(D2547_Y), .Y(D14523_Y),     .A1(D14524_Y), .B0(D14532_Y), .A0(D14503_Y));
KC_AOI32_X1 D14522 ( .B1(D12173_Y), .A2(D14497_Y), .Y(D14522_Y),     .A1(D12173_Y), .B0(D14499_Y), .A0(D14518_Q));
KC_AOI32_X1 D14195 ( .B1(D14194_Y), .A2(D14168_Q), .Y(D14195_Y),     .A1(D14194_Y), .B0(D13985_Y), .A0(D14109_Q));
KC_AOI32_X1 D14111 ( .B1(D13323_Y), .A2(D14025_Y), .Y(D14111_Y),     .A1(D13328_Y), .B0(D754_Y), .A0(D14020_Y));
KC_AOI32_X1 D14000 ( .B1(D13928_Y), .A2(D14785_Y), .Y(D14000_Y),     .A1(D13928_Y), .B0(D14005_Y), .A0(D573_Y));
KC_AOI32_X1 D13769 ( .B1(D13752_Y), .A2(D13725_Y), .Y(D13769_Y),     .A1(D10266_Y), .B0(D13725_Y), .A0(D13730_Y));
KC_AOI32_X1 D13709 ( .B1(D2332_Y), .A2(D13672_Y), .Y(D13709_Y),     .A1(D2332_Y), .B0(D2411_Y), .A0(D13770_Q));
KC_AOI32_X1 D13708 ( .B1(D13706_Q), .A2(D12968_Y), .Y(D13708_Y),     .A1(D13706_Q), .B0(D13451_Y), .A0(D2435_Y));
KC_AOI32_X1 D13707 ( .B1(D1147_Q), .A2(D13029_Y), .Y(D13707_Y),     .A1(D1147_Q), .B0(D13558_Y), .A0(D13543_Y));
KC_AOI32_X1 D13633 ( .B1(D2391_Q), .A2(D13497_Y), .Y(D13633_Y),     .A1(D2391_Q), .B0(D13558_Y), .A0(D13543_Y));
KC_AOI32_X1 D13632 ( .B1(D14238_Q), .A2(D12972_Y), .Y(D13632_Y),     .A1(D14238_Q), .B0(D13457_Y), .A0(D13458_Y));
KC_AOI32_X1 D13631 ( .B1(D13703_Q), .A2(D2382_Y), .Y(D13631_Y),     .A1(D13703_Q), .B0(D2427_Y), .A0(D13466_Y));
KC_AOI32_X1 D13630 ( .B1(D13711_Q), .A2(D12969_Y), .Y(D13630_Y),     .A1(D13711_Q), .B0(D13459_Y), .A0(D2438_Y));
KC_AOI32_X1 D13629 ( .B1(D13590_Y), .A2(D13545_Y), .Y(D13629_Y),     .A1(D13590_Y), .B0(D13409_Y), .A0(D13588_Y));
KC_AOI32_X1 D13523 ( .B1(D13476_Y), .A2(D13323_Y), .Y(D13523_Y),     .A1(D13476_Y), .B0(D13477_Y), .A0(D7669_Y));
KC_AOI32_X1 D13522 ( .B1(D930_Q), .A2(D13497_Y), .Y(D13522_Y),     .A1(D930_Q), .B0(D13459_Y), .A0(D2438_Y));
KC_AOI32_X1 D13521 ( .B1(D13530_Q), .A2(D13442_Y), .Y(D13521_Y),     .A1(D13530_Q), .B0(D13454_Y), .A0(D13513_Y));
KC_AOI32_X1 D13520 ( .B1(D14165_Q), .A2(D13442_Y), .Y(D13520_Y),     .A1(D14165_Q), .B0(D13454_Y), .A0(D13461_Y));
KC_AOI32_X1 D13519 ( .B1(D928_Q), .A2(D13497_Y), .Y(D13519_Y),     .A1(D928_Q), .B0(D13457_Y), .A0(D13458_Y));
KC_AOI32_X1 D13518 ( .B1(D954_Q), .A2(D13497_Y), .Y(D13518_Y),     .A1(D954_Q), .B0(D13451_Y), .A0(D2435_Y));
KC_AOI32_X1 D13517 ( .B1(D12921_Q), .A2(D13442_Y), .Y(D13517_Y),     .A1(D12921_Q), .B0(D13454_Y), .A0(D886_Y));
KC_AOI32_X1 D13405 ( .B1(D13475_Y), .A2(D14017_Y), .Y(D13405_Y),     .A1(D13475_Y), .B0(D13314_Y), .A0(D14111_Y));
KC_AOI32_X1 D13278 ( .B1(D13241_Y), .A2(D13178_Y), .Y(D13278_Y),     .A1(D13231_Y), .B0(D13235_Y), .A0(D13938_Y));
KC_AOI32_X1 D13053 ( .B1(D13050_Q), .A2(D2381_Y), .Y(D13053_Y),     .A1(D13050_Q), .B0(D13571_Y), .A0(D13567_Y));
KC_AOI32_X1 D13008 ( .B1(D12996_Q), .A2(D13442_Y), .Y(D13008_Y),     .A1(D12996_Q), .B0(D13454_Y), .A0(D988_Y));
KC_AOI32_X1 D13007 ( .B1(D12994_Q), .A2(D13442_Y), .Y(D13007_Y),     .A1(D12994_Q), .B0(D13454_Y), .A0(D2373_Y));
KC_AOI32_X1 D13006 ( .B1(D12993_Q), .A2(D13442_Y), .Y(D13006_Y),     .A1(D12993_Q), .B0(D13454_Y), .A0(D12960_Y));
KC_AOI32_X1 D13005 ( .B1(D12997_Q), .A2(D13497_Y), .Y(D13005_Y),     .A1(D12997_Q), .B0(D13560_Y), .A0(D13548_Y));
KC_AOI32_X1 D13004 ( .B1(D12992_Q), .A2(D13578_Y), .Y(D13004_Y),     .A1(D12992_Q), .B0(D12946_Y), .A0(D12974_Y));
KC_AOI32_X1 D13003 ( .B1(D12973_Y), .A2(D13702_Y), .Y(D13003_Y),     .A1(D12973_Y), .B0(D13001_Y), .A0(D12970_Y));
KC_AOI32_X1 D13002 ( .B1(D12991_Q), .A2(D13497_Y), .Y(D13002_Y),     .A1(D12991_Q), .B0(D13571_Y), .A0(D13567_Y));
KC_AOI32_X1 D13001 ( .B1(D12952_Y), .A2(D12873_Y), .Y(D13001_Y),     .A1(D12952_Y), .B0(D12991_Q), .A0(D956_Q));
KC_AOI32_X1 D13000 ( .B1(D13051_Q), .A2(D12967_Y), .Y(D13000_Y),     .A1(D13051_Q), .B0(D13560_Y), .A0(D13548_Y));
KC_AOI32_X1 D12933 ( .B1(D12870_Y), .A2(D12875_Y), .Y(D12933_Y),     .A1(D12870_Y), .B0(D12919_Q), .A0(D146_Q));
KC_AOI32_X1 D12862 ( .B1(D13370_Y), .A2(D12858_Q), .Y(D12862_Y),     .A1(D12815_Y), .B0(D12748_Q), .A0(D12855_Q));
KC_AOI32_X1 D11670 ( .B1(D11657_Y), .A2(D10177_Y), .Y(D11670_Y),     .A1(D11657_Y), .B0(D11655_Y), .A0(D9371_Y));
KC_AOI32_X1 D10064 ( .B1(D347_Y), .A2(D10052_Y), .Y(D10064_Y),     .A1(D347_Y), .B0(D2122_Y), .A0(D10135_Y));
KC_AOI32_X1 D10063 ( .B1(D9078_Y), .A2(D10629_Y), .Y(D10063_Y),     .A1(D9078_Y), .B0(D10092_Y), .A0(D11623_Y));
KC_AOI32_X1 D9949 ( .B1(D183_Y), .A2(D9948_Y), .Y(D9949_Y),     .A1(D183_Y), .B0(D8769_Y), .A0(D9924_Y));
KC_AOI32_X1 D9948 ( .B1(D175_Y), .A2(D8669_Y), .Y(D9948_Y),     .A1(D175_Y), .B0(D9923_Y), .A0(D205_Y));
KC_AOI32_X1 D9589 ( .B1(D9522_Y), .A2(D9508_Y), .Y(D9589_Y),     .A1(D9578_Q), .B0(D9509_Y), .A0(D9511_Y));
KC_AOI32_X1 D9588 ( .B1(D9579_Q), .A2(D2039_Y), .Y(D9588_Y),     .A1(D9579_Q), .B0(D9532_Y), .A0(D9501_Y));
KC_AOI32_X1 D9587 ( .B1(D9577_Q), .A2(D2039_Y), .Y(D9587_Y),     .A1(D9577_Q), .B0(D9498_Y), .A0(D9597_Y));
KC_AOI32_X1 D9586 ( .B1(D9597_Y), .A2(D9502_Y), .Y(D9586_Y),     .A1(D9574_Q), .B0(D9543_Y), .A0(D9539_Y));
KC_AOI32_X1 D9339 ( .B1(D490_Y), .A2(D9266_Y), .Y(D9339_Y),     .A1(D490_Y), .B0(D1862_Y), .A0(D9237_Y));
KC_AOI32_X1 D9338 ( .B1(D7896_Q), .A2(D481_Y), .Y(D9338_Y),     .A1(D7896_Q), .B0(D1862_Y), .A0(D9237_Y));
KC_AOI32_X1 D9337 ( .B1(D13287_Y), .A2(D9306_Y), .Y(D9337_Y),     .A1(D13287_Y), .B0(D7779_Y), .A0(D9237_Y));
KC_AOI32_X1 D9292 ( .B1(D13289_Y), .A2(D9235_Y), .Y(D9292_Y),     .A1(D13289_Y), .B0(D7779_Y), .A0(D9237_Y));
KC_AOI32_X1 D9291 ( .B1(D724_Y), .A2(D9236_Y), .Y(D9291_Y),     .A1(D724_Y), .B0(D7779_Y), .A0(D9237_Y));
KC_AOI32_X1 D9290 ( .B1(D9275_Q), .A2(D9269_Y), .Y(D9290_Y),     .A1(D9275_Q), .B0(D1862_Y), .A0(D9237_Y));
KC_AOI32_X1 D9289 ( .B1(D154_Q), .A2(D7730_Y), .Y(D9289_Y),     .A1(D154_Q), .B0(D1862_Y), .A0(D9237_Y));
KC_AOI32_X1 D9288 ( .B1(D12764_Y), .A2(D1998_Y), .Y(D9288_Y),     .A1(D12764_Y), .B0(D7779_Y), .A0(D9237_Y));
KC_AOI32_X1 D9287 ( .B1(D723_Q), .A2(D1997_Y), .Y(D9287_Y),     .A1(D723_Q), .B0(D7779_Y), .A0(D9237_Y));
KC_AOI32_X1 D9162 ( .B1(D7497_Y), .A2(D6075_Y), .Y(D9162_Y),     .A1(D9166_Y), .B0(D9159_Q), .A0(D13171_Y));
KC_AOI32_X1 D9098 ( .B1(D8070_Y), .A2(D8985_Y), .Y(D9098_Y),     .A1(D8070_Y), .B0(D308_Y), .A0(D9059_Y));
KC_AOI32_X1 D9097 ( .B1(D8066_Y), .A2(D9109_Y), .Y(D9097_Y),     .A1(D8066_Y), .B0(D308_Y), .A0(D9059_Y));
KC_AOI32_X1 D9096 ( .B1(D615_Y), .A2(D9056_Y), .Y(D9096_Y),     .A1(D615_Y), .B0(D308_Y), .A0(D9059_Y));
KC_AOI32_X1 D9095 ( .B1(D8065_Y), .A2(D338_Y), .Y(D9095_Y),     .A1(D8065_Y), .B0(D308_Y), .A0(D9059_Y));
KC_AOI32_X1 D9094 ( .B1(D8067_Y), .A2(D9122_Y), .Y(D9094_Y),     .A1(D8067_Y), .B0(D308_Y), .A0(D9059_Y));
KC_AOI32_X1 D9026 ( .B1(D8979_Y), .A2(D1866_Y), .Y(D9026_Y),     .A1(D8979_Y), .B0(D7361_Y), .A0(D9002_Y));
KC_AOI32_X1 D8834 ( .B1(D8739_Y), .A2(D8823_Q), .Y(D8834_Y),     .A1(D8739_Y), .B0(D8737_Y), .A0(D227_Q));
KC_AOI32_X1 D8833 ( .B1(D8740_Y), .A2(D8784_Y), .Y(D8833_Y),     .A1(D8740_Y), .B0(D8746_Y), .A0(D233_Q));
KC_AOI32_X1 D8832 ( .B1(D9477_Y), .A2(D2027_Y), .Y(D8832_Y),     .A1(D9477_Y), .B0(D8743_Y), .A0(D8831_Y));
KC_AOI32_X1 D8831 ( .B1(D8877_Y), .A2(D7183_Y), .Y(D8831_Y),     .A1(D8877_Y), .B0(D9479_Y), .A0(D9480_Y));
KC_AOI32_X1 D8727 ( .B1(D8682_Y), .A2(D8771_Y), .Y(D8727_Y),     .A1(D8682_Y), .B0(D8820_Y), .A0(D8770_Y));
KC_AOI32_X1 D8726 ( .B1(D8724_Y), .A2(D8770_Y), .Y(D8726_Y),     .A1(D8771_Y), .B0(D8785_Y), .A0(D8724_Y));
KC_AOI32_X1 D8475 ( .B1(D8413_Y), .A2(D8419_Y), .Y(D8475_Y),     .A1(D8413_Y), .B0(D8400_Y), .A0(D8387_Y));
KC_AOI32_X1 D8474 ( .B1(D8368_Y), .A2(D8403_Y), .Y(D8474_Y),     .A1(D8388_Y), .B0(D8382_Y), .A0(D8387_Y));
KC_AOI32_X1 D7903 ( .B1(D7842_Y), .A2(D7859_Y), .Y(D7903_Y),     .A1(D7842_Y), .B0(D7857_Y), .A0(D7885_Q));
KC_AOI32_X1 D7902 ( .B1(D7842_Y), .A2(D7854_Y), .Y(D7902_Y),     .A1(D7842_Y), .B0(D7845_Y), .A0(D7889_Q));
KC_AOI32_X1 D7901 ( .B1(D7904_Y), .A2(D480_Q), .Y(D7901_Y),     .A1(D7904_Y), .B0(D7846_Y), .A0(D7886_Q));
KC_AOI32_X1 D7900 ( .B1(D7843_Y), .A2(D7849_Y), .Y(D7900_Y),     .A1(D7843_Y), .B0(D7869_Y), .A0(D7877_Y));
KC_AOI32_X1 D7899 ( .B1(D7842_Y), .A2(D7580_Y), .Y(D7899_Y),     .A1(D7842_Y), .B0(D7851_Y), .A0(D7887_Q));
KC_AOI32_X1 D7817 ( .B1(D13171_Y), .A2(D7783_Y), .Y(D7817_Y),     .A1(D13171_Y), .B0(D7779_Y), .A0(D9237_Y));
KC_AOI32_X1 D7816 ( .B1(D465_Y), .A2(D10162_Y), .Y(D7816_Y),     .A1(D465_Y), .B0(D1862_Y), .A0(D9237_Y));
KC_AOI32_X1 D7815 ( .B1(D7823_Y), .A2(D10161_Y), .Y(D7815_Y),     .A1(D7823_Y), .B0(D1862_Y), .A0(D9237_Y));
KC_AOI32_X1 D7744 ( .B1(D7751_Q), .A2(D1904_Y), .Y(D7744_Y),     .A1(D7751_Q), .B0(D7645_Y), .A0(D6075_Y));
KC_AOI32_X1 D7743 ( .B1(D7742_Q), .A2(D7629_Y), .Y(D7743_Y),     .A1(D7742_Q), .B0(D7645_Y), .A0(D6075_Y));
KC_AOI32_X1 D7538 ( .B1(D7496_Y), .A2(D9102_Y), .Y(D7538_Y),     .A1(D7739_Y), .B0(D7443_Y), .A0(D7501_Y));
KC_AOI32_X1 D7486 ( .B1(D6021_Y), .A2(D6035_Y), .Y(D7486_Y),     .A1(D7436_Y), .B0(D7435_Y), .A0(D7984_Y));
KC_AOI32_X1 D7485 ( .B1(D7430_Y), .A2(D5984_Y), .Y(D7485_Y),     .A1(D7430_Y), .B0(D177_Y), .A0(D6039_Y));
KC_AOI32_X1 D7484 ( .B1(D5991_Y), .A2(D382_Y), .Y(D7484_Y),     .A1(D5991_Y), .B0(D7421_Y), .A0(D7420_Y));
KC_AOI32_X1 D7399 ( .B1(D7337_Y), .A2(D7323_Y), .Y(D7399_Y),     .A1(D7337_Y), .B0(D7334_Y), .A0(D7204_Y));
KC_AOI32_X1 D7398 ( .B1(D1877_Y), .A2(D4116_Y), .Y(D7398_Y),     .A1(D1877_Y), .B0(D7210_Y), .A0(D7263_Y));
KC_AOI32_X1 D7301 ( .B1(D7183_Y), .A2(D7168_Y), .Y(D7301_Y),     .A1(D7183_Y), .B0(D7165_Y), .A0(D203_Y));
KC_AOI32_X1 D7300 ( .B1(D7184_Y), .A2(D8841_Y), .Y(D7300_Y),     .A1(D7184_Y), .B0(D1956_Y), .A0(D8822_Q));
KC_AOI32_X1 D7299 ( .B1(D7234_Y), .A2(D7218_Y), .Y(D7299_Y),     .A1(D7234_Y), .B0(D1885_Y), .A0(D7634_Y));
KC_AOI32_X1 D7159 ( .B1(D7244_Y), .A2(D5864_Y), .Y(D7159_Y),     .A1(D7244_Y), .B0(D7163_Y), .A0(D7106_Y));
KC_AOI32_X1 D6566 ( .B1(D7920_Y), .A2(D1694_Y), .Y(D6566_Y),     .A1(D7920_Y), .B0(D6514_Y), .A0(D1786_Q));
KC_AOI32_X1 D6403 ( .B1(D4949_Y), .A2(D6362_Y), .Y(D6403_Y),     .A1(D4949_Y), .B0(D4951_Y), .A0(D441_Y));
KC_AOI32_X1 D6404 ( .B1(D4949_Y), .A2(D1698_Y), .Y(D6404_Y),     .A1(D4949_Y), .B0(D4951_Y), .A0(D6363_Y));
KC_AOI32_X1 D6280 ( .B1(D6276_Y), .A2(D14498_Y), .Y(D6280_Y),     .A1(D6247_Y), .B0(D6254_Y), .A0(D6218_Y));
KC_AOI32_X1 D6201 ( .B1(D6180_Y), .A2(D6178_Y), .Y(D6201_Y),     .A1(D6163_Y), .B0(D6179_Y), .A0(D7784_Y));
KC_AOI32_X1 D6131 ( .B1(D6086_Y), .A2(D7531_Y), .Y(D6131_Y),     .A1(D16143_Y), .B0(D7531_Y), .A0(D6105_Y));
KC_AOI32_X1 D6130 ( .B1(D34_Y), .A2(D6088_Y), .Y(D6130_Y),     .A1(D1957_Y), .B0(D6129_Y), .A0(D6131_Y));
KC_AOI32_X1 D6083 ( .B1(D6039_Y), .A2(D5976_Y), .Y(D6083_Y),     .A1(D6039_Y), .B0(D6080_Y), .A0(D6008_Y));
KC_AOI32_X1 D6082 ( .B1(D6033_Y), .A2(D12305_Y), .Y(D6082_Y),     .A1(D6033_Y), .B0(D7687_Y), .A0(D266_Y));
KC_AOI32_X1 D6081 ( .B1(D6047_Y), .A2(D5977_Y), .Y(D6081_Y),     .A1(D6047_Y), .B0(D6094_Y), .A0(D5965_Y));
KC_AOI32_X1 D5943 ( .B1(D8865_Y), .A2(D5840_Y), .Y(D5943_Y),     .A1(D8865_Y), .B0(D7295_Y), .A0(D5846_Y));
KC_AOI32_X1 D5942 ( .B1(D5698_Y), .A2(D249_Y), .Y(D5942_Y),     .A1(D5698_Y), .B0(D5917_Y), .A0(D5889_Y));
KC_AOI32_X1 D5941 ( .B1(D7295_Y), .A2(D10050_Y), .Y(D5941_Y),     .A1(D7295_Y), .B0(D8865_Y), .A0(D5738_Y));
KC_AOI32_X1 D5940 ( .B1(D7310_Y), .A2(D1718_Y), .Y(D5940_Y),     .A1(D7310_Y), .B0(D5685_Y), .A0(D6027_Y));
KC_AOI32_X1 D5939 ( .B1(D177_Y), .A2(D5903_Y), .Y(D5939_Y),     .A1(D177_Y), .B0(D7232_Y), .A0(D6032_Y));
KC_AOI32_X1 D5821 ( .B1(D210_Y), .A2(D5729_Y), .Y(D5821_Y),     .A1(D210_Y), .B0(D5648_Y), .A0(D1734_Y));
KC_AOI32_X1 D5820 ( .B1(D20_Y), .A2(D1733_Y), .Y(D5820_Y), .A1(D235_Y),     .B0(D4186_Y), .A0(D5742_Y));
KC_AOI32_X1 D5819 ( .B1(D1730_Y), .A2(D5836_Y), .Y(D5819_Y),     .A1(D1730_Y), .B0(D5847_Y), .A0(D5782_Y));
KC_AOI32_X1 D5090 ( .B1(D4999_Y), .A2(D5041_Y), .Y(D5090_Y),     .A1(D4999_Y), .B0(D1567_Y), .A0(D4889_Y));
KC_AOI32_X1 D5089 ( .B1(D4877_Y), .A2(D4867_Y), .Y(D5089_Y),     .A1(D4877_Y), .B0(D5038_Y), .A0(D3446_Y));
KC_AOI32_X1 D5088 ( .B1(D4993_Y), .A2(D5001_Y), .Y(D5088_Y),     .A1(D3484_Q), .B0(D4926_Y), .A0(D5021_Y));
KC_AOI32_X1 D5087 ( .B1(D6427_Y), .A2(D4987_Y), .Y(D5087_Y),     .A1(D7935_Y), .B0(D6417_Y), .A0(D5089_Y));
KC_AOI32_X1 D5086 ( .B1(D5006_Y), .A2(D3556_Y), .Y(D5086_Y),     .A1(D5006_Y), .B0(D3484_Q), .A0(D3506_Y));
KC_AOI32_X1 D5085 ( .B1(D3400_Y), .A2(D1570_Y), .Y(D5085_Y),     .A1(D3400_Y), .B0(D5038_Y), .A0(D4874_Y));
KC_AOI32_X1 D4974 ( .B1(D4960_Y), .A2(D7966_Q), .Y(D4974_Y),     .A1(D4960_Y), .B0(D7968_Q), .A0(D3599_Y));
KC_AOI32_X1 D4973 ( .B1(D1537_Y), .A2(D3430_Y), .Y(D4973_Y),     .A1(D1537_Y), .B0(D4885_Y), .A0(D4875_Y));
KC_AOI32_X1 D4972 ( .B1(D3499_Y), .A2(D4926_Y), .Y(D4972_Y),     .A1(D3499_Y), .B0(D4877_Y), .A0(D4891_Y));
KC_AOI32_X1 D4971 ( .B1(D3499_Y), .A2(D1570_Y), .Y(D4971_Y),     .A1(D3416_Y), .B0(D3599_Y), .A0(D4952_Y));
KC_AOI32_X1 D4970 ( .B1(D4973_Y), .A2(D4933_Y), .Y(D4970_Y),     .A1(D4973_Y), .B0(D4926_Y), .A0(D4910_Y));
KC_AOI32_X1 D4969 ( .B1(D4884_Y), .A2(D4971_Y), .Y(D4969_Y),     .A1(D4884_Y), .B0(D4869_Y), .A0(D3371_Y));
KC_AOI32_X1 D4968 ( .B1(D3484_Q), .A2(D4916_Y), .Y(D4968_Y),     .A1(D3484_Q), .B0(D4967_Y), .A0(D4874_Y));
KC_AOI32_X1 D4967 ( .B1(D4913_Y), .A2(D4867_Y), .Y(D4967_Y),     .A1(D4913_Y), .B0(D4871_Y), .A0(D4906_Y));
KC_AOI32_X1 D4838 ( .B1(D1570_Y), .A2(D402_Y), .Y(D4838_Y),     .A1(D1570_Y), .B0(D3336_Y), .A0(D4906_Y));
KC_AOI32_X1 D4734 ( .B1(D4689_Y), .A2(D4706_Y), .Y(D4734_Y),     .A1(D4689_Y), .B0(D4691_Y), .A0(D1606_Y));
KC_AOI32_X1 D4733 ( .B1(D4638_Q), .A2(D4619_Y), .Y(D4733_Y),     .A1(D3243_Y), .B0(D4591_Y), .A0(D273_Y));
KC_AOI32_X1 D4732 ( .B1(D4577_Y), .A2(D4572_Y), .Y(D4732_Y),     .A1(D4577_Y), .B0(D3097_Y), .A0(D4709_Y));
KC_AOI32_X1 D4731 ( .B1(D4636_Q), .A2(D4619_Y), .Y(D4731_Y),     .A1(D3243_Y), .B0(D4591_Y), .A0(D7_Y));
KC_AOI32_X1 D4494 ( .B1(D4428_Y), .A2(D4516_Y), .Y(D4494_Y),     .A1(D4428_Y), .B0(D5677_Y), .A0(D4743_Q));
KC_AOI32_X1 D4493 ( .B1(D8313_Q), .A2(D4409_Y), .Y(D4493_Y),     .A1(D8313_Q), .B0(D4149_Q), .A0(D165_Y));
KC_AOI32_X1 D4398 ( .B1(D4185_Y), .A2(D5990_Y), .Y(D4398_Y),     .A1(D4185_Y), .B0(D1721_Y), .A0(D286_Y));
KC_AOI32_X1 D4397 ( .B1(D4327_Y), .A2(D4319_Y), .Y(D4397_Y),     .A1(D1629_Y), .B0(D148_Q), .A0(D4289_Y));
KC_AOI32_X1 D4249 ( .B1(D4118_Q), .A2(D4172_Y), .Y(D4249_Y),     .A1(D4118_Q), .B0(D4178_Y), .A0(D6039_Y));
KC_AOI32_X1 D4248 ( .B1(D4233_Y), .A2(D5753_Y), .Y(D4248_Y),     .A1(D4233_Y), .B0(D4211_Y), .A0(D8838_Y));
KC_AOI32_X1 D4247 ( .B1(D4233_Y), .A2(D5753_Y), .Y(D4247_Y),     .A1(D4233_Y), .B0(D4212_Y), .A0(D4150_Y));
KC_AOI32_X1 D4246 ( .B1(D4233_Y), .A2(D5753_Y), .Y(D4246_Y),     .A1(D4233_Y), .B0(D4217_Y), .A0(D239_Q));
KC_AOI32_X1 D4135 ( .B1(D5645_Y), .A2(D4197_Y), .Y(D4135_Y),     .A1(D5645_Y), .B0(D4092_Y), .A0(D4121_Q));
KC_AOI32_X1 D3585 ( .B1(D3594_Y), .A2(D3502_Y), .Y(D3585_Y),     .A1(D4925_Y), .B0(D3388_Q), .A0(D3498_Y));
KC_AOI32_X1 D3584 ( .B1(D3518_Y), .A2(D3575_Q), .Y(D3584_Y),     .A1(D3518_Y), .B0(D3539_Y), .A0(D68_Y));
KC_AOI32_X1 D3489 ( .B1(D4923_Y), .A2(D3363_Y), .Y(D3489_Y),     .A1(D4923_Y), .B0(D4938_Y), .A0(D3388_Q));
KC_AOI32_X1 D3488 ( .B1(D3388_Q), .A2(D3443_Y), .Y(D3488_Y),     .A1(D4925_Y), .B0(D3430_Y), .A0(D3400_Y));
KC_AOI32_X1 D3487 ( .B1(D4882_Y), .A2(D3304_Y), .Y(D3487_Y),     .A1(D4882_Y), .B0(D3405_Y), .A0(D4925_Y));
KC_AOI32_X1 D3486 ( .B1(D4960_Y), .A2(D4916_Y), .Y(D3486_Y),     .A1(D4960_Y), .B0(D3437_Y), .A0(D3446_Y));
KC_AOI32_X1 D3395 ( .B1(D1671_Y), .A2(D3339_Y), .Y(D3395_Y),     .A1(D1671_Y), .B0(D4749_Y), .A0(D3338_Y));
KC_AOI32_X1 D3394 ( .B1(D3309_Y), .A2(D3373_Q), .Y(D3394_Y),     .A1(D3309_Y), .B0(D3308_Y), .A0(D3375_Q));
KC_AOI32_X1 D3393 ( .B1(D3306_Y), .A2(D3540_Y), .Y(D3393_Y),     .A1(D3374_Q), .B0(D3442_Y), .A0(D3446_Y));
KC_AOI32_X1 D3294 ( .B1(D1456_Y), .A2(D3232_Y), .Y(D3294_Y),     .A1(D1456_Y), .B0(D1425_Y), .A0(D3283_Q));
KC_AOI32_X1 D3293 ( .B1(D9345_Y), .A2(D1428_Y), .Y(D3293_Y),     .A1(D9345_Y), .B0(D371_Y), .A0(D3252_Y));
KC_AOI32_X1 D3292 ( .B1(D3204_Y), .A2(D3207_Y), .Y(D3292_Y),     .A1(D3259_Y), .B0(D3290_Y), .A0(D3223_Y));
KC_AOI32_X1 D3092 ( .B1(D3032_Y), .A2(D31_Y), .Y(D3092_Y),     .A1(D4627_Y), .B0(D3063_Y), .A0(D2948_Y));
KC_AOI32_X1 D3007 ( .B1(D2931_Y), .A2(D2933_Y), .Y(D3007_Y),     .A1(D2931_Y), .B0(D4435_Y), .A0(D2981_Y));
KC_AOI32_X1 D3006 ( .B1(D2924_Y), .A2(D2933_Y), .Y(D3006_Y),     .A1(D2924_Y), .B0(D2947_Y), .A0(D2977_Y));
KC_AOI32_X1 D3005 ( .B1(D2923_Y), .A2(D2933_Y), .Y(D3005_Y),     .A1(D2923_Y), .B0(D2936_Y), .A0(D2980_Y));
KC_AOI32_X1 D2898 ( .B1(D2808_Y), .A2(D1437_Y), .Y(D2898_Y),     .A1(D2808_Y), .B0(D2738_Y), .A0(D2816_Q));
KC_AOI32_X1 D2897 ( .B1(D2849_Y), .A2(D2808_Y), .Y(D2897_Y),     .A1(D2849_Y), .B0(D2851_Y), .A0(D2738_Y));
KC_AOI32_X1 D2807 ( .B1(D2773_Y), .A2(D2793_Y), .Y(D2807_Y),     .A1(D2773_Y), .B0(D2747_Y), .A0(D2738_Y));
KC_AOI32_X1 D2806 ( .B1(D2751_Y), .A2(D2758_Y), .Y(D2806_Y),     .A1(D2751_Y), .B0(D2672_Y), .A0(D2765_Y));
KC_AOI32_X1 D2805 ( .B1(D2758_Y), .A2(D2833_Y), .Y(D2805_Y),     .A1(D2758_Y), .B0(D2765_Y), .A0(D2816_Q));
KC_AOI32_X1 D2683 ( .B1(D2650_Y), .A2(D2651_Y), .Y(D2683_Y),     .A1(D16049_Y), .B0(D16084_Y), .A0(D2590_Y));
KC_AOI32_X1 D2648 ( .B1(D15462_Y), .A2(D2607_Y), .Y(D2648_Y),     .A1(D15462_Y), .B0(D15622_Y), .A0(D2614_Y));
KC_AOI32_X1 D2473 ( .B1(D12919_Q), .A2(D13497_Y), .Y(D2473_Y),     .A1(D12919_Q), .B0(D2427_Y), .A0(D13466_Y));
KC_AOI32_X1 D2399 ( .B1(D1152_Q), .A2(D12949_Y), .Y(D2399_Y),     .A1(D1152_Q), .B0(D12946_Y), .A0(D13442_Y));
KC_AOI32_X1 D2398 ( .B1(D2375_Y), .A2(D12874_Y), .Y(D2398_Y),     .A1(D2375_Y), .B0(D12997_Q), .A0(D12926_Q));
KC_AOI32_X1 D2397 ( .B1(D2374_Y), .A2(D12874_Y), .Y(D2397_Y),     .A1(D2374_Y), .B0(D2391_Q), .A0(D929_Q));
KC_AOI32_X1 D2396 ( .B1(D12918_Q), .A2(D13442_Y), .Y(D2396_Y),     .A1(D12918_Q), .B0(D13454_Y), .A0(D12893_Y));
KC_AOI32_X1 D2358 ( .B1(D2311_Y), .A2(D2353_Y), .Y(D2358_Y),     .A1(D2311_Y), .B0(D552_Y), .A0(D2360_Y));
KC_AOI32_X1 D1963 ( .B1(D12301_Y), .A2(D5958_Y), .Y(D1963_Y),     .A1(D12301_Y), .B0(D5960_Y), .A0(D5872_Y));
KC_AOI32_X1 D1962 ( .B1(D7504_Y), .A2(D6040_Y), .Y(D1962_Y),     .A1(D7504_Y), .B0(D6091_Y), .A0(D73_Y));
KC_AOI32_X1 D1812 ( .B1(D1960_Y), .A2(D1935_Y), .Y(D1812_Y),     .A1(D1960_Y), .B0(D1826_Y), .A0(D1826_Y));
KC_AOI32_X1 D1811 ( .B1(D1729_Y), .A2(D252_Y), .Y(D1811_Y),     .A1(D1729_Y), .B0(D5847_Y), .A0(D5946_Y));
KC_AOI32_X1 D1810 ( .B1(D6427_Y), .A2(D4968_Y), .Y(D1810_Y),     .A1(D7935_Y), .B0(D6448_Y), .A0(D1559_Y));
KC_AOI32_X1 D1809 ( .B1(D6517_Y), .A2(D6419_Y), .Y(D1809_Y),     .A1(D6517_Y), .B0(D6512_Y), .A0(D1694_Y));
KC_AOI32_X1 D1670 ( .B1(D4233_Y), .A2(D4398_Y), .Y(D1670_Y),     .A1(D4233_Y), .B0(D4213_Y), .A0(D6039_Y));
KC_AOI32_X1 D1669 ( .B1(D4271_Y), .A2(D4470_Y), .Y(D1669_Y),     .A1(D4271_Y), .B0(D4280_Y), .A0(D1584_Y));
KC_AOI32_X1 D1668 ( .B1(D1572_Y), .A2(D4572_Y), .Y(D1668_Y),     .A1(D1572_Y), .B0(D3097_Y), .A0(D4681_Y));
KC_AOI32_X1 D1526 ( .B1(D1512_Y), .A2(D3447_Y), .Y(D1526_Y),     .A1(D3371_Y), .B0(D3498_Y), .A0(D3529_Y));
KC_AOI32_X1 D841 ( .B1(D13343_Y), .A2(D12793_Y), .Y(D841_Y),     .A1(D13349_Y), .B0(D819_Q), .A0(D12794_Y));
KC_AOI32_X1 D489 ( .B1(D6427_Y), .A2(D5018_Y), .Y(D489_Y),     .A1(D7935_Y), .B0(D6423_Y), .A0(D5088_Y));
KC_AOI32_X1 D234 ( .B1(D8751_Y), .A2(D8749_Y), .Y(D234_Y),     .A1(D8876_Y), .B0(D9476_Y), .A0(D9482_Y));
KC_AOI32_X1 D163 ( .B1(D9243_Y), .A2(D9168_Y), .Y(D163_Y),     .A1(D2120_Y), .B0(D10105_Y), .A0(D407_Y));
KC_AO22_X1 D12932 ( .Y(D12932_Y), .B1(D12915_Q), .B0(D12803_Y),     .A1(D2383_Y), .A0(D12917_Q));
KC_AO22_X1 D12931 ( .Y(D12931_Y), .B1(D12934_Q), .B0(D12803_Y),     .A1(D12907_Y), .A0(D12936_Q));
KC_AO22_X1 D12930 ( .Y(D12930_Y), .B1(D12914_Q), .B0(D12803_Y),     .A1(D12907_Y), .A0(D12923_Q));
KC_AO22_X1 D12929 ( .Y(D12929_Y), .B1(D12920_Q), .B0(D12803_Y),     .A1(D12902_Y), .A0(D12925_Q));
KC_AO22_X1 D12928 ( .Y(D12928_Y), .B1(D12922_Q), .B0(D12803_Y),     .A1(D12902_Y), .A0(D12924_Q));
KC_AO22_X1 D12861 ( .Y(D12861_Y), .B1(D12851_Q), .B0(D12803_Y),     .A1(D12830_Y), .A0(D12853_Q));
KC_AO22_X1 D12422 ( .Y(D12422_Y), .B1(D12794_Y), .B0(D12935_Q),     .A1(D12773_Y), .A0(D12415_Q));
KC_AO22_X1 D12421 ( .Y(D12421_Y), .B1(D12794_Y), .B0(D931_Q),     .A1(D12773_Y), .A0(D12414_Q));
KC_AO22_X1 D12420 ( .Y(D12420_Y), .B1(D12794_Y), .B0(D927_Q),     .A1(D12773_Y), .A0(D12418_Q));
KC_AO22_X1 D12305 ( .Y(D12305_Y), .B1(D12244_Y), .B0(D9345_Y),     .A1(D12660_Y), .A0(D14003_Y));
KC_AO22_X1 D12294 ( .Y(D12294_Y), .B1(D12295_Y), .B0(D9345_Y),     .A1(D12660_Y), .A0(D13950_Y));
KC_AO22_X1 D9286 ( .Y(D9286_Y), .B1(D9420_Y), .B0(D5966_Y),     .A1(D9240_Y), .A0(D9277_Q));
KC_AO22_X1 D9284 ( .Y(D9284_Y), .B1(D624_Y), .B0(D5966_Y),     .A1(D2002_Y), .A0(D9273_Q));
KC_AO22_X1 D9283 ( .Y(D9283_Y), .B1(D9490_Y), .B0(D5966_Y),     .A1(D9180_Y), .A0(D9274_Q));
KC_AO22_X1 D9225 ( .Y(D9225_Y), .B1(D9231_Q), .B0(D5966_Y),     .A1(D9167_Y), .A0(D9280_Q));
KC_AO22_X1 D9161 ( .Y(D9161_Y), .B1(D11116_Y), .B0(D5966_Y),     .A1(D9129_Y), .A0(D387_Q));
KC_AO22_X1 D9093 ( .Y(D9093_Y), .B1(D9276_Q), .B0(D9054_Y),     .A1(D8067_Y), .A0(D7473_Y));
KC_AO22_X1 D8725 ( .Y(D8725_Y), .B1(D7132_Y), .B0(D8690_Y),     .A1(D8688_Y), .A0(D7133_Y));
KC_AO22_X1 D8072 ( .Y(D8072_Y), .B1(D8275_Y), .B0(D8019_Y),     .A1(D6585_Y), .A0(D620_Y));
KC_AO22_X1 D8071 ( .Y(D8071_Y), .B1(D8390_Y), .B0(D8019_Y),     .A1(D5268_Y), .A0(D620_Y));
KC_AO22_X1 D8070 ( .Y(D8070_Y), .B1(D8274_Y), .B0(D8019_Y),     .A1(D5180_Y), .A0(D620_Y));
KC_AO22_X1 D8069 ( .Y(D8069_Y), .B1(D1834_Y), .B0(D8019_Y),     .A1(D5172_Y), .A0(D620_Y));
KC_AO22_X1 D8068 ( .Y(D8068_Y), .B1(D8409_Y), .B0(D8019_Y),     .A1(D740_Y), .A0(D620_Y));
KC_AO22_X1 D8067 ( .Y(D8067_Y), .B1(D8375_Y), .B0(D8019_Y),     .A1(D3776_Y), .A0(D620_Y));
KC_AO22_X1 D8066 ( .Y(D8066_Y), .B1(D8380_Y), .B0(D8019_Y),     .A1(D5293_Y), .A0(D620_Y));
KC_AO22_X1 D8065 ( .Y(D8065_Y), .B1(D8391_Y), .B0(D8019_Y),     .A1(D5288_Y), .A0(D620_Y));
KC_AO22_X1 D8064 ( .Y(D8064_Y), .B1(D8273_Y), .B0(D8019_Y),     .A1(D6580_Y), .A0(D620_Y));
KC_AO22_X1 D8061 ( .Y(D8061_Y), .B1(D8399_Y), .B0(D8019_Y),     .A1(D3792_Y), .A0(D620_Y));
KC_AO22_X1 D7482 ( .Y(D7482_Y), .B1(D4137_Q), .B0(D285_Y),     .A1(D7424_Y), .A0(D7426_Y));
KC_AO22_X1 D6277 ( .Y(D6277_Y), .B1(D6235_Y), .B0(D6212_Y),     .A1(D6269_Y), .A0(D6256_Y));
KC_AO22_X1 D6200 ( .Y(D6200_Y), .B1(D1795_Y), .B0(D6148_Y),     .A1(D6208_Co), .A0(D6199_Y));
KC_AO22_X1 D4837 ( .Y(D4837_Y), .B1(D4776_Y), .B0(D4821_Q),     .A1(D4777_Y), .A0(D4822_Q));
KC_AO22_X1 D4565 ( .Y(D4565_Y), .B1(D4466_Y), .B0(D4517_Y),     .A1(D4481_Y), .A0(D4517_Y));
KC_AO22_X1 D4134 ( .Y(D4134_Y), .B1(D4106_Y), .B0(D4145_Y),     .A1(D2716_Y), .A0(D4547_Y));
KC_AO22_X1 D3392 ( .Y(D3392_Y), .B1(D6369_Y), .B0(D3337_Y),     .A1(D3313_Y), .A0(D3307_Y));
KC_AO22_X1 D3289 ( .Y(D3289_Y), .B1(D3259_Y), .B0(D3259_Y),     .A1(D1469_Y), .A0(D3259_Y));
KC_AO22_X1 D2682 ( .Y(D2682_Y), .B1(D16085_Y), .B0(D16118_Y),     .A1(D2673_Y), .A0(D16178_Y));
KC_AO22_X1 D2472 ( .Y(D2472_Y), .B1(D2406_Y), .B0(D13257_Y),     .A1(D13400_Y), .A0(D999_Y));
KC_AO22_X1 D2395 ( .Y(D2395_Y), .B1(D12848_Q), .B0(D12803_Y),     .A1(D2383_Y), .A0(D12850_Q));
KC_AO22_X1 D2394 ( .Y(D2394_Y), .B1(D2392_Q), .B0(D12803_Y),     .A1(D12830_Y), .A0(D12852_Q));
KC_AO22_X1 D2173 ( .Y(D2173_Y), .B1(D12287_Y), .B0(D5966_Y),     .A1(D2044_Y), .A0(D353_Q));
KC_AO22_X1 D1808 ( .Y(D1808_Y), .B1(D1935_Y), .B0(D1826_Y),     .A1(D1827_Y), .A0(D1827_Y));
KC_AO22_X1 D950 ( .Y(D950_Y), .B1(D12794_Y), .B0(D12916_Q),     .A1(D12773_Y), .A0(D12417_Q));
KC_AO22_X1 D949 ( .Y(D949_Y), .B1(D12794_Y), .B0(D932_Q),     .A1(D12773_Y), .A0(D12419_Q));
KC_AO22_X1 D715 ( .Y(D715_Y), .B1(D8836_Q), .B0(D8120_Y), .A1(D8139_Y),     .A0(D703_Q));
KC_AO22_X1 D615 ( .Y(D615_Y), .B1(D8269_Y), .B0(D8019_Y), .A1(D6589_Y),     .A0(D620_Y));
KC_AO22_X1 D162 ( .Y(D162_Y), .B1(D12794_Y), .B0(D842_Q),     .A1(D12773_Y), .A0(D12340_Q));
KC_AO21_X1 D15592 ( .B(D15549_Y), .A1(D15599_Y), .Y(D15592_Y),     .A0(D14750_Y));
KC_AO21_X1 D14904 ( .B(D14860_Y), .A1(D15598_Y), .Y(D14904_Y),     .A0(D14829_Y));
KC_AO21_X1 D161 ( .B(D4489_Q), .A1(D1610_Y), .Y(D161_Y), .A0(D6239_Y));
KC_BUF_X13 D16731 ( .Y(D16731_Y), .A(D16728_Y));
KC_BUF_X13 D16711 ( .Y(D16711_Y), .A(D16703_Y));
KC_BUF_X13 D16636 ( .Y(D16636_Y), .A(D16630_Y));
KC_BUF_X13 D16618 ( .Y(D16618_Y), .A(D16620_Y));
KC_BUF_X13 D16334 ( .Y(D16334_Y), .A(D16133_Y));
KC_BUF_X13 D16333 ( .Y(D16333_Y), .A(D16323_Y));
KC_BUF_X13 D15155 ( .Y(D15155_Y), .A(D15136_Y));
KC_BUF_X13 D15154 ( .Y(D15154_Y), .A(D15137_Y));
KC_BUF_X13 D13838 ( .Y(D13838_Y), .A(D13831_Y));
KC_BUF_X13 D13623 ( .Y(D13623_Y), .A(D13617_Y));
KC_BUF_X13 D12513 ( .Y(D12513_Y), .A(D2402_Y));
KC_BUF_X13 D12292 ( .Y(D12292_Y), .A(D12282_Y));
KC_BUF_X13 D11607 ( .Y(D11607_Y), .A(D11599_Y));
KC_BUF_X13 D10827 ( .Y(D10827_Y), .A(D10816_Y));
KC_BUF_X13 D9920 ( .Y(D9920_Y), .A(D9916_Y));
KC_BUF_X13 D9919 ( .Y(D9919_Y), .A(D9913_Y));
KC_BUF_X13 D9583 ( .Y(D9583_Y), .A(D9625_Q));
KC_BUF_X13 D6564 ( .Y(D6564_Y), .A(D6560_Y));
KC_BUF_X13 D6126 ( .Y(D6126_Y), .A(D27_Y));
KC_BUF_X13 D5700 ( .Y(D5700_Y), .A(D5697_Y));
KC_BUF_X13 D4648 ( .Y(D4648_Y), .A(D4643_Y));
KC_BUF_X13 D4087 ( .Y(D4087_Y), .A(D4053_Y));
KC_BUF_X13 D4067 ( .Y(D4067_Y), .A(D4056_Y));
KC_BUF_X13 D4025 ( .Y(D4025_Y), .A(D1521_Y));
KC_BUF_X13 D3984 ( .Y(D3984_Y), .A(D3980_Y));
KC_BUF_X13 D3759 ( .Y(D3759_Y), .A(D3752_Y));
KC_BUF_X13 D2257 ( .Y(D2257_Y), .A(D11345_Y));
KC_BUF_X13 D1807 ( .Y(D1807_Y), .A(D1796_Y));
KC_BUF_X13 D1397 ( .Y(D1397_Y), .A(D13833_Y));
KC_BUF_X13 D1329 ( .Y(D1329_Y), .A(D16702_Y));
KC_BUF_X13 D1328 ( .Y(D1328_Y), .A(D16723_Y));
KC_BUF_X13 D1244 ( .Y(D1244_Y), .A(D13090_Y));
KC_BUF_X13 D713 ( .Y(D713_Y), .A(D6677_Y));
KC_BUF_X13 D712 ( .Y(D712_Y), .A(D6679_Y));
KC_BUF_X13 D711 ( .Y(D711_Y), .A(D707_Y));
KC_BUF_X13 D362 ( .Y(D362_Y), .A(D1794_Y));
KC_BUF_X13 D160 ( .Y(D160_Y), .A(D9627_Y));
KC_AOI22_X2 D15954 ( .A1(D15948_Q), .B0(D14886_Y), .B1(D15949_Q),     .Y(D15954_Y), .A0(D14883_Y));
KC_AOI22_X2 D15953 ( .A1(D15947_Q), .B0(D14884_Y), .B1(D16388_Q),     .Y(D15953_Y), .A0(D14885_Y));
KC_AOI22_X2 D15951 ( .A1(D15992_Q), .B0(D14884_Y), .B1(D1326_Q),     .Y(D15951_Y), .A0(D14885_Y));
KC_AOI22_X2 D15950 ( .A1(D1230_Q), .B0(D14886_Y), .B1(D15994_Q),     .Y(D15950_Y), .A0(D14883_Y));
KC_AOI22_X2 D15876 ( .A1(D15868_Q), .B0(D14886_Y), .B1(D1149_Q),     .Y(D15876_Y), .A0(D14883_Y));
KC_AOI22_X2 D15875 ( .A1(D1148_Q), .B0(D14884_Y), .B1(D16357_Q),     .Y(D15875_Y), .A0(D14885_Y));
KC_AOI22_X2 D15805 ( .A1(D2639_Q), .B0(D1070_Q), .B1(D14884_Y),     .Y(D15805_Y), .A0(D14885_Y));
KC_AOI22_X2 D15804 ( .A1(D14883_Y), .B0(D14886_Y), .B1(D15795_Q),     .Y(D15804_Y), .A0(D14871_Q));
KC_AOI22_X2 D15802 ( .A1(D15668_Q), .B0(D14886_Y), .B1(D1053_Q),     .Y(D15802_Y), .A0(D14883_Y));
KC_AOI22_X2 D15801 ( .A1(D2640_Q), .B0(D14884_Y), .B1(D15796_Q),     .Y(D15801_Y), .A0(D14885_Y));
KC_AOI22_X2 D15799 ( .A1(D15791_Q), .B0(D14886_Y), .B1(D1050_Q),     .Y(D15799_Y), .A0(D14883_Y));
KC_AOI22_X2 D15798 ( .A1(D15792_Q), .B0(D14884_Y), .B1(D16346_Q),     .Y(D15798_Y), .A0(D14885_Y));
KC_AOI22_X2 D15681 ( .A1(D15634_Y), .B0(D879_Y), .B1(D14829_Y),     .Y(D15681_Y), .A0(D2569_Y));
KC_AOI22_X2 D15679 ( .A1(D15634_Y), .B0(D14840_Y), .B1(D13156_Y),     .Y(D15679_Y), .A0(D15629_Y));
KC_AOI22_X2 D15677 ( .A1(D2870_Y), .B0(D14387_Y), .B1(D15616_Y),     .Y(D15677_Y), .A0(D14840_Y));
KC_AOI22_X2 D15676 ( .A1(D15634_Y), .B0(D15662_Y), .B1(D14829_Y),     .Y(D15676_Y), .A0(D15709_Y));
KC_AOI22_X2 D15675 ( .A1(D14829_Y), .B0(D15598_Y), .B1(D15634_Y),     .Y(D15675_Y), .A0(D15659_Y));
KC_AOI22_X2 D15672 ( .A1(D14840_Y), .B0(D15616_Y), .B1(D14187_Y),     .Y(D15672_Y), .A0(D16166_Y));
KC_AOI22_X2 D15671 ( .A1(D15634_Y), .B0(D15660_Y), .B1(D14829_Y),     .Y(D15671_Y), .A0(D2648_Y));
KC_AOI22_X2 D15580 ( .A1(D8886_Y), .B0(D15146_Y), .B1(D15506_Y),     .Y(D15580_Y), .A0(D15529_Y));
KC_AOI22_X2 D15579 ( .A1(D15506_Y), .B0(D9553_Y), .B1(D15529_Y),     .Y(D15579_Y), .A0(D14314_Y));
KC_AOI22_X2 D15578 ( .A1(D755_Y), .B0(D15552_Y), .B1(D14750_Y),     .Y(D15578_Y), .A0(D15416_Y));
KC_AOI22_X2 D15577 ( .A1(D755_Y), .B0(D15416_Y), .B1(D14750_Y),     .Y(D15577_Y), .A0(D15553_Y));
KC_AOI22_X2 D15574 ( .A1(D15529_Y), .B0(D15506_Y), .B1(D14184_Y),     .Y(D15574_Y), .A0(D8997_Y));
KC_AOI22_X2 D15573 ( .A1(D15529_Y), .B0(D15952_Y), .B1(D15506_Y),     .Y(D15573_Y), .A0(D2871_Y));
KC_AOI22_X2 D15572 ( .A1(D14750_Y), .B0(D15599_Y), .B1(D755_Y),     .Y(D15572_Y), .A0(D15410_Y));
KC_AOI22_X2 D15571 ( .A1(D14750_Y), .B0(D15410_Y), .B1(D755_Y),     .Y(D15571_Y), .A0(D15497_Y));
KC_AOI22_X2 D15570 ( .A1(D755_Y), .B0(D15415_Y), .B1(D14750_Y),     .Y(D15570_Y), .A0(D15459_Y));
KC_AOI22_X2 D15148 ( .A1(D15134_Q), .B0(D14886_Y), .B1(D1327_Q),     .Y(D15148_Y), .A0(D14885_Y));
KC_AOI22_X2 D15147 ( .A1(D1377_Q), .B0(D14883_Y), .B1(D15991_Q),     .Y(D15147_Y), .A0(D14884_Y));
KC_AOI22_X2 D15145 ( .A1(D1232_Q), .B0(D14880_Y), .B1(D15217_Q),     .Y(D15145_Y), .A0(D14881_Y));
KC_AOI22_X2 D15081 ( .A1(D1157_Q), .B0(D14886_Y), .B1(D15084_Q),     .Y(D15081_Y), .A0(D14885_Y));
KC_AOI22_X2 D15080 ( .A1(D1163_Q), .B0(D14883_Y), .B1(D15870_Q),     .Y(D15080_Y), .A0(D14884_Y));
KC_AOI22_X2 D15078 ( .A1(D1151_Q), .B0(D14886_Y), .B1(D1153_Q),     .Y(D15078_Y), .A0(D14885_Y));
KC_AOI22_X2 D15077 ( .A1(D14300_Q), .B0(D14883_Y), .B1(D15869_Q),     .Y(D15077_Y), .A0(D14884_Y));
KC_AOI22_X2 D15075 ( .A1(D1158_Q), .B0(D14886_Y), .B1(D15133_Q),     .Y(D15075_Y), .A0(D14885_Y));
KC_AOI22_X2 D15074 ( .A1(D2572_Q), .B0(D14883_Y), .B1(D16010_Q),     .Y(D15074_Y), .A0(D14884_Y));
KC_AOI22_X2 D15002 ( .A1(D14875_Q), .B0(D14886_Y), .B1(D14995_Q),     .Y(D15002_Y), .A0(D14885_Y));
KC_AOI22_X2 D15001 ( .A1(D1052_Q), .B0(D14883_Y), .B1(D924_Q),     .Y(D15001_Y), .A0(D14884_Y));
KC_AOI22_X2 D14999 ( .A1(D14873_Q), .B0(D14886_Y), .B1(D14996_Q),     .Y(D14999_Y), .A0(D14885_Y));
KC_AOI22_X2 D14998 ( .A1(D1051_Q), .B0(D14883_Y), .B1(D15793_Q),     .Y(D14998_Y), .A0(D14884_Y));
KC_AOI22_X2 D14901 ( .A1(D853_Q), .B0(D14879_Y), .B1(D14878_Q),     .Y(D14901_Y), .A0(D14882_Y));
KC_AOI22_X2 D14900 ( .A1(D818_Q), .B0(D14881_Y), .B1(D14814_Q),     .Y(D14900_Y), .A0(D14880_Y));
KC_AOI22_X2 D14897 ( .A1(D14886_Y), .B0(D14815_Q), .B1(D14883_Y),     .Y(D14897_Y), .A0(D14808_Q));
KC_AOI22_X2 D14896 ( .A1(D14886_Y), .B0(D14787_Q), .B1(D14883_Y),     .Y(D14896_Y), .A0(D14788_Q));
KC_AOI22_X2 D14895 ( .A1(D14840_Y), .B0(D14262_Y), .B1(D15616_Y),     .Y(D14895_Y), .A0(D10205_Y));
KC_AOI22_X2 D14894 ( .A1(D14789_Q), .B0(D14884_Y), .B1(D14877_Q),     .Y(D14894_Y), .A0(D14885_Y));
KC_AOI22_X2 D14893 ( .A1(D815_Q), .B0(D14884_Y), .B1(D2573_Q),     .Y(D14893_Y), .A0(D14885_Y));
KC_AOI22_X2 D14891 ( .A1(D14094_Q), .B0(D14879_Y), .B1(D14169_Q),     .Y(D14891_Y), .A0(D14882_Y));
KC_AOI22_X2 D14890 ( .A1(D856_Q), .B0(D14881_Y), .B1(D14091_Q),     .Y(D14890_Y), .A0(D14880_Y));
KC_AOI22_X2 D14888 ( .A1(D14886_Y), .B0(D14883_Y), .B1(D2517_Q),     .Y(D14888_Y), .A0(D820_Q));
KC_AOI22_X2 D14887 ( .A1(D14790_Q), .B0(D14884_Y), .B1(D14876_Q),     .Y(D14887_Y), .A0(D14885_Y));
KC_AOI22_X2 D14798 ( .A1(D14750_Y), .B0(D14380_Y), .B1(D15506_Y),     .Y(D14798_Y), .A0(D14672_Y));
KC_AOI22_X2 D14797 ( .A1(D755_Y), .B0(D15529_Y), .B1(D16132_Y),     .Y(D14797_Y), .A0(D757_Y));
KC_AOI22_X2 D14795 ( .A1(D15529_Y), .B0(D2578_Y), .B1(D15506_Y),     .Y(D14795_Y), .A0(D15437_Y));
KC_AOI22_X2 D14794 ( .A1(D755_Y), .B0(D15424_Y), .B1(D14750_Y),     .Y(D14794_Y), .A0(D14672_Y));
KC_AOI22_X2 D14395 ( .A1(D15216_Q), .B0(D14879_Y), .B1(D15232_Q),     .Y(D14395_Y), .A0(D14882_Y));
KC_AOI22_X2 D14394 ( .A1(D14490_Q), .B0(D14881_Y), .B1(D14475_Q),     .Y(D14394_Y), .A0(D14879_Y));
KC_AOI22_X2 D14393 ( .A1(D14374_Q), .B0(D14880_Y), .B1(D15214_Q),     .Y(D14393_Y), .A0(D14881_Y));
KC_AOI22_X2 D14391 ( .A1(D14375_Q), .B0(D14880_Y), .B1(D13771_Q),     .Y(D14391_Y), .A0(D14882_Y));
KC_AOI22_X2 D14389 ( .A1(D13762_Q), .B0(D14880_Y), .B1(D13816_Q),     .Y(D14389_Y), .A0(D14881_Y));
KC_AOI22_X2 D14388 ( .A1(D13809_Q), .B0(D14879_Y), .B1(D13807_Q),     .Y(D14388_Y), .A0(D14882_Y));
KC_AOI22_X2 D14385 ( .A1(D2524_Q), .B0(D14880_Y), .B1(D15218_Q),     .Y(D14385_Y), .A0(D14882_Y));
KC_AOI22_X2 D14384 ( .A1(D2523_Q), .B0(D14880_Y), .B1(D15215_Q),     .Y(D14384_Y), .A0(D14882_Y));
KC_AOI22_X2 D14383 ( .A1(D1376_Q), .B0(D14881_Y), .B1(D1323_Q),     .Y(D14383_Y), .A0(D14879_Y));
KC_AOI22_X2 D14382 ( .A1(D15229_Q), .B0(D14881_Y), .B1(D15212_Q),     .Y(D14382_Y), .A0(D14879_Y));
KC_AOI22_X2 D14379 ( .A1(D13804_Q), .B0(D14881_Y), .B1(D13811_Q),     .Y(D14379_Y), .A0(D14879_Y));
KC_AOI22_X2 D14378 ( .A1(D13761_Q), .B0(D14880_Y), .B1(D13815_Q),     .Y(D14378_Y), .A0(D14881_Y));
KC_AOI22_X2 D14377 ( .A1(D13814_Q), .B0(D14879_Y), .B1(D1321_Q),     .Y(D14377_Y), .A0(D14882_Y));
KC_AOI22_X2 D14376 ( .A1(D13764_Q), .B0(D14880_Y), .B1(D13760_Q),     .Y(D14376_Y), .A0(D14882_Y));
KC_AOI22_X2 D14313 ( .A1(D13705_Q), .B0(D14879_Y), .B1(D13704_Q),     .Y(D14313_Y), .A0(D14882_Y));
KC_AOI22_X2 D14312 ( .A1(D1159_Q), .B0(D14880_Y), .B1(D164_Q),     .Y(D14312_Y), .A0(D14881_Y));
KC_AOI22_X2 D14310 ( .A1(D13765_Q), .B0(D14880_Y), .B1(D2468_Q),     .Y(D14310_Y), .A0(D14882_Y));
KC_AOI22_X2 D14309 ( .A1(D1235_Q), .B0(D14881_Y), .B1(D1150_Q),     .Y(D14309_Y), .A0(D14879_Y));
KC_AOI22_X2 D14261 ( .A1(D14238_Q), .B0(D14879_Y), .B1(D13051_Q),     .Y(D14261_Y), .A0(D14882_Y));
KC_AOI22_X2 D14260 ( .A1(D13050_Q), .B0(D14881_Y), .B1(D13703_Q),     .Y(D14260_Y), .A0(D14880_Y));
KC_AOI22_X2 D14190 ( .A1(D14093_Q), .B0(D14881_Y), .B1(D14117_Q),     .Y(D14190_Y), .A0(D14880_Y));
KC_AOI22_X2 D14189 ( .A1(D14880_Y), .B0(D14118_Q), .B1(D14881_Y),     .Y(D14189_Y), .A0(D817_Q));
KC_AOI22_X2 D14188 ( .A1(D14092_Q), .B0(D14879_Y), .B1(D14170_Q),     .Y(D14188_Y), .A0(D14882_Y));
KC_AOI22_X2 D14186 ( .A1(D928_Q), .B0(D14880_Y), .B1(D12991_Q),     .Y(D14186_Y), .A0(D14882_Y));
KC_AOI22_X2 D14185 ( .A1(D12997_Q), .B0(D14881_Y), .B1(D12919_Q),     .Y(D14185_Y), .A0(D14879_Y));
KC_AOI22_X2 D14183 ( .A1(D930_Q), .B0(D14879_Y), .B1(D2391_Q),     .Y(D14183_Y), .A0(D14882_Y));
KC_AOI22_X2 D14182 ( .A1(D954_Q), .B0(D14880_Y), .B1(D12995_Q),     .Y(D14182_Y), .A0(D14881_Y));
KC_AOI22_X2 D14180 ( .A1(D13530_Q), .B0(D14879_Y), .B1(D12994_Q),     .Y(D14180_Y), .A0(D14882_Y));
KC_AOI22_X2 D14179 ( .A1(D12921_Q), .B0(D14880_Y), .B1(D12992_Q),     .Y(D14179_Y), .A0(D14881_Y));
KC_AOI22_X2 D11667 ( .A1(D11665_Y), .B0(D11652_Y), .B1(D11669_Y),     .Y(D11667_Y), .A0(D612_Y));
KC_AOI22_X2 D11666 ( .A1(D11674_Y), .B0(D12201_Y), .B1(D11675_Y),     .Y(D11666_Y), .A0(D11651_Y));
KC_AOI22_X2 D9335 ( .A1(D490_Y), .B0(D6077_Y), .B1(D9353_Q),     .Y(D9335_Y), .A0(D9181_Y));
KC_AOI22_X2 D9331 ( .A1(D9319_Q), .B0(D9114_Y), .B1(D483_Q),     .Y(D9331_Y), .A0(D7631_Y));
KC_AOI22_X2 D9330 ( .A1(D7822_Y), .B0(D6077_Y), .B1(D9323_Q),     .Y(D9330_Y), .A0(D9181_Y));
KC_AOI22_X2 D9329 ( .A1(D9336_Q), .B0(D9114_Y), .B1(D482_Q),     .Y(D9329_Y), .A0(D7631_Y));
KC_AOI22_X2 D9328 ( .A1(D9324_Q), .B0(D9114_Y), .B1(D7894_Q),     .Y(D9328_Y), .A0(D7631_Y));
KC_AOI22_X2 D9327 ( .A1(D465_Y), .B0(D6077_Y), .B1(D9318_Q),     .Y(D9327_Y), .A0(D9181_Y));
KC_AOI22_X2 D9157 ( .A1(D7638_Y), .B0(D9114_Y), .B1(D9278_Q),     .Y(D9157_Y), .A0(D386_Q));
KC_AOI22_X2 D9156 ( .A1(D9260_Q), .B0(D9102_Y), .B1(D8711_Q),     .Y(D9156_Y), .A0(D7631_Y));
KC_AOI22_X2 D9154 ( .A1(D7638_Y), .B0(D9114_Y), .B1(D2092_Q),     .Y(D9154_Y), .A0(D7667_Q));
KC_AOI22_X2 D9153 ( .A1(D9209_Q), .B0(D9102_Y), .B1(D8709_Q),     .Y(D9153_Y), .A0(D7631_Y));
KC_AOI22_X2 D8957 ( .A1(D2070_Y), .B0(D7479_Q), .B1(D7393_Y),     .Y(D8957_Y), .A0(D8954_Q));
KC_AOI22_X2 D8956 ( .A1(D727_Y), .B0(D10006_Q), .B1(D9990_Y),     .Y(D8956_Y), .A0(D8900_Y));
KC_AOI22_X2 D8720 ( .A1(D8689_S), .B0(D8716_Y), .B1(D8677_Y),     .Y(D8720_Y), .A0(D8694_Y));
KC_AOI22_X2 D8719 ( .A1(D8733_Y), .B0(D8678_Y), .B1(D8684_Y),     .Y(D8719_Y), .A0(D8685_Y));
KC_AOI22_X2 D8252 ( .A1(D8225_Y), .B0(D8239_Y), .B1(D8226_Y),     .Y(D8252_Y), .A0(D9559_Y));
KC_AOI22_X2 D8251 ( .A1(D8224_Y), .B0(D8241_Y), .B1(D8215_Y),     .Y(D8251_Y), .A0(D8234_Y));
KC_AOI22_X2 D7665 ( .A1(D343_Y), .B0(D7545_Y), .B1(D6175_Y),     .Y(D7665_Y), .A0(D12764_Y));
KC_AOI22_X2 D7664 ( .A1(D1923_Y), .B0(D6264_Y), .B1(D7654_Y),     .Y(D7664_Y), .A0(D6177_Y));
KC_AOI22_X2 D7663 ( .A1(D343_Y), .B0(D7545_Y), .B1(D9210_Y),     .Y(D7663_Y), .A0(D13280_Q));
KC_AOI22_X2 D7661 ( .A1(D7135_Y), .B0(D6264_Y), .B1(D4720_Y),     .Y(D7661_Y), .A0(D6177_Y));
KC_AOI22_X2 D7611 ( .A1(D343_Y), .B0(D7545_Y), .B1(D1925_Y),     .Y(D7611_Y), .A0(D12763_Y));
KC_AOI22_X2 D7607 ( .A1(D343_Y), .B0(D6177_Y), .B1(D7522_Y),     .Y(D7607_Y), .A0(D13289_Y));
KC_AOI22_X2 D7606 ( .A1(D4630_Y), .B0(D7545_Y), .B1(D8703_Y),     .Y(D7606_Y), .A0(D6264_Y));
KC_AOI22_X2 D7605 ( .A1(D343_Y), .B0(D7545_Y), .B1(D6174_Y),     .Y(D7605_Y), .A0(D12300_Y));
KC_AOI22_X2 D7602 ( .A1(D7581_Y), .B0(D6264_Y), .B1(D6286_Y),     .Y(D7602_Y), .A0(D6177_Y));
KC_AOI22_X2 D7601 ( .A1(D7521_Y), .B0(D6264_Y), .B1(D7617_Y),     .Y(D7601_Y), .A0(D6177_Y));
KC_AOI22_X2 D7600 ( .A1(D343_Y), .B0(D7545_Y), .B1(D4551_Y),     .Y(D7600_Y), .A0(D723_Q));
KC_AOI22_X2 D7598 ( .A1(D343_Y), .B0(D7545_Y), .B1(D6185_Y),     .Y(D7598_Y), .A0(D13288_Y));
KC_AOI22_X2 D7597 ( .A1(D7656_Y), .B0(D6264_Y), .B1(D7584_Y),     .Y(D7597_Y), .A0(D6177_Y));
KC_AOI22_X2 D7596 ( .A1(D343_Y), .B0(D7545_Y), .B1(D5949_Y),     .Y(D7596_Y), .A0(D725_Y));
KC_AOI22_X2 D7594 ( .A1(D6170_Y), .B0(D6264_Y), .B1(D1825_Y),     .Y(D7594_Y), .A0(D6177_Y));
KC_AOI22_X2 D7593 ( .A1(D343_Y), .B0(D7545_Y), .B1(D1677_Y),     .Y(D7593_Y), .A0(D724_Y));
KC_AOI22_X2 D7591 ( .A1(D4807_Y), .B0(D6264_Y), .B1(D9264_Y),     .Y(D7591_Y), .A0(D6177_Y));
KC_AOI22_X2 D7590 ( .A1(D343_Y), .B0(D7545_Y), .B1(D7588_Y),     .Y(D7590_Y), .A0(D12762_Y));
KC_AOI22_X2 D7157 ( .A1(D182_Y), .B0(D7114_Y), .B1(D181_Y),     .Y(D7157_Y), .A0(D8704_Y));
KC_AOI22_X2 D7155 ( .A1(D181_Y), .B0(D7160_Y), .B1(D8704_Y),     .Y(D7155_Y), .A0(D7160_Y));
KC_AOI22_X2 D7154 ( .A1(D7113_Y), .B0(D8704_Y), .B1(D7125_Y),     .Y(D7154_Y), .A0(D7160_Y));
KC_AOI22_X2 D6347 ( .A1(D6315_Y), .B0(D6325_Y), .B1(D6268_Y),     .Y(D6347_Y), .A0(D6330_Y));
KC_AOI22_X2 D6346 ( .A1(D7564_Y), .B0(D6326_Y), .B1(D6305_Y),     .Y(D6346_Y), .A0(D6296_Y));
KC_AOI22_X2 D6270 ( .A1(D7136_Y), .B0(D6264_Y), .B1(D9223_Y),     .Y(D6270_Y), .A0(D6177_Y));
KC_AOI22_X2 D6195 ( .A1(D4804_Y), .B0(D6264_Y), .B1(D1771_Y),     .Y(D6195_Y), .A0(D6177_Y));
KC_AOI22_X2 D6193 ( .A1(D6184_Y), .B0(D6117_Y), .B1(D6182_Y),     .Y(D6193_Y), .A0(D6151_Y));
KC_AOI22_X2 D6192 ( .A1(D6253_Y), .B0(D6145_Y), .B1(D6147_Y),     .Y(D6192_Y), .A0(D6204_Y));
KC_AOI22_X2 D6190 ( .A1(D6171_Y), .B0(D6264_Y), .B1(D6173_Y),     .Y(D6190_Y), .A0(D6177_Y));
KC_AOI22_X2 D6189 ( .A1(D6209_Y), .B0(D6264_Y), .B1(D6169_Y),     .Y(D6189_Y), .A0(D6177_Y));
KC_AOI22_X2 D6187 ( .A1(D4628_Y), .B0(D6264_Y), .B1(D16754_Y),     .Y(D6187_Y), .A0(D6177_Y));
KC_AOI22_X2 D5081 ( .A1(D3446_Y), .B0(D3406_Y), .B1(D4900_Y),     .Y(D5081_Y), .A0(D4891_Y));
KC_AOI22_X2 D4126 ( .A1(D4421_Y), .B0(D4149_Q), .B1(D4097_Y),     .Y(D4126_Y), .A0(D4120_Q));
KC_AOI22_X2 D4125 ( .A1(D4118_Q), .B0(D8313_Q), .B1(D4096_Y),     .Y(D4125_Y), .A0(D4440_Y));
KC_AOI22_X2 D3581 ( .A1(D3409_Y), .B0(D5044_Y), .B1(D3553_Y),     .Y(D3581_Y), .A0(D4916_Y));
KC_AOI22_X2 D3286 ( .A1(D3289_Y), .B0(D3242_Y), .B1(D3292_Y),     .Y(D3286_Y), .A0(D3207_Y));
KC_AOI22_X2 D3285 ( .A1(D3260_S), .B0(D3291_Y), .B1(D3244_Y),     .Y(D3285_Y), .A0(D3223_Y));
KC_AOI22_X2 D3089 ( .A1(D3042_Y), .B0(D3042_Y), .B1(D3021_Y),     .Y(D3089_Y), .A0(D3019_Y));
KC_AOI22_X2 D3088 ( .A1(D3053_Y), .B0(D3053_Y), .B1(D3062_Y),     .Y(D3088_Y), .A0(D3064_Y));
KC_AOI22_X2 D2646 ( .A1(D15873_Q), .B0(D14886_Y), .B1(D16363_Q),     .Y(D2646_Y), .A0(D14883_Y));
KC_AOI22_X2 D2645 ( .A1(D144_Q), .B0(D14884_Y), .B1(D1156_Q),     .Y(D2645_Y), .A0(D14885_Y));
KC_AOI22_X2 D2643 ( .A1(D1233_Q), .B0(D14884_Y), .B1(D142_Q),     .Y(D2643_Y), .A0(D14885_Y));
KC_AOI22_X2 D2642 ( .A1(D2638_Q), .B0(D14886_Y), .B1(D1234_Q),     .Y(D2642_Y), .A0(D14883_Y));
KC_AOI22_X2 D2582 ( .A1(D14885_Y), .B0(D14266_Q), .B1(D14886_Y),     .Y(D2582_Y), .A0(D952_Q));
KC_AOI22_X2 D2581 ( .A1(D1065_Q), .B0(D14883_Y), .B1(D14903_Q),     .Y(D2581_Y), .A0(D14884_Y));
KC_AOI22_X2 D2580 ( .A1(D143_Q), .B0(D14883_Y), .B1(D15874_Q),     .Y(D2580_Y), .A0(D14884_Y));
KC_AOI22_X2 D2577 ( .A1(D14263_Q), .B0(D14886_Y), .B1(D1048_Q),     .Y(D2577_Y), .A0(D14885_Y));
KC_AOI22_X2 D2576 ( .A1(D13706_Q), .B0(D14886_Y), .B1(D1152_Q),     .Y(D2576_Y), .A0(D14883_Y));
KC_AOI22_X2 D2575 ( .A1(D13711_Q), .B0(D14884_Y), .B1(D1147_Q),     .Y(D2575_Y), .A0(D14885_Y));
KC_AOI22_X2 D2520 ( .A1(D12996_Q), .B0(D14881_Y), .B1(D12918_Q),     .Y(D2520_Y), .A0(D14880_Y));
KC_AOI22_X2 D2097 ( .A1(D382_Y), .B0(D8665_Y), .B1(D8732_Y),     .Y(D2097_Y), .A0(D8806_Y));
KC_AOI22_X2 D2096 ( .A1(D8666_Y), .B0(D8787_Y), .B1(D8666_Y),     .Y(D2096_Y), .A0(D8665_Y));
KC_AOI22_X2 D1951 ( .A1(D7134_Y), .B0(D6264_Y), .B1(D7652_Y),     .Y(D1951_Y), .A0(D6177_Y));
KC_AOI22_X2 D1950 ( .A1(D343_Y), .B0(D7545_Y), .B1(D7723_Y),     .Y(D1950_Y), .A0(D12301_Y));
KC_AOI22_X2 D1948 ( .A1(D7727_Y), .B0(D6264_Y), .B1(D6261_Y),     .Y(D1948_Y), .A0(D6177_Y));
KC_AOI22_X2 D1803 ( .A1(D1008_Y), .B0(D6264_Y), .B1(D107_Y),     .Y(D1803_Y), .A0(D6177_Y));
KC_AOI22_X2 D1802 ( .A1(D343_Y), .B0(D7545_Y), .B1(D6360_Y),     .Y(D1802_Y), .A0(D12761_Y));
KC_AOI22_X2 D1239 ( .A1(D1325_Q), .B0(D14879_Y), .B1(D15213_Q),     .Y(D1239_Y), .A0(D14882_Y));
KC_AOI22_X2 D939 ( .A1(D14109_Q), .B0(D14879_Y), .B1(D14168_Q),     .Y(D939_Y), .A0(D14882_Y));
KC_AOI22_X2 D938 ( .A1(D14829_Y), .B0(D14392_Y), .B1(D15616_Y),     .Y(D938_Y), .A0(D2569_Y));
KC_AOI22_X2 D937 ( .A1(D12139_Y), .B0(D14386_Y), .B1(D15616_Y),     .Y(D937_Y), .A0(D14840_Y));
KC_AOI22_X2 D832 ( .A1(D15438_Y), .B0(D14396_Y), .B1(D15506_Y),     .Y(D832_Y), .A0(D15529_Y));
KC_AOI22_X2 D388 ( .A1(D343_Y), .B0(D7545_Y), .B1(D378_Y), .Y(D388_Y),     .A0(D13171_Y));
KC_AOI22_X2 D359 ( .A1(D343_Y), .B0(D7545_Y), .B1(D5930_Y), .Y(D359_Y),     .A0(D13287_Y));
KC_AOI22_X2 D357 ( .A1(D343_Y), .B0(D7545_Y), .B1(D6337_Y), .Y(D357_Y),     .A0(D12863_Y));
KC_AOI22_X2 D197 ( .A1(D7127_Y), .B0(D7125_Y), .B1(D182_Y), .Y(D197_Y),     .A0(D7160_Y));
KC_AOI22_X2 D159 ( .A1(D343_Y), .B0(D7545_Y), .B1(D6257_Y), .Y(D159_Y),     .A0(D13285_Y));
KC_AOI22_X2 D158 ( .A1(D14165_Q), .B0(D14879_Y), .B1(D12993_Q),     .Y(D158_Y), .A0(D14882_Y));
KC_NOR2_X5 D16728 ( .Y(D16728_Y), .B(D16725_Y), .A(D16726_Y));
KC_NOR2_X5 D16723 ( .Y(D16723_Y), .B(D16725_Y), .A(D16721_Y));
KC_NOR2_X5 D16703 ( .Y(D16703_Y), .B(D16714_Y), .A(D16698_Y));
KC_NOR2_X5 D16702 ( .Y(D16702_Y), .B(D16714_Y), .A(D16699_Y));
KC_NOR2_X5 D16630 ( .Y(D16630_Y), .B(D16644_Y), .A(D16637_Y));
KC_NOR2_X5 D16620 ( .Y(D16620_Y), .B(D16644_Y), .A(D16621_Y));
KC_NOR2_X5 D16593 ( .Y(D16593_Y), .B(D16589_Y), .A(D16584_Y));
KC_NOR2_X5 D16580 ( .Y(D16580_Y), .B(D16589_Y), .A(D16577_Y));
KC_NOR2_X5 D16327 ( .Y(D16327_Y), .B(D16342_Y), .A(D16312_Y));
KC_NOR2_X5 D16323 ( .Y(D16323_Y), .B(D16342_Y), .A(GND));
KC_NOR2_X5 D15137 ( .Y(D15137_Y), .B(D15157_Y), .A(D15130_Y));
KC_NOR2_X5 D15136 ( .Y(D15136_Y), .B(D15157_Y), .A(D15129_Y));
KC_NOR2_X5 D14793 ( .Y(D14793_Y), .B(D14804_Y), .A(D14784_Y));
KC_NOR2_X5 D14792 ( .Y(D14792_Y), .B(D14804_Y), .A(D14680_Y));
KC_NOR2_X5 D14247 ( .Y(D14247_Y), .B(D14134_Y), .A(D874_Y));
KC_NOR2_X5 D13833 ( .Y(D13833_Y), .B(D13844_Y), .A(D13821_Y));
KC_NOR2_X5 D13831 ( .Y(D13831_Y), .B(D13844_Y), .A(D13822_Y));
KC_NOR2_X5 D13617 ( .Y(D13617_Y), .B(D13009_Y), .A(D13608_Y));
KC_NOR2_X5 D13613 ( .Y(D13613_Y), .B(D13009_Y), .A(D13606_Y));
KC_NOR2_X5 D13090 ( .Y(D13090_Y), .B(D13093_Y), .A(D13084_Y));
KC_NOR2_X5 D12365 ( .Y(D12365_Y), .B(D12308_Y), .A(D12271_Y));
KC_NOR2_X5 D12282 ( .Y(D12282_Y), .B(D12308_Y), .A(D12338_Y));
KC_NOR2_X5 D12125 ( .Y(D12125_Y), .B(D11611_Y), .A(D12118_Y));
KC_NOR2_X5 D12051 ( .Y(D12051_Y), .B(D11964_Y), .A(D11957_Y));
KC_NOR2_X5 D12050 ( .Y(D12050_Y), .B(D11965_Y), .A(D11957_Y));
KC_NOR2_X5 D11930 ( .Y(D11930_Y), .B(D11959_Y), .A(D11941_Y));
KC_NOR2_X5 D11929 ( .Y(D11929_Y), .B(D1108_Y), .A(D11946_Y));
KC_NOR2_X5 D11599 ( .Y(D11599_Y), .B(D11611_Y), .A(D11596_Y));
KC_NOR2_X5 D11345 ( .Y(D11345_Y), .B(D11418_Y), .A(D11332_Y));
KC_NOR2_X5 D11040 ( .Y(D11040_Y), .B(D11054_Y), .A(D11028_Y));
KC_NOR2_X5 D11038 ( .Y(D11038_Y), .B(D11054_Y), .A(D11032_Y));
KC_NOR2_X5 D11009 ( .Y(D11009_Y), .B(D10983_Y), .A(D10964_Y));
KC_NOR2_X5 D10816 ( .Y(D10816_Y), .B(D10829_Y), .A(D10798_Y));
KC_NOR2_X5 D10812 ( .Y(D10812_Y), .B(D10829_Y), .A(D10795_Y));
KC_NOR2_X5 D10809 ( .Y(D10809_Y), .B(D10761_Y), .A(D10729_Y));
KC_NOR2_X5 D10808 ( .Y(D10808_Y), .B(D10762_Y), .A(D10729_Y));
KC_NOR2_X5 D10634 ( .Y(D10634_Y), .B(D9012_Y), .A(D2162_Y));
KC_NOR2_X5 D10559 ( .Y(D10559_Y), .B(D10479_Y), .A(D10965_Y));
KC_NOR2_X5 D10558 ( .Y(D10558_Y), .B(D10486_Y), .A(D10965_Y));
KC_NOR2_X5 D10169 ( .Y(D10169_Y), .B(D208_Y), .A(D2162_Y));
KC_NOR2_X5 D10151 ( .Y(D10151_Y), .B(D2162_Y), .A(D10152_Y));
KC_NOR2_X5 D10127 ( .Y(D10127_Y), .B(D10057_Y), .A(D10128_Y));
KC_NOR2_X5 D10124 ( .Y(D10124_Y), .B(D10057_Y), .A(D10125_Y));
KC_NOR2_X5 D10122 ( .Y(D10122_Y), .B(D10057_Y), .A(D10123_Y));
KC_NOR2_X5 D10121 ( .Y(D10121_Y), .B(D10057_Y), .A(D10120_Y));
KC_NOR2_X5 D10119 ( .Y(D10119_Y), .B(D10057_Y), .A(D10118_Y));
KC_NOR2_X5 D9916 ( .Y(D9916_Y), .B(D8662_Y), .A(D9907_Y));
KC_NOR2_X5 D9913 ( .Y(D9913_Y), .B(D8662_Y), .A(D9901_Y));
KC_NOR2_X5 D9718 ( .Y(D9718_Y), .B(D9721_Y), .A(D9715_Y));
KC_NOR2_X5 D9627 ( .Y(D9627_Y), .B(D9721_Y), .A(D9716_Y));
KC_NOR2_X5 D8600 ( .Y(D8600_Y), .B(D8608_Y), .A(D8586_Y));
KC_NOR2_X5 D8599 ( .Y(D8599_Y), .B(D8608_Y), .A(D8592_Y));
KC_NOR2_X5 D8346 ( .Y(D8346_Y), .B(D8351_Y), .A(D8048_Y));
KC_NOR2_X5 D8345 ( .Y(D8345_Y), .B(D8351_Y), .A(D8290_Y));
KC_NOR2_X5 D8344 ( .Y(D8344_Y), .B(D8289_Y), .A(D8288_Y));
KC_NOR2_X5 D8153 ( .Y(D8153_Y), .B(D9518_Y), .A(D8254_Y));
KC_NOR2_X5 D7660 ( .Y(D7660_Y), .B(D481_Y), .A(D346_Y));
KC_NOR2_X5 D7393 ( .Y(D7393_Y), .B(D7323_Y), .A(D7460_Y));
KC_NOR2_X5 D6974 ( .Y(D6974_Y), .B(D6942_Y), .A(D6923_Y));
KC_NOR2_X5 D6973 ( .Y(D6973_Y), .B(D6943_Y), .A(D6923_Y));
KC_NOR2_X5 D6760 ( .Y(D6760_Y), .B(D5294_Y), .A(D5260_Y));
KC_NOR2_X5 D6679 ( .Y(D6679_Y), .B(D8165_Y), .A(D6664_Y));
KC_NOR2_X5 D6677 ( .Y(D6677_Y), .B(D8165_Y), .A(D6654_Y));
KC_NOR2_X5 D6560 ( .Y(D6560_Y), .B(D6567_Y), .A(D6545_Y));
KC_NOR2_X5 D6559 ( .Y(D6559_Y), .B(D6567_Y), .A(D6541_Y));
KC_NOR2_X5 D6396 ( .Y(D6396_Y), .B(D6413_Y), .A(D6378_Y));
KC_NOR2_X5 D6393 ( .Y(D6393_Y), .B(D6413_Y), .A(D6377_Y));
KC_NOR2_X5 D6268 ( .Y(D6268_Y), .B(D10162_Y), .A(D7563_Y));
KC_NOR2_X5 D6186 ( .Y(D6186_Y), .B(D7785_Y), .A(D7564_Y));
KC_NOR2_X5 D27 ( .Y(D27_Y), .B(D30_Y), .A(D4478_Y));
KC_NOR2_X5 D6075 ( .Y(D6075_Y), .B(D243_Y), .A(D1872_Y));
KC_NOR2_X5 D5809 ( .Y(D5809_Y), .B(D5822_Y), .A(D5801_Y));
KC_NOR2_X5 D5697 ( .Y(D5697_Y), .B(D5822_Y), .A(D5681_Y));
KC_NOR2_X5 D5542 ( .Y(D5542_Y), .B(D1597_Y), .A(D5510_Y));
KC_NOR2_X5 D5484 ( .Y(D5484_Y), .B(D5490_Y), .A(D5473_Y));
KC_NOR2_X5 D4643 ( .Y(D4643_Y), .B(D1818_Y), .A(D1646_Y));
KC_NOR2_X5 D4056 ( .Y(D4056_Y), .B(D4073_Y), .A(D4046_Y));
KC_NOR2_X5 D4053 ( .Y(D4053_Y), .B(D4073_Y), .A(D4084_Y));
KC_NOR2_X5 D3980 ( .Y(D3980_Y), .B(D1535_Y), .A(D3970_Y));
KC_NOR2_X5 D3752 ( .Y(D3752_Y), .B(D5253_Y), .A(D3730_Y));
KC_NOR2_X5 D2402 ( .Y(D2402_Y), .B(D13093_Y), .A(D2386_Y));
KC_NOR2_X5 D1945 ( .Y(D1945_Y), .B(D8017_Y), .A(D2343_Y));
KC_NOR2_X5 D1801 ( .Y(D1801_Y), .B(D5372_Y), .A(D6782_Y));
KC_NOR2_X5 D1796 ( .Y(D1796_Y), .B(D30_Y), .A(D4479_Y));
KC_NOR2_X5 D1794 ( .Y(D1794_Y), .B(D1818_Y), .A(D6262_Y));
KC_NOR2_X5 D1660 ( .Y(D1660_Y), .B(D5490_Y), .A(D5477_Y));
KC_NOR2_X5 D1521 ( .Y(D1521_Y), .B(D1535_Y), .A(D1492_Y));
KC_NOR2_X5 D935 ( .Y(D935_Y), .B(D11418_Y), .A(D11331_Y));
KC_NOR2_X5 D707 ( .Y(D707_Y), .B(D5253_Y), .A(D3729_Y));
KC_NOR2_X5 D157 ( .Y(D157_Y), .B(D6795_Y), .A(D5259_Y));
KC_OR2_X2 D16727 ( .Y(D16727_Y), .B(D16715_Y), .A(D16732_Y));
KC_OR2_X2 D16706 ( .Y(D16706_Y), .B(D16772_Y), .A(D16707_Y));
KC_OR2_X2 D16631 ( .Y(D16631_Y), .B(D16639_Y), .A(D16628_Y));
KC_OR2_X2 D16616 ( .Y(D16616_Y), .B(D16639_Y), .A(D16619_Y));
KC_OR2_X2 D16552 ( .Y(D16552_Y), .B(D16588_Y), .A(D16553_Y));
KC_OR2_X2 D16324 ( .Y(D16324_Y), .B(D16469_Y), .A(D16294_Y));
KC_OR2_X2 D16322 ( .Y(D16322_Y), .B(D16341_Y), .A(D16326_Y));
KC_OR2_X2 D15141 ( .Y(D15141_Y), .B(D15159_Y), .A(D15142_Y));
KC_OR2_X2 D15140 ( .Y(D15140_Y), .B(D15159_Y), .A(D15135_Y));
KC_OR2_X2 D14696 ( .Y(D14696_Y), .B(D14712_Y), .A(D14791_Y));
KC_OR2_X2 D14695 ( .Y(D14695_Y), .B(D14712_Y), .A(D14697_Y));
KC_OR2_X2 D13829 ( .Y(D13829_Y), .B(D13843_Y), .A(D13830_Y));
KC_OR2_X2 D13828 ( .Y(D13828_Y), .B(D13843_Y), .A(D13832_Y));
KC_OR2_X2 D13614 ( .Y(D13614_Y), .B(D1076_Y), .A(D13615_Y));
KC_OR2_X2 D13611 ( .Y(D13611_Y), .B(D1076_Y), .A(D13612_Y));
KC_OR2_X2 D12549 ( .Y(D12549_Y), .B(D13094_Y), .A(D12548_Y));
KC_OR2_X2 D12285 ( .Y(D12285_Y), .B(D12304_Y), .A(D12284_Y));
KC_OR2_X2 D12283 ( .Y(D12283_Y), .B(D12304_Y), .A(D12293_Y));
KC_OR2_X2 D11629 ( .Y(D11629_Y), .B(D11673_Q), .A(D11639_Q));
KC_OR2_X2 D11604 ( .Y(D11604_Y), .B(D11612_Y), .A(D11603_Y));
KC_OR2_X2 D11600 ( .Y(D11600_Y), .B(D11612_Y), .A(D11598_Y));
KC_OR2_X2 D11408 ( .Y(D11408_Y), .B(D11417_Y), .A(D11407_Y));
KC_OR2_X2 D11346 ( .Y(D11346_Y), .B(D11417_Y), .A(D11347_Y));
KC_OR2_X2 D11046 ( .Y(D11046_Y), .B(D11055_Y), .A(D11037_Y));
KC_OR2_X2 D11042 ( .Y(D11042_Y), .B(D11055_Y), .A(D11041_Y));
KC_OR2_X2 D10817 ( .Y(D10817_Y), .B(D16082_Y), .A(D10810_Y));
KC_OR2_X2 D10813 ( .Y(D10813_Y), .B(D16082_Y), .A(D10814_Y));
KC_OR2_X2 D9915 ( .Y(D9915_Y), .B(D8663_Y), .A(D9914_Y));
KC_OR2_X2 D9719 ( .Y(D9719_Y), .B(D8478_Y), .A(D9720_Y));
KC_OR2_X2 D8659 ( .Y(D8659_Y), .B(D8663_Y), .A(D8660_Y));
KC_OR2_X2 D8598 ( .Y(D8598_Y), .B(D8607_Y), .A(D1238_Y));
KC_OR2_X2 D8467 ( .Y(D8467_Y), .B(D8478_Y), .A(D8468_Y));
KC_OR2_X2 D7974 ( .Y(D7974_Y), .B(D7975_Y), .A(D7929_Y));
KC_OR2_X2 D7016 ( .Y(D7016_Y), .B(D8607_Y), .A(D7015_Y));
KC_OR2_X2 D6678 ( .Y(D6678_Y), .B(D16753_Y), .A(D6680_Y));
KC_OR2_X2 D6676 ( .Y(D6676_Y), .B(D16753_Y), .A(D6682_Y));
KC_OR2_X2 D6557 ( .Y(D6557_Y), .B(D16696_Y), .A(D6565_Y));
KC_OR2_X2 D6397 ( .Y(D6397_Y), .B(D14591_Y), .A(D6395_Y));
KC_OR2_X2 D6394 ( .Y(D6394_Y), .B(D14591_Y), .A(D6388_Y));
KC_OR2_X2 D6124 ( .Y(D6124_Y), .B(D6128_Y), .A(D6121_Y));
KC_OR2_X2 D5810 ( .Y(D5810_Y), .B(D6275_Y), .A(D5696_Y));
KC_OR2_X2 D5694 ( .Y(D5694_Y), .B(D6275_Y), .A(D5695_Y));
KC_OR2_X2 D5482 ( .Y(D5482_Y), .B(D5489_Y), .A(D5483_Y));
KC_OR2_X2 D4644 ( .Y(D4644_Y), .B(D6197_Y), .A(D4646_Y));
KC_OR2_X2 D4058 ( .Y(D4058_Y), .B(D4072_Y), .A(D4055_Y));
KC_OR2_X2 D4054 ( .Y(D4054_Y), .B(D4072_Y), .A(D4052_Y));
KC_OR2_X2 D4020 ( .Y(D4020_Y), .B(D4571_Y), .A(D4021_Y));
KC_OR2_X2 D3981 ( .Y(D3981_Y), .B(D4571_Y), .A(D3982_Y));
KC_OR2_X2 D3753 ( .Y(D3753_Y), .B(D4406_Y), .A(D3760_Y));
KC_OR2_X2 D3750 ( .Y(D3750_Y), .B(D4406_Y), .A(D3751_Y));
KC_OR2_X2 D2696 ( .Y(D2696_Y), .B(D16715_Y), .A(D16724_Y));
KC_OR2_X2 D2359 ( .Y(D2359_Y), .B(D13094_Y), .A(D12511_Y));
KC_OR2_X2 D1798 ( .Y(D1798_Y), .B(D16696_Y), .A(D6558_Y));
KC_OR2_X2 D1659 ( .Y(D1659_Y), .B(D5489_Y), .A(D5486_Y));
KC_OR2_X2 D1657 ( .Y(D1657_Y), .B(D6197_Y), .A(D1656_Y));
KC_OR2_X2 D1387 ( .Y(D1387_Y), .B(D16772_Y), .A(D16683_Y));
KC_OR2_X2 D156 ( .Y(D156_Y), .B(D6128_Y), .A(D6074_Y));
KC_DFFRNHQ_X1 D16684 ( .Q(D16684_Q), .D(D16680_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D16682 ( .Q(D16682_Q), .D(D16678_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D16681 ( .Q(D16681_Q), .D(D16679_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D16677 ( .Q(D16677_Q), .D(D16675_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D16660 ( .Q(D16660_Q), .D(D16651_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D16650 ( .Q(D16650_Q), .D(D16648_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D16613 ( .Q(D16613_Q), .D(D16602_Y), .RN(D16579_Y),     .CK(D16581_Y));
KC_DFFRNHQ_X1 D16611 ( .Q(D16611_Q), .D(D16606_Y), .RN(D16579_Y),     .CK(D16581_Y));
KC_DFFRNHQ_X1 D16599 ( .Q(D16599_Q), .D(D16627_Y), .RN(D16579_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D16598 ( .Q(D16598_Q), .D(D16601_Y), .RN(D16579_Y),     .CK(D16581_Y));
KC_DFFRNHQ_X1 D16590 ( .Q(D16590_Q), .D(D16569_Y), .RN(D16579_Y),     .CK(D16581_Y));
KC_DFFRNHQ_X1 D16564 ( .Q(D16564_Q), .D(D16562_Y), .RN(D16579_Y),     .CK(D16581_Y));
KC_DFFRNHQ_X1 D16558 ( .Q(D16558_Q), .D(D16520_Y), .RN(D16579_Y),     .CK(D16515_QN));
KC_DFFRNHQ_X1 D16557 ( .Q(D16557_Q), .D(D16522_Y), .RN(D16579_Y),     .CK(D16515_QN));
KC_DFFRNHQ_X1 D16556 ( .Q(D16556_Q), .D(D16516_Y), .RN(D16579_Y),     .CK(D16515_QN));
KC_DFFRNHQ_X1 D16555 ( .Q(D16555_Q), .D(D16532_Y), .RN(D16376_Y),     .CK(D16455_Y));
KC_DFFRNHQ_X1 D16475 ( .Q(D16475_Q), .D(D16526_Y), .RN(D16376_Y),     .CK(D16515_QN));
KC_DFFRNHQ_X1 D16474 ( .Q(D16474_Q), .D(D16486_Y), .RN(D16377_Y),     .CK(D16455_Y));
KC_DFFRNHQ_X1 D16473 ( .Q(D16473_Q), .D(D16465_Y), .RN(D16377_Y),     .CK(D16476_Y));
KC_DFFRNHQ_X1 D16472 ( .Q(D16472_Q), .D(D16480_Y), .RN(D16377_Y),     .CK(D16455_Y));
KC_DFFRNHQ_X1 D16471 ( .Q(D16471_Q), .D(D16445_Y), .RN(D16377_Y),     .CK(D16476_Y));
KC_DFFRNHQ_X1 D16470 ( .Q(D16470_Q), .D(D16468_Y), .RN(D16377_Y),     .CK(D16476_Y));
KC_DFFRNHQ_X1 D16459 ( .Q(D16459_Q), .D(D16406_Y), .RN(D16376_Y),     .CK(D16476_Y));
KC_DFFRNHQ_X1 D16393 ( .Q(D16393_Q), .D(D16351_Y), .RN(D965_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16392 ( .Q(D16392_Q), .D(D16309_Y), .RN(D16384_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16391 ( .Q(D16391_Q), .D(D16309_Y), .RN(D16384_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D16390 ( .Q(D16390_Q), .D(D16309_Y), .RN(D16384_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D16389 ( .Q(D16389_Q), .D(D16309_Y), .RN(D16384_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D16388 ( .Q(D16388_Q), .D(D15925_Y), .RN(D16384_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D16387 ( .Q(D16387_Q), .D(D16307_Y), .RN(D16376_Y),     .CK(D16455_Y));
KC_DFFRNHQ_X1 D16386 ( .Q(D16386_Q), .D(D16373_Y), .RN(D16376_Y),     .CK(D15663_Y));
KC_DFFRNHQ_X1 D16385 ( .Q(D16385_Q), .D(D15927_Y), .RN(D16384_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16369 ( .Q(D16369_Q), .D(D15586_Y), .RN(D16352_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D16365 ( .Q(D16365_Q), .D(D16351_Y), .RN(D16352_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D16364 ( .Q(D16364_Q), .D(D16351_Y), .RN(D16352_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D16363 ( .Q(D16363_Q), .D(D2625_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D16362 ( .Q(D16362_Q), .D(D15592_Y), .RN(D2627_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D16361 ( .Q(D16361_Q), .D(D16278_Y), .RN(D2627_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D16360 ( .Q(D16360_Q), .D(D16278_Y), .RN(D2627_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16359 ( .Q(D16359_Q), .D(D16278_Y), .RN(D2627_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D16358 ( .Q(D16358_Q), .D(D15586_Y), .RN(D16352_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D16357 ( .Q(D16357_Q), .D(D1106_Y), .RN(D16352_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D16356 ( .Q(D16356_Q), .D(D15688_Y), .RN(D16352_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16355 ( .Q(D16355_Q), .D(D15586_Y), .RN(D16352_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16354 ( .Q(D16354_Q), .D(D15586_Y), .RN(D2627_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D16353 ( .Q(D16353_Q), .D(D16278_Y), .RN(D2627_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D16346 ( .Q(D16346_Q), .D(D15748_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D16340 ( .Q(D16340_Q), .D(D15587_Y), .RN(D2677_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D16319 ( .Q(D16319_Q), .D(D2666_Y), .RN(D2627_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16318 ( .Q(D16318_Q), .D(D15592_Y), .RN(D2677_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D16317 ( .Q(D16317_Q), .D(D14904_Y), .RN(D2677_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D16316 ( .Q(D16316_Q), .D(D15592_Y), .RN(D2627_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D16315 ( .Q(D16315_Q), .D(D15592_Y), .RN(D2627_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D16314 ( .Q(D16314_Q), .D(D14904_Y), .RN(D2627_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D16293 ( .Q(D16293_Q), .D(D16262_Y), .RN(D16383_Y),     .CK(D2513_QN));
KC_DFFRNHQ_X1 D16292 ( .Q(D16292_Q), .D(D16284_Y), .RN(D16383_Y),     .CK(D2513_QN));
KC_DFFRNHQ_X1 D16291 ( .Q(D16291_Q), .D(D16282_Y), .RN(D16383_Y),     .CK(D2513_QN));
KC_DFFRNHQ_X1 D16290 ( .Q(D16290_Q), .D(D16248_Y), .RN(D16383_Y),     .CK(D2513_QN));
KC_DFFRNHQ_X1 D16289 ( .Q(D16289_Q), .D(D16254_Y), .RN(D16383_Y),     .CK(D2513_QN));
KC_DFFRNHQ_X1 D16288 ( .Q(D16288_Q), .D(D16296_Y), .RN(D16383_Y),     .CK(D2586_Y));
KC_DFFRNHQ_X1 D16287 ( .Q(D16287_Q), .D(D2656_Y), .RN(D16383_Y),     .CK(D2586_Y));
KC_DFFRNHQ_X1 D16242 ( .Q(D16242_Q), .D(D16204_Y), .RN(D16383_Y),     .CK(D2568_Y));
KC_DFFRNHQ_X1 D16225 ( .Q(D16225_Q), .D(D16138_Y), .RN(D15652_Y),     .CK(D2568_Y));
KC_DFFRNHQ_X1 D16014 ( .Q(D16014_Q), .D(D15789_Y), .RN(D15990_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D16013 ( .Q(D16013_Q), .D(D877_Y), .RN(D15990_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D16012 ( .Q(D16012_Q), .D(D15684_Y), .RN(D15990_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D16011 ( .Q(D16011_Q), .D(D15684_Y), .RN(D15990_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D16010 ( .Q(D16010_Q), .D(D15974_Y), .RN(D15990_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D16009 ( .Q(D16009_Q), .D(D15684_Y), .RN(D15990_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D16008 ( .Q(D16008_Q), .D(D15684_Y), .RN(D15990_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D15999 ( .Q(D15999_Q), .D(D877_Y), .RN(D16383_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D15998 ( .Q(D15998_Q), .D(D15927_Y), .RN(D16384_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D15997 ( .Q(D15997_Q), .D(D877_Y), .RN(D15990_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D15996 ( .Q(D15996_Q), .D(D15927_Y), .RN(D16384_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D15995 ( .Q(D15995_Q), .D(D16381_Y), .RN(D16384_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D15994 ( .Q(D15994_Q), .D(D15981_Y), .RN(D16383_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D15993 ( .Q(D15993_Q), .D(D877_Y), .RN(D15990_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D15992 ( .Q(D15992_Q), .D(D15973_Y), .RN(D15990_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15991 ( .Q(D15991_Q), .D(D16002_Y), .RN(D15990_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15949 ( .Q(D15949_Q), .D(D15918_Y), .RN(D16384_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D15948 ( .Q(D15948_Q), .D(D15926_Y), .RN(D16352_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D15947 ( .Q(D15947_Q), .D(D15921_Y), .RN(D16384_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D15874 ( .Q(D15874_Q), .D(D2621_Y), .RN(D14296_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15873 ( .Q(D15873_Q), .D(D2620_Y), .RN(D16352_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15872 ( .Q(D15872_Q), .D(D15688_Y), .RN(D16352_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D15871 ( .Q(D15871_Q), .D(D15688_Y), .RN(D16352_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D15870 ( .Q(D15870_Q), .D(D15836_Y), .RN(D16352_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D15869 ( .Q(D15869_Q), .D(D15837_Y), .RN(D16352_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D15868 ( .Q(D15868_Q), .D(D15847_Y), .RN(D16352_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15797 ( .Q(D15797_Q), .D(D2666_Y), .RN(D2677_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D15796 ( .Q(D15796_Q), .D(D15762_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15795 ( .Q(D15795_Q), .D(D15764_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15794 ( .Q(D15794_Q), .D(D14904_Y), .RN(D2677_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D15793 ( .Q(D15793_Q), .D(D15746_Y), .RN(D15790_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15792 ( .Q(D15792_Q), .D(D15755_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15791 ( .Q(D15791_Q), .D(D15754_Y), .RN(D15790_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D15711 ( .Q(D15711_Q), .D(D15664_Y), .RN(D15790_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D15670 ( .Q(D15670_Q), .D(D15587_Y), .RN(D15790_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D15669 ( .Q(D15669_Q), .D(D15664_Y), .RN(D2677_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D15668 ( .Q(D15668_Q), .D(D15770_Y), .RN(D15790_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D15238 ( .Q(D15238_Q), .D(D15838_Y), .RN(D15990_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D15237 ( .Q(D15237_Q), .D(D15128_Y), .RN(D15990_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D15236 ( .Q(D15236_Q), .D(D15838_Y), .RN(D15990_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D15235 ( .Q(D15235_Q), .D(D15789_Y), .RN(D15990_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D15234 ( .Q(D15234_Q), .D(D15838_Y), .RN(D14489_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D15233 ( .Q(D15233_Q), .D(D15128_Y), .RN(D14489_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D15232 ( .Q(D15232_Q), .D(D15183_Y), .RN(D14489_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15231 ( .Q(D15231_Q), .D(D15128_Y), .RN(D15990_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D15230 ( .Q(D15230_Q), .D(D15789_Y), .RN(D14489_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D15229 ( .Q(D15229_Q), .D(D15184_Y), .RN(D14489_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15218 ( .Q(D15218_Q), .D(D2549_Y), .RN(D14291_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15217 ( .Q(D15217_Q), .D(D15195_Y), .RN(D14291_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15216 ( .Q(D15216_Q), .D(D15210_Y), .RN(D14489_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15215 ( .Q(D15215_Q), .D(D15202_Y), .RN(D14291_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15214 ( .Q(D15214_Q), .D(D15191_Y), .RN(D14489_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15213 ( .Q(D15213_Q), .D(D15209_Y), .RN(D14291_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15212 ( .Q(D15212_Q), .D(D15198_Y), .RN(D14291_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D15134 ( .Q(D15134_Q), .D(D15116_Y), .RN(D14291_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D15133 ( .Q(D15133_Q), .D(D15920_Y), .RN(D14291_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D15084 ( .Q(D15084_Q), .D(D15049_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D14997 ( .Q(D14997_Q), .D(D15664_Y), .RN(D14869_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14996 ( .Q(D14996_Q), .D(D14966_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D14995 ( .Q(D14995_Q), .D(D14967_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D14903 ( .Q(D14903_Q), .D(D2556_Y), .RN(D15790_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D14878 ( .Q(D14878_Q), .D(D2561_Y), .RN(D15790_Y),     .CK(D14162_QN));
KC_DFFRNHQ_X1 D14877 ( .Q(D14877_Q), .D(D2562_Y), .RN(D15790_Y),     .CK(D14162_QN));
KC_DFFRNHQ_X1 D14876 ( .Q(D14876_Q), .D(D14761_Y), .RN(D15790_Y),     .CK(D14162_QN));
KC_DFFRNHQ_X1 D14875 ( .Q(D14875_Q), .D(D2557_Y), .RN(D15790_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D14874 ( .Q(D14874_Q), .D(D15683_Y), .RN(D15790_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14873 ( .Q(D14873_Q), .D(D14855_Y), .RN(D15790_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D14872 ( .Q(D14872_Q), .D(D14904_Y), .RN(D15790_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D14871 ( .Q(D14871_Q), .D(D2626_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D14870 ( .Q(D14870_Q), .D(D15664_Y), .RN(D14869_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D14815 ( .Q(D14815_Q), .D(D14755_Y), .RN(D15790_Y),     .CK(D14112_QN));
KC_DFFRNHQ_X1 D14814 ( .Q(D14814_Q), .D(D14757_Y), .RN(D15790_Y),     .CK(D14112_QN));
KC_DFFRNHQ_X1 D14808 ( .Q(D14808_Q), .D(D14765_Y), .RN(D14474_Y),     .CK(D13261_QN));
KC_DFFRNHQ_X1 D14790 ( .Q(D14790_Q), .D(D14770_Y), .RN(D13265_Y),     .CK(D14080_QN));
KC_DFFRNHQ_X1 D14789 ( .Q(D14789_Q), .D(D14768_Y), .RN(D13265_Y),     .CK(D14080_QN));
KC_DFFRNHQ_X1 D14788 ( .Q(D14788_Q), .D(D14764_Y), .RN(D14474_Y),     .CK(D13261_QN));
KC_DFFRNHQ_X1 D14787 ( .Q(D14787_Q), .D(D14756_Y), .RN(D15790_Y),     .CK(D14112_QN));
KC_DFFRNHQ_X1 D14689 ( .Q(D14689_Q), .D(D14659_Y), .RN(D13265_Y),     .CK(D13263_QN));
KC_DFFRNHQ_X1 D14688 ( .Q(D14688_Q), .D(D14636_Y), .RN(D13265_Y),     .CK(D15663_Y));
KC_DFFRNHQ_X1 D14687 ( .Q(D14687_Q), .D(D14709_Y), .RN(D13265_Y),     .CK(D15663_Y));
KC_DFFRNHQ_X1 D14686 ( .Q(D14686_Q), .D(D14617_Y), .RN(D13265_Y),     .CK(D13263_QN));
KC_DFFRNHQ_X1 D14685 ( .Q(D14685_Q), .D(D14658_Y), .RN(D13265_Y),     .CK(D13263_QN));
KC_DFFRNHQ_X1 D14601 ( .Q(D14601_Q), .D(D14561_Y), .RN(D13185_Y),     .CK(D14579_Y));
KC_DFFRNHQ_X1 D14520 ( .Q(D14520_Q), .D(D14565_Y), .RN(D13185_Y),     .CK(D14579_Y));
KC_DFFRNHQ_X1 D14519 ( .Q(D14519_Q), .D(D14559_Y), .RN(D13185_Y),     .CK(D14579_Y));
KC_DFFRNHQ_X1 D14518 ( .Q(D14518_Q), .D(D14600_Y), .RN(D13185_Y),     .CK(D14579_Y));
KC_DFFRNHQ_X1 D14496 ( .Q(D14496_Q), .D(D14760_Y), .RN(D14489_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D14495 ( .Q(D14495_Q), .D(D15113_Y), .RN(D14489_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D14494 ( .Q(D14494_Q), .D(D14856_Y), .RN(D14489_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D14493 ( .Q(D14493_Q), .D(D14760_Y), .RN(D14489_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D14492 ( .Q(D14492_Q), .D(D15113_Y), .RN(D14489_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D14491 ( .Q(D14491_Q), .D(D15648_Y), .RN(D14489_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D14490 ( .Q(D14490_Q), .D(D14456_Y), .RN(D14474_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D14475 ( .Q(D14475_Q), .D(D14458_Y), .RN(D14474_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D14375 ( .Q(D14375_Q), .D(D14368_Y), .RN(D14288_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D14374 ( .Q(D14374_Q), .D(D14367_Y), .RN(D14288_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D14316 ( .Q(D14316_Q), .D(D15691_Y), .RN(D14288_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14308 ( .Q(D14308_Q), .D(D15691_Y), .RN(D14288_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14307 ( .Q(D14307_Q), .D(D14786_Y), .RN(D14296_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D14306 ( .Q(D14306_Q), .D(D14859_Y), .RN(D14296_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14305 ( .Q(D14305_Q), .D(D14859_Y), .RN(D14288_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D14304 ( .Q(D14304_Q), .D(D2676_Y), .RN(D14296_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14303 ( .Q(D14303_Q), .D(D14786_Y), .RN(D14288_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D14302 ( .Q(D14302_Q), .D(D14859_Y), .RN(D14288_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14301 ( .Q(D14301_Q), .D(D15691_Y), .RN(D14288_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D14300 ( .Q(D14300_Q), .D(D15058_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D14299 ( .Q(D14299_Q), .D(D15691_Y), .RN(D14288_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D14298 ( .Q(D14298_Q), .D(D762_Y), .RN(D14288_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14297 ( .Q(D14297_Q), .D(D762_Y), .RN(D14288_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14266 ( .Q(D14266_Q), .D(D998_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D14265 ( .Q(D14265_Q), .D(D15774_Y), .RN(D14869_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D14264 ( .Q(D14264_Q), .D(D15765_Y), .RN(D14474_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D14263 ( .Q(D14263_Q), .D(D994_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D14246 ( .Q(D14246_Q), .D(D15583_Y), .RN(D14474_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14245 ( .Q(D14245_Q), .D(D15774_Y), .RN(D14869_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14244 ( .Q(D14244_Q), .D(D15765_Y), .RN(D14869_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14243 ( .Q(D14243_Q), .D(D15774_Y), .RN(D14869_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14242 ( .Q(D14242_Q), .D(D15765_Y), .RN(D14869_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14241 ( .Q(D14241_Q), .D(D15694_Y), .RN(D14869_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D14240 ( .Q(D14240_Q), .D(D14786_Y), .RN(D14296_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14239 ( .Q(D14239_Q), .D(D15694_Y), .RN(D14474_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D14238 ( .Q(D14238_Q), .D(D13583_Y), .RN(D14474_Y),     .CK(D13511_Y));
KC_DFFRNHQ_X1 D14237 ( .Q(D14237_Q), .D(D14859_Y), .RN(D14296_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D14236 ( .Q(D14236_Q), .D(D15774_Y), .RN(D14869_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D14196 ( .Q(D14196_Q), .D(D15583_Y), .RN(D14474_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D14170 ( .Q(D14170_Q), .D(D14150_Y), .RN(D14163_Y),     .CK(D14162_QN));
KC_DFFRNHQ_X1 D14169 ( .Q(D14169_Q), .D(D14153_Y), .RN(D14163_Y),     .CK(D14162_QN));
KC_DFFRNHQ_X1 D14168 ( .Q(D14168_Q), .D(D14151_Y), .RN(D14163_Y),     .CK(D14162_QN));
KC_DFFRNHQ_X1 D14167 ( .Q(D14167_Q), .D(D15583_Y), .RN(D14163_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14166 ( .Q(D14166_Q), .D(D15694_Y), .RN(D14163_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D14165 ( .Q(D14165_Q), .D(D13494_Y), .RN(D2510_Y),     .CK(D13511_Y));
KC_DFFRNHQ_X1 D14164 ( .Q(D14164_Q), .D(D15694_Y), .RN(D14474_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D14118 ( .Q(D14118_Q), .D(D14048_Y), .RN(D14163_Y),     .CK(D14112_QN));
KC_DFFRNHQ_X1 D14117 ( .Q(D14117_Q), .D(D14152_Y), .RN(D14163_Y),     .CK(D14112_QN));
KC_DFFRNHQ_X1 D14109 ( .Q(D14109_Q), .D(D14055_Y), .RN(D14163_Y),     .CK(D14080_QN));
KC_DFFRNHQ_X1 D14094 ( .Q(D14094_Q), .D(D14052_Y), .RN(D13265_Y),     .CK(D14080_QN));
KC_DFFRNHQ_X1 D14093 ( .Q(D14093_Q), .D(D14056_Y), .RN(D14163_Y),     .CK(D13261_QN));
KC_DFFRNHQ_X1 D14092 ( .Q(D14092_Q), .D(D14053_Y), .RN(D14163_Y),     .CK(D14080_QN));
KC_DFFRNHQ_X1 D14091 ( .Q(D14091_Q), .D(D14049_Y), .RN(D14163_Y),     .CK(D14112_QN));
KC_DFFRNHQ_X1 D13998 ( .Q(D13998_Q), .D(D14069_Y), .RN(D13242_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D13997 ( .Q(D13997_Q), .D(D14078_Y), .RN(D13266_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13996 ( .Q(D13996_Q), .D(D14075_Y), .RN(D13265_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13995 ( .Q(D13995_Q), .D(D14612_Y), .RN(D13265_Y),     .CK(D13263_QN));
KC_DFFRNHQ_X1 D13994 ( .Q(D13994_Q), .D(D14069_Y), .RN(D13242_Y),     .CK(D13214_QN));
KC_DFFRNHQ_X1 D13993 ( .Q(D13993_Q), .D(D14069_Y), .RN(D13265_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13992 ( .Q(D13992_Q), .D(D14075_Y), .RN(D13242_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13991 ( .Q(D13991_Q), .D(D14078_Y), .RN(D13266_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13990 ( .Q(D13990_Q), .D(D14069_Y), .RN(D13242_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13989 ( .Q(D13989_Q), .D(D14075_Y), .RN(D13266_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D13921 ( .Q(D13921_Q), .D(D12741_Y), .RN(D13194_Y),     .CK(D13193_QN));
KC_DFFRNHQ_X1 D13920 ( .Q(D13920_Q), .D(D12741_Y), .RN(D13194_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13918 ( .Q(D13918_Q), .D(D12666_Y), .RN(D13194_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13909 ( .Q(D13909_Q), .D(D12672_Y), .RN(D13194_Y),     .CK(D13193_QN));
KC_DFFRNHQ_X1 D13908 ( .Q(D13908_Q), .D(D12671_Y), .RN(D13265_Y),     .CK(D13193_QN));
KC_DFFRNHQ_X1 D13907 ( .Q(D13907_Q), .D(D12666_Y), .RN(D13194_Y),     .CK(D13193_QN));
KC_DFFRNHQ_X1 D13872 ( .Q(D13872_Q), .D(D13851_Y), .RN(D13185_Y),     .CK(D506_QN));
KC_DFFRNHQ_X1 D13865 ( .Q(D13865_Q), .D(D13850_Y), .RN(D13185_Y),     .CK(D506_QN));
KC_DFFRNHQ_X1 D13864 ( .Q(D13864_Q), .D(D13853_Y), .RN(D13185_Y),     .CK(D506_QN));
KC_DFFRNHQ_X1 D13860 ( .Q(D13860_Q), .D(D12673_Y), .RN(D13194_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13827 ( .Q(D13827_Q), .D(D2500_Y), .RN(D13825_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D13826 ( .Q(D13826_Q), .D(D14856_Y), .RN(D14474_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D13816 ( .Q(D13816_Q), .D(D13785_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13815 ( .Q(D13815_Q), .D(D2439_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13814 ( .Q(D13814_Q), .D(D1283_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13813 ( .Q(D13813_Q), .D(D15648_Y), .RN(D13825_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D13812 ( .Q(D13812_Q), .D(D2500_Y), .RN(D13825_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D13811 ( .Q(D13811_Q), .D(D13782_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13810 ( .Q(D13810_Q), .D(D15648_Y), .RN(D13825_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D13809 ( .Q(D13809_Q), .D(D13790_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13808 ( .Q(D13808_Q), .D(D14856_Y), .RN(D13825_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D13807 ( .Q(D13807_Q), .D(D13791_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13806 ( .Q(D13806_Q), .D(D15648_Y), .RN(D13825_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D13805 ( .Q(D13805_Q), .D(D2500_Y), .RN(D13825_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D13804 ( .Q(D13804_Q), .D(D13788_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13771 ( .Q(D13771_Q), .D(D13733_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13770 ( .Q(D13770_Q), .D(D762_Y), .RN(D13758_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D13765 ( .Q(D13765_Q), .D(D13742_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D13764 ( .Q(D13764_Q), .D(D13743_Y), .RN(D13758_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13762 ( .Q(D13762_Q), .D(D13735_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13761 ( .Q(D13761_Q), .D(D13737_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13760 ( .Q(D13760_Q), .D(D13731_Y), .RN(D13825_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D13759 ( .Q(D13759_Q), .D(D14856_Y), .RN(D13825_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D13711 ( .Q(D13711_Q), .D(D13687_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D13706 ( .Q(D13706_Q), .D(D13686_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D13705 ( .Q(D13705_Q), .D(D13685_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D13704 ( .Q(D13704_Q), .D(D13683_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D13703 ( .Q(D13703_Q), .D(D2440_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D13530 ( .Q(D13530_Q), .D(D13500_Y), .RN(D12901_Y),     .CK(D13511_Y));
KC_DFFRNHQ_X1 D13515 ( .Q(D13515_Q), .D(D2450_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D13398 ( .Q(D13398_Q), .D(D13233_Y), .RN(D13242_Y),     .CK(D13264_QN));
KC_DFFRNHQ_X1 D13397 ( .Q(D13397_Q), .D(D13351_Y), .RN(D13242_Y),     .CK(D13264_QN));
KC_DFFRNHQ_X1 D13396 ( .Q(D13396_Q), .D(D13341_Y), .RN(D13242_Y),     .CK(D13264_QN));
KC_DFFRNHQ_X1 D13395 ( .Q(D13395_Q), .D(D13371_Y), .RN(D13242_Y),     .CK(D13264_QN));
KC_DFFRNHQ_X1 D13279 ( .Q(D13279_Q), .D(D13250_Y), .RN(D13266_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D13275 ( .Q(D13275_Q), .D(D13386_Y), .RN(D13266_Y),     .CK(D2460_Y));
KC_DFFRNHQ_X1 D13274 ( .Q(D13274_Q), .D(D13244_Y), .RN(D13266_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X1 D13273 ( .Q(D13273_Q), .D(D13250_Y), .RN(D13242_Y),     .CK(D2460_Y));
KC_DFFRNHQ_X1 D13272 ( .Q(D13272_Q), .D(D13386_Y), .RN(D13266_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D13271 ( .Q(D13271_Q), .D(D13386_Y), .RN(D13266_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13270 ( .Q(D13270_Q), .D(D13232_Y), .RN(D13266_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X1 D13269 ( .Q(D13269_Q), .D(D627_Y), .RN(D13242_Y),     .CK(D13264_QN));
KC_DFFRNHQ_X1 D13268 ( .Q(D13268_Q), .D(D12723_Y), .RN(D13242_Y),     .CK(D12746_QN));
KC_DFFRNHQ_X1 D13267 ( .Q(D13267_Q), .D(D632_Y), .RN(D13242_Y),     .CK(D13264_QN));
KC_DFFRNHQ_X1 D13195 ( .Q(D13195_Q), .D(D13179_Y), .RN(D12679_Y),     .CK(D13193_QN));
KC_DFFRNHQ_X1 D13216 ( .Q(D13216_Q), .D(D13399_Y), .RN(D13266_Y),     .CK(D13214_QN));
KC_DFFRNHQ_X1 D13213 ( .Q(D13213_Q), .D(D13278_Y), .RN(D12679_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X1 D13212 ( .Q(D13212_Q), .D(D13384_Y), .RN(D13266_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13211 ( .Q(D13211_Q), .D(D12671_Y), .RN(D12679_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13210 ( .Q(D13210_Q), .D(D12665_Y), .RN(D12679_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13209 ( .Q(D13209_Q), .D(D12741_Y), .RN(D13194_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13208 ( .Q(D13208_Q), .D(D14079_Y), .RN(D13194_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13203 ( .Q(D13203_Q), .D(D12672_Y), .RN(D12679_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13202 ( .Q(D13202_Q), .D(D13384_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D13201 ( .Q(D13201_Q), .D(D12671_Y), .RN(D13194_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13200 ( .Q(D13200_Q), .D(D12671_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D13199 ( .Q(D13199_Q), .D(D13384_Y), .RN(D12679_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D13198 ( .Q(D13198_Q), .D(D13384_Y), .RN(D13266_Y),     .CK(D2460_Y));
KC_DFFRNHQ_X1 D13197 ( .Q(D13197_Q), .D(D14079_Y), .RN(D13194_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D13196 ( .Q(D13196_Q), .D(D13399_Y), .RN(D13266_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D13175 ( .Q(D13175_Q), .D(D500_Y), .RN(D13185_Y),     .CK(D506_QN));
KC_DFFRNHQ_X1 D13051 ( .Q(D13051_Q), .D(D13025_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D13050 ( .Q(D13050_Q), .D(D13026_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D12997 ( .Q(D12997_Q), .D(D12959_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12996 ( .Q(D12996_Q), .D(D13638_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12995 ( .Q(D12995_Q), .D(D12954_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12994 ( .Q(D12994_Q), .D(D13594_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12993 ( .Q(D12993_Q), .D(D13589_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12992 ( .Q(D12992_Q), .D(D13593_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12991 ( .Q(D12991_Q), .D(D12948_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12936 ( .Q(D12936_Q), .D(D12883_Y), .RN(D12900_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12935 ( .Q(D12935_Q), .D(D12890_Y), .RN(D12900_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D12934 ( .Q(D12934_Q), .D(D12832_Y), .RN(D12900_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D12926 ( .Q(D12926_Q), .D(D2452_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D12925 ( .Q(D12925_Q), .D(D12891_Y), .RN(D12846_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12924 ( .Q(D12924_Q), .D(D12885_Y), .RN(D12900_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12923 ( .Q(D12923_Q), .D(D12884_Y), .RN(D12900_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12922 ( .Q(D12922_Q), .D(D12906_Y), .RN(D12900_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D12921 ( .Q(D12921_Q), .D(D13483_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12920 ( .Q(D12920_Q), .D(D12832_Y), .RN(D12900_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D12919 ( .Q(D12919_Q), .D(D13418_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12918 ( .Q(D12918_Q), .D(D13480_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D12917 ( .Q(D12917_Q), .D(D12882_Y), .RN(D12846_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12916 ( .Q(D12916_Q), .D(D12868_Y), .RN(D12900_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D12915 ( .Q(D12915_Q), .D(D12906_Y), .RN(D12846_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D12914 ( .Q(D12914_Q), .D(D12906_Y), .RN(D12900_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D12858 ( .Q(D12858_Q), .D(D12839_Y), .RN(D12846_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D12857 ( .Q(D12857_Q), .D(D12817_Y), .RN(D12846_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D12856 ( .Q(D12856_Q), .D(D12840_Y), .RN(D12846_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X1 D12855 ( .Q(D12855_Q), .D(D12828_Y), .RN(D12846_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D12854 ( .Q(D12854_Q), .D(D12822_Y), .RN(D12846_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12853 ( .Q(D12853_Q), .D(D12812_Y), .RN(D12846_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12852 ( .Q(D12852_Q), .D(D12811_Y), .RN(D12846_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12851 ( .Q(D12851_Q), .D(D12832_Y), .RN(D12846_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D12850 ( .Q(D12850_Q), .D(D2378_Y), .RN(D12846_Y),     .CK(D12903_Y));
KC_DFFRNHQ_X1 D12849 ( .Q(D12849_Q), .D(D12890_Y), .RN(D12846_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D12848 ( .Q(D12848_Q), .D(D12832_Y), .RN(D12846_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D12756 ( .Q(D12756_Q), .D(D12721_Y), .RN(D12258_Y),     .CK(D12746_QN));
KC_DFFRNHQ_X1 D12755 ( .Q(D12755_Q), .D(D12724_Y), .RN(D12258_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D12754 ( .Q(D12754_Q), .D(D12709_Y), .RN(D12258_Y),     .CK(D12746_QN));
KC_DFFRNHQ_X1 D12753 ( .Q(D12753_Q), .D(D13223_Y), .RN(D12258_Y),     .CK(D12746_QN));
KC_DFFRNHQ_X1 D12752 ( .Q(D12752_Q), .D(D12727_Y), .RN(D12258_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D12749 ( .Q(D12749_Q), .D(D12818_Y), .RN(D12258_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D12748 ( .Q(D12748_Q), .D(D12802_Y), .RN(D12258_Y),     .CK(D12740_Y));
KC_DFFRNHQ_X1 D12689 ( .Q(D12689_Q), .D(D12673_Y), .RN(D12679_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D12688 ( .Q(D12688_Q), .D(D12666_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D12687 ( .Q(D12687_Q), .D(D2365_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D12686 ( .Q(D12686_Q), .D(D12741_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D12685 ( .Q(D12685_Q), .D(D13179_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D12684 ( .Q(D12684_Q), .D(D12665_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D12683 ( .Q(D12683_Q), .D(D13179_Y), .RN(D12662_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D12682 ( .Q(D12682_Q), .D(D12673_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D12681 ( .Q(D12681_Q), .D(D12672_Y), .RN(D12679_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D12680 ( .Q(D12680_Q), .D(D12666_Y), .RN(D12679_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D12419 ( .Q(D12419_Q), .D(D12393_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12418 ( .Q(D12418_Q), .D(D12394_Y), .RN(D12900_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12417 ( .Q(D12417_Q), .D(D2335_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12416 ( .Q(D12416_Q), .D(D2333_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12415 ( .Q(D12415_Q), .D(D12395_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12414 ( .Q(D12414_Q), .D(D12396_Y), .RN(D12900_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12368 ( .Q(D12368_Q), .D(D12322_Y), .RN(D10725_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D12367 ( .Q(D12367_Q), .D(D12330_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12360 ( .Q(D12360_Q), .D(D12326_Y), .RN(D10725_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D12359 ( .Q(D12359_Q), .D(D12317_Y), .RN(D12339_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D12358 ( .Q(D12358_Q), .D(D12322_Y), .RN(D12339_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D12357 ( .Q(D12357_Q), .D(D12326_Y), .RN(D10725_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D12356 ( .Q(D12356_Q), .D(D12326_Y), .RN(D10725_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D12355 ( .Q(D12355_Q), .D(D12806_Y), .RN(D12258_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D12353 ( .Q(D12353_Q), .D(D12322_Y), .RN(D12339_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D12352 ( .Q(D12352_Q), .D(D12317_Y), .RN(D12339_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D12351 ( .Q(D12351_Q), .D(D12328_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12350 ( .Q(D12350_Q), .D(D12317_Y), .RN(D12339_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D12349 ( .Q(D12349_Q), .D(D12322_Y), .RN(D12339_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D12348 ( .Q(D12348_Q), .D(D12333_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12346 ( .Q(D12346_Q), .D(D12370_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12344 ( .Q(D12344_Q), .D(D12327_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12343 ( .Q(D12343_Q), .D(D12329_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12342 ( .Q(D12342_Q), .D(D2334_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12341 ( .Q(D12341_Q), .D(D2331_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12340 ( .Q(D12340_Q), .D(D12332_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D12279 ( .Q(D12279_Q), .D(D2307_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D12278 ( .Q(D12278_Q), .D(D2308_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D12277 ( .Q(D12277_Q), .D(D2309_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D12275 ( .Q(D12275_Q), .D(D12326_Y), .RN(D10725_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D12274 ( .Q(D12274_Q), .D(D12317_Y), .RN(D10725_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D12237 ( .Q(D12237_Q), .D(D12217_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D12236 ( .Q(D12236_Q), .D(D12220_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D12235 ( .Q(D12235_Q), .D(D12216_Y), .RN(D12662_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D12234 ( .Q(D12234_Q), .D(D12219_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D12177 ( .Q(D12177_Q), .D(D16761_Y), .RN(D12177_RN),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D11672 ( .Q(D11672_Q), .D(D141_Q), .RN(D11636_SN),     .CK(D12174_Y));
KC_DFFRNHQ_X1 D10368 ( .Q(D10368_Q), .D(D10363_Q), .RN(D9538_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10365 ( .Q(D10365_Q), .D(D2168_Q), .RN(D9538_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10364 ( .Q(D10364_Q), .D(D946_Q), .RN(D9538_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10363 ( .Q(D10363_Q), .D(D10371_Q), .RN(D9538_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10362 ( .Q(D10362_Q), .D(D10367_Y), .RN(D10325_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10361 ( .Q(D10361_Q), .D(D10322_Y), .RN(D10330_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10360 ( .Q(D10360_Q), .D(D10319_Y), .RN(D10341_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10359 ( .Q(D10359_Q), .D(D10346_Y), .RN(D10327_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D10311 ( .Q(D10311_Q), .D(D10262_Y), .RN(D9381_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10308 ( .Q(D10308_Q), .D(D10732_Y), .RN(D10369_Y),     .CK(D10746_Y));
KC_DFFRNHQ_X1 D10307 ( .Q(D10307_Q), .D(D10313_Y), .RN(D10285_Y),     .CK(D10821_Y));
KC_DFFRNHQ_X1 D10306 ( .Q(D10306_Q), .D(D10746_Y), .RN(D10369_Y),     .CK(D10735_Y));
KC_DFFRNHQ_X1 D10305 ( .Q(D10305_Q), .D(D10304_Q), .RN(D10357_Y),     .CK(D10821_Y));
KC_DFFRNHQ_X1 D10304 ( .Q(D10304_Q), .D(D10292_Y), .RN(D10369_Y),     .CK(D10732_Y));
KC_DFFRNHQ_X1 D10303 ( .Q(D10303_Q), .D(D10261_Y), .RN(D9381_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10302 ( .Q(D10302_Q), .D(D10260_Y), .RN(D9381_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10301 ( .Q(D10301_Q), .D(D10312_Y), .RN(D9381_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10300 ( .Q(D10300_Q), .D(D849_Y), .RN(D12838_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10299 ( .Q(D10299_Q), .D(D10314_Y), .RN(D10725_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10298 ( .Q(D10298_Q), .D(D10269_Y), .RN(D10357_Y),     .CK(D709_Y));
KC_DFFRNHQ_X1 D10297 ( .Q(D10297_Q), .D(D9561_Y), .RN(D9538_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D10296 ( .Q(D10296_Q), .D(D2143_Y), .RN(D10725_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10295 ( .Q(D10295_Q), .D(D10735_Y), .RN(D10369_Y),     .CK(D11632_Y));
KC_DFFRNHQ_X1 D10294 ( .Q(D10294_Q), .D(D10263_Y), .RN(D10725_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D10293 ( .Q(D10293_Q), .D(D10270_Y), .RN(D2149_Y),     .CK(D10821_Y));
KC_DFFRNHQ_X1 D10231 ( .Q(D10231_Q), .D(D10240_Co), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10229 ( .Q(D10229_Q), .D(D9943_Y), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10228 ( .Q(D10228_Q), .D(D10229_Q), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10227 ( .Q(D10227_Q), .D(D10228_Q), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10226 ( .Q(D10226_Q), .D(D8453_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D10225 ( .Q(D10225_Q), .D(D10784_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D10224 ( .Q(D10224_Q), .D(D9942_Y), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10223 ( .Q(D10223_Q), .D(D10224_Q), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10222 ( .Q(D10222_Q), .D(D9985_Y), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10221 ( .Q(D10221_Q), .D(D16759_Co), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10220 ( .Q(D10220_Q), .D(D10223_Q), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D10219 ( .Q(D10219_Q), .D(D698_Q), .RN(D10726_Y),     .CK(D10821_Y));
KC_DFFRNHQ_X1 D10218 ( .Q(D10218_Q), .D(D10217_Q), .RN(D10726_Y),     .CK(D10821_Y));
KC_DFFRNHQ_X1 D10217 ( .Q(D10217_Q), .D(D16758_Co), .RN(D10726_Y),     .CK(D10821_Y));
KC_DFFRNHQ_X1 D10147 ( .Q(D10147_Q), .D(D9176_Y), .RN(D9271_Y),     .CK(D9212_QN));
KC_DFFRNHQ_X1 D10146 ( .Q(D10146_Q), .D(D9238_Y), .RN(D9271_Y),     .CK(D10107_QN));
KC_DFFRNHQ_X1 D10145 ( .Q(D10145_Q), .D(D9238_Y), .RN(D9271_Y),     .CK(D9212_QN));
KC_DFFRNHQ_X1 D10109 ( .Q(D10109_Q), .D(D16745_Y), .RN(D9271_Y),     .CK(D9140_QN));
KC_DFFRNHQ_X1 D10108 ( .Q(D10108_Q), .D(D422_Y), .RN(D9128_Y),     .CK(D9139_QN));
KC_DFFRNHQ_X1 D10062 ( .Q(D10062_Q), .D(D1921_Y), .RN(D324_Y),     .CK(D443_QN));
KC_DFFRNHQ_X1 D10061 ( .Q(D10061_Q), .D(D9089_Y), .RN(D324_Y),     .CK(D9141_QN));
KC_DFFRNHQ_X1 D10060 ( .Q(D10060_Q), .D(D9088_Y), .RN(D324_Y),     .CK(D9141_QN));
KC_DFFRNHQ_X1 D10059 ( .Q(D10059_Q), .D(D10056_Y), .RN(D324_Y),     .CK(D443_QN));
KC_DFFRNHQ_X1 D10058 ( .Q(D10058_Q), .D(D10063_Y), .RN(D324_Y),     .CK(D443_QN));
KC_DFFRNHQ_X1 D10051 ( .Q(D10051_Q), .D(D2142_Y), .RN(D324_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10049 ( .Q(D10049_Q), .D(D10038_Y), .RN(D324_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10048 ( .Q(D10048_Q), .D(D10042_Y), .RN(D324_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10047 ( .Q(D10047_Q), .D(D10041_Y), .RN(D324_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10033 ( .Q(D10033_Q), .D(D10022_Y), .RN(D8894_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10032 ( .Q(D10032_Q), .D(D10025_Y), .RN(D324_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10031 ( .Q(D10031_Q), .D(D10023_Y), .RN(D324_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10009 ( .Q(D10009_Q), .D(D10020_Y), .RN(D8894_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10008 ( .Q(D10008_Q), .D(D10004_Y), .RN(D8818_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10007 ( .Q(D10007_Q), .D(D256_Y), .RN(D8894_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D10006 ( .Q(D10006_Q), .D(D10003_Y), .RN(D8894_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D9984 ( .Q(D9984_Q), .D(D9959_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D9983 ( .Q(D9983_Q), .D(D9994_Y), .RN(D8818_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D9982 ( .Q(D9982_Q), .D(D8884_Y), .RN(D8818_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D9981 ( .Q(D9981_Q), .D(D9987_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D9980 ( .Q(D9980_Q), .D(D9969_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D9950 ( .Q(D9950_Q), .D(D9930_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D9941 ( .Q(D9941_Q), .D(D9929_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D9625 ( .Q(D9625_Q), .D(D9624_Q), .RN(D10357_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D9624 ( .Q(D9624_Q), .D(D2072_Y), .RN(D10357_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D9623 ( .Q(D9623_Q), .D(D9635_Q), .RN(D10357_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D9622 ( .Q(D9622_Q), .D(D9629_Q), .RN(D10357_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D9621 ( .Q(D9621_Q), .D(D9636_Y), .RN(D10357_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D9620 ( .Q(D9620_Q), .D(D947_Q), .RN(D10357_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D9582 ( .Q(D9582_Q), .D(D9471_Q), .RN(D9381_Y),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D9581 ( .Q(D9581_Q), .D(D9433_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D9580 ( .Q(D9580_Q), .D(D10786_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D9579 ( .Q(D9579_Q), .D(D9500_Y), .RN(D12838_Y),     .CK(D775_QN));
KC_DFFRNHQ_X1 D9578 ( .Q(D9578_Q), .D(D9589_Y), .RN(D12838_Y),     .CK(D775_QN));
KC_DFFRNHQ_X1 D9577 ( .Q(D9577_Q), .D(D9537_Y), .RN(D12838_Y),     .CK(D775_QN));
KC_DFFRNHQ_X1 D9576 ( .Q(D9576_Q), .D(D9541_Y), .RN(D12838_Y),     .CK(D775_QN));
KC_DFFRNHQ_X1 D9575 ( .Q(D9575_Q), .D(D9557_Y), .RN(D12838_Y),     .CK(D775_QN));
KC_DFFRNHQ_X1 D9574 ( .Q(D9574_Q), .D(D9586_Y), .RN(D12838_Y),     .CK(D775_QN));
KC_DFFRNHQ_X1 D9472 ( .Q(D9472_Q), .D(D9435_Y), .RN(D9446_Y),     .CK(D9321_Y));
KC_DFFRNHQ_X1 D9471 ( .Q(D9471_Q), .D(D654_Y), .RN(D9381_Y),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D9470 ( .Q(D9470_Q), .D(D10203_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D9356 ( .Q(D9356_Q), .D(D9351_Y), .RN(D12302_Y),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D9355 ( .Q(D9355_Q), .D(D1995_Y), .RN(D9375_Y),     .CK(D9346_Y));
KC_DFFRNHQ_X1 D9325 ( .Q(D9325_Q), .D(D9253_Y), .RN(D7892_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D9280 ( .Q(D9280_Q), .D(D9225_Y), .RN(D9271_Y),     .CK(D7530_QN));
KC_DFFRNHQ_X1 D9279 ( .Q(D9279_Q), .D(D9262_Y), .RN(D9271_Y),     .CK(D9141_QN));
KC_DFFRNHQ_X1 D9278 ( .Q(D9278_Q), .D(D9296_Y), .RN(D7788_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D9277 ( .Q(D9277_Q), .D(D9286_Y), .RN(D9271_Y),     .CK(D7530_QN));
KC_DFFRNHQ_X1 D9276 ( .Q(D9276_Q), .D(D9261_Y), .RN(D9271_Y),     .CK(D9141_QN));
KC_DFFRNHQ_X1 D9275 ( .Q(D9275_Q), .D(D9298_Y), .RN(D7788_Y),     .CK(D416_QN));
KC_DFFRNHQ_X1 D9274 ( .Q(D9274_Q), .D(D9283_Y), .RN(D9271_Y),     .CK(D7530_QN));
KC_DFFRNHQ_X1 D9273 ( .Q(D9273_Q), .D(D9284_Y), .RN(D9271_Y),     .CK(D7530_QN));
KC_DFFRNHQ_X1 D9272 ( .Q(D9272_Q), .D(D9197_Y), .RN(D7892_Y),     .CK(D9212_QN));
KC_DFFRNHQ_X1 D9221 ( .Q(D9221_Q), .D(D9187_Y), .RN(D9128_Y),     .CK(D9142_QN));
KC_DFFRNHQ_X1 D9220 ( .Q(D9220_Q), .D(D9182_Y), .RN(D9271_Y),     .CK(D9142_QN));
KC_DFFRNHQ_X1 D9219 ( .Q(D9219_Q), .D(D9195_Y), .RN(D7788_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D9218 ( .Q(D9218_Q), .D(D424_Y), .RN(D9214_Y),     .CK(D9139_QN));
KC_DFFRNHQ_X1 D9217 ( .Q(D9217_Q), .D(D9201_Y), .RN(D9214_Y),     .CK(D9212_QN));
KC_DFFRNHQ_X1 D9216 ( .Q(D9216_Q), .D(D9192_Y), .RN(D9214_Y),     .CK(D7530_QN));
KC_DFFRNHQ_X1 D9215 ( .Q(D9215_Q), .D(D9191_Y), .RN(D9128_Y),     .CK(D9142_QN));
KC_DFFRNHQ_X1 D9150 ( .Q(D9150_Q), .D(D9137_Y), .RN(D9214_Y),     .CK(D9141_QN));
KC_DFFRNHQ_X1 D9149 ( .Q(D9149_Q), .D(D9134_Y), .RN(D9128_Y),     .CK(D9141_QN));
KC_DFFRNHQ_X1 D9148 ( .Q(D9148_Q), .D(D389_Y), .RN(D9214_Y),     .CK(D9139_QN));
KC_DFFRNHQ_X1 D9023 ( .Q(D9023_Q), .D(D313_Y), .RN(D324_Y),     .CK(D7466_QN));
KC_DFFRNHQ_X1 D9021 ( .Q(D9021_Q), .D(D319_Y), .RN(D4461_Y),     .CK(D7468_QN));
KC_DFFRNHQ_X1 D9019 ( .Q(D9019_Q), .D(D2015_Y), .RN(D324_Y),     .CK(D7466_QN));
KC_DFFRNHQ_X1 D8955 ( .Q(D8955_Q), .D(D8940_Y), .RN(D8894_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8954 ( .Q(D8954_Q), .D(D8915_Y), .RN(D8894_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8953 ( .Q(D8953_Q), .D(D8929_Y), .RN(D4461_Y),     .CK(D7468_QN));
KC_DFFRNHQ_X1 D8952 ( .Q(D8952_Q), .D(D7414_Y), .RN(D8894_Y),     .CK(D9139_QN));
KC_DFFRNHQ_X1 D8951 ( .Q(D8951_Q), .D(D2048_Y), .RN(D4461_Y),     .CK(D7468_QN));
KC_DFFRNHQ_X1 D8899 ( .Q(D8899_Q), .D(D8875_Y), .RN(D8818_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8898 ( .Q(D8898_Q), .D(D2051_Y), .RN(D8818_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8897 ( .Q(D8897_Q), .D(D2021_Y), .RN(D8818_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8896 ( .Q(D8896_Q), .D(D8862_Y), .RN(D8818_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8895 ( .Q(D8895_Q), .D(D8880_Y), .RN(D8894_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8825 ( .Q(D8825_Q), .D(D9958_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D8824 ( .Q(D8824_Q), .D(D2023_Y), .RN(D8818_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D8823 ( .Q(D8823_Q), .D(D9986_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D8822 ( .Q(D8822_Q), .D(D8759_Y), .RN(D8779_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D8821 ( .Q(D8821_Q), .D(D8834_Y), .RN(D8779_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D8712 ( .Q(D8712_Q), .D(D8680_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D8711 ( .Q(D8711_Q), .D(D2717_Y), .RN(D7795_Y),     .CK(D9140_QN));
KC_DFFRNHQ_X1 D8709 ( .Q(D8709_Q), .D(D8696_Y), .RN(D7795_Y),     .CK(D9140_QN));
KC_DFFRNHQ_X1 D8343 ( .Q(D8343_Q), .D(D9621_Q), .RN(D8300_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D8342 ( .Q(D8342_Q), .D(D8343_Q), .RN(D8300_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D8341 ( .Q(D8341_Q), .D(D896_Y), .RN(D8322_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D8250 ( .Q(D8250_Q), .D(D6647_Y), .RN(D12838_Y),     .CK(D8235_QN));
KC_DFFRNHQ_X1 D8249 ( .Q(D8249_Q), .D(D1896_Y), .RN(D12838_Y),     .CK(D8235_QN));
KC_DFFRNHQ_X1 D8248 ( .Q(D8248_Q), .D(D1841_Y), .RN(D12838_Y),     .CK(D8235_QN));
KC_DFFRNHQ_X1 D8247 ( .Q(D8247_Q), .D(D2040_Y), .RN(D12838_Y),     .CK(D8235_QN));
KC_DFFRNHQ_X1 D8246 ( .Q(D8246_Q), .D(D9427_Y), .RN(D12838_Y),     .CK(D8235_QN));
KC_DFFRNHQ_X1 D8245 ( .Q(D8245_Q), .D(D8236_Y), .RN(D8229_Y),     .CK(D9458_QN));
KC_DFFRNHQ_X1 D8244 ( .Q(D8244_Q), .D(D8191_Y), .RN(D8229_Y),     .CK(D9458_QN));
KC_DFFRNHQ_X1 D8243 ( .Q(D8243_Q), .D(D8265_Y), .RN(D8229_Y),     .CK(D9458_QN));
KC_DFFRNHQ_X1 D8151 ( .Q(D8151_Q), .D(D8143_Y), .RN(D9375_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D8150 ( .Q(D8150_Q), .D(D8101_Y), .RN(D12838_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D8149 ( .Q(D8149_Q), .D(D16774_Y), .RN(D12838_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D8148 ( .Q(D8148_Q), .D(D8133_Y), .RN(D12838_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D8147 ( .Q(D8147_Q), .D(D8131_Y), .RN(D12838_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D8058 ( .Q(D8058_Q), .D(D9341_Y), .RN(D9374_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D7973 ( .Q(D7973_Q), .D(D1967_Y), .RN(D9374_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D7896 ( .Q(D7896_Q), .D(D9309_Y), .RN(D7892_Y),     .CK(D416_QN));
KC_DFFRNHQ_X1 D7894 ( .Q(D7894_Q), .D(D9313_Y), .RN(D7892_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D7794 ( .Q(D7794_Q), .D(D7811_Y), .RN(D7788_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D7793 ( .Q(D7793_Q), .D(D7807_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D7791 ( .Q(D7791_Q), .D(D7805_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D7790 ( .Q(D7790_Q), .D(D7801_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D7789 ( .Q(D7789_Q), .D(D7802_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D7745 ( .Q(D7745_Q), .D(D7747_Y), .RN(D7788_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7737 ( .Q(D7737_Q), .D(D7719_Y), .RN(D7788_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7736 ( .Q(D7736_Q), .D(D1965_Y), .RN(D7788_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7735 ( .Q(D7735_Q), .D(D7748_Y), .RN(D7788_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7734 ( .Q(D7734_Q), .D(D7746_Y), .RN(D7788_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7733 ( .Q(D7733_Q), .D(D7699_Y), .RN(D7788_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7732 ( .Q(D7732_Q), .D(D7698_Y), .RN(D7788_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7659 ( .Q(D7659_Q), .D(D6264_Y), .RN(VDD),     .CK(D7575_Y));
KC_DFFRNHQ_X1 D7587 ( .Q(D7587_Q), .D(D7562_Y), .RN(D7521_Y),     .CK(D7575_Y));
KC_DFFRNHQ_X1 D7586 ( .Q(D7586_Q), .D(D7587_Q), .RN(D7521_Y),     .CK(D7575_Y));
KC_DFFRNHQ_X1 D7534 ( .Q(D7534_Q), .D(D7536_Y), .RN(D4461_Y),     .CK(D7530_QN));
KC_DFFRNHQ_X1 D7533 ( .Q(D7533_Q), .D(D1926_Y), .RN(D4483_Y),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D7481 ( .Q(D7481_Q), .D(D7432_Y), .RN(D8894_Y),     .CK(D7468_QN));
KC_DFFRNHQ_X1 D7480 ( .Q(D7480_Q), .D(D7440_Y), .RN(D9358_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D7479 ( .Q(D7479_Q), .D(D7448_Y), .RN(D4461_Y),     .CK(D7466_QN));
KC_DFFRNHQ_X1 D7478 ( .Q(D7478_Q), .D(D7462_Y), .RN(D4483_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D7476 ( .Q(D7476_Q), .D(D7484_Y), .RN(D9358_Y),     .CK(D7530_QN));
KC_DFFRNHQ_X1 D7475 ( .Q(D7475_Q), .D(D17_Y), .RN(D9358_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D7409 ( .Q(D7409_Q), .D(D7388_Y), .RN(D8894_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D7391 ( .Q(D7391_Q), .D(D5897_Y), .RN(D8894_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D7152 ( .Q(D7152_Q), .D(D7230_Y), .RN(D7795_Y),     .CK(D5799_Y));
KC_DFFRNHQ_X1 D7151 ( .Q(D7151_Q), .D(D7121_Y), .RN(D5683_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D7150 ( .Q(D7150_Q), .D(D7122_Y), .RN(D7795_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D7149 ( .Q(D7149_Q), .D(D7102_Y), .RN(D7795_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D7148 ( .Q(D7148_Q), .D(D7128_Y), .RN(D5683_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D7147 ( .Q(D7147_Q), .D(D7298_Y), .RN(D5683_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D7146 ( .Q(D7146_Q), .D(D7117_Y), .RN(D5683_Y),     .CK(D191_QN));
KC_DFFRNHQ_X1 D7145 ( .Q(D7145_Q), .D(D7118_Y), .RN(D5683_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D7144 ( .Q(D7144_Q), .D(D7130_Y), .RN(D5683_Y),     .CK(D191_QN));
KC_DFFRNHQ_X1 D6481 ( .Q(D6481_Q), .D(D6440_Y), .RN(D6463_Y),     .CK(D6462_Y));
KC_DFFRNHQ_X1 D6480 ( .Q(D6480_Q), .D(D5072_Y), .RN(D6463_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D6387 ( .Q(D6387_Q), .D(D457_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D6386 ( .Q(D6386_Q), .D(D7810_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D6385 ( .Q(D6385_Q), .D(D7814_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D6384 ( .Q(D6384_Q), .D(D7809_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D6383 ( .Q(D6383_Q), .D(D7806_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D6382 ( .Q(D6382_Q), .D(D7812_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D6381 ( .Q(D6381_Q), .D(D1953_Y), .RN(D7786_Y),     .CK(D6462_Y));
KC_DFFRNHQ_X1 D6351 ( .Q(D6351_Q), .D(D6323_Y), .RN(D7893_Y),     .CK(D6321_Y));
KC_DFFRNHQ_X1 D6345 ( .Q(D6345_Q), .D(D6317_Y), .RN(D7893_Y),     .CK(D6321_Y));
KC_DFFRNHQ_X1 D6344 ( .Q(D6344_Q), .D(D1958_Y), .RN(D965_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D6073 ( .Q(D6073_Q), .D(D6051_Y), .RN(D4483_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D5693 ( .Q(D5693_Q), .D(D5794_Y), .RN(D5683_Y),     .CK(D5799_Y));
KC_DFFRNHQ_X1 D5692 ( .Q(D5692_Q), .D(D7126_Y), .RN(D5683_Y),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D5691 ( .Q(D5691_Q), .D(D5819_Y), .RN(D5683_Y),     .CK(D5800_QN));
KC_DFFRNHQ_X1 D5690 ( .Q(D5690_Q), .D(D5781_Y), .RN(D5683_Y),     .CK(D5800_QN));
KC_DFFRNHQ_X1 D5689 ( .Q(D5689_Q), .D(D5750_Y), .RN(D5683_Y),     .CK(D5800_QN));
KC_DFFRNHQ_X1 D5688 ( .Q(D5688_Q), .D(D5914_Y), .RN(D5683_Y),     .CK(D5800_QN));
KC_DFFRNHQ_X1 D5687 ( .Q(D5687_Q), .D(D5785_Y), .RN(D5683_Y),     .CK(D5800_QN));
KC_DFFRNHQ_X1 D5686 ( .Q(D5686_Q), .D(D5784_Y), .RN(D5683_Y),     .CK(D5800_QN));
KC_DFFRNHQ_X1 D4826 ( .Q(D4826_Q), .D(D4795_Y), .RN(D4827_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D4825 ( .Q(D4825_Q), .D(D4794_Y), .RN(D965_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D4824 ( .Q(D4824_Q), .D(D4790_Y), .RN(D965_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D4823 ( .Q(D4823_Q), .D(D4792_Y), .RN(D965_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D4822 ( .Q(D4822_Q), .D(D4776_Y), .RN(D4827_Y),     .CK(D380_QN));
KC_DFFRNHQ_X1 D4821 ( .Q(D4821_Q), .D(D4837_Y), .RN(D965_Y),     .CK(D380_QN));
KC_DFFRNHQ_X1 D4820 ( .Q(D4820_Q), .D(D4810_Y), .RN(D965_Y),     .CK(D380_QN));
KC_DFFRNHQ_X1 D4819 ( .Q(D4819_Q), .D(D4766_Y), .RN(D4827_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D4818 ( .Q(D4818_Q), .D(D4809_Y), .RN(D965_Y),     .CK(D380_QN));
KC_DFFRNHQ_X1 D4817 ( .Q(D4817_Q), .D(D4800_Y), .RN(D4827_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D4729 ( .Q(D4729_Q), .D(D4667_Y), .RN(D4827_Y),     .CK(D4799_Y));
KC_DFFRNHQ_X1 D4728 ( .Q(D4728_Q), .D(D4722_Y), .RN(D4827_Y),     .CK(D4799_Y));
KC_DFFRNHQ_X1 D4727 ( .Q(D4727_Q), .D(D4723_Y), .RN(D4827_Y),     .CK(D4799_Y));
KC_DFFRNHQ_X1 D4641 ( .Q(D4641_Q), .D(D341_Y), .RN(D1934_Y),     .CK(D4527_Y));
KC_DFFRNHQ_X1 D4640 ( .Q(D4640_Q), .D(D4597_Y), .RN(D4634_Y),     .CK(D3178_QN));
KC_DFFRNHQ_X1 D4639 ( .Q(D4639_Q), .D(D4624_Y), .RN(D1934_Y),     .CK(D4527_Y));
KC_DFFRNHQ_X1 D4638 ( .Q(D4638_Q), .D(D4584_Y), .RN(D4634_Y),     .CK(D3178_QN));
KC_DFFRNHQ_X1 D4637 ( .Q(D4637_Q), .D(D4609_Y), .RN(D4634_Y),     .CK(D3178_QN));
KC_DFFRNHQ_X1 D4636 ( .Q(D4636_Q), .D(D4583_Y), .RN(D4634_Y),     .CK(D3178_QN));
KC_DFFRNHQ_X1 D4556 ( .Q(D4556_Q), .D(D4529_Y), .RN(D1934_Y),     .CK(D4527_Y));
KC_DFFRNHQ_X1 D4555 ( .Q(D4555_Q), .D(D4536_Y), .RN(D1934_Y),     .CK(D4527_Y));
KC_DFFRNHQ_X1 D4488 ( .Q(D4488_Q), .D(D4494_Y), .RN(D1652_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D4491 ( .Q(D4491_Q), .D(D16773_Y), .RN(D1652_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D4490 ( .Q(D4490_Q), .D(D4463_Y), .RN(D1652_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D4489 ( .Q(D4489_Q), .D(D4433_Y), .RN(D1652_Y),     .CK(D5931_QN));
KC_DFFRNHQ_X1 D4487 ( .Q(D4487_Q), .D(D4464_Y), .RN(D1652_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D4486 ( .Q(D4486_Q), .D(D2957_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D4485 ( .Q(D4485_Q), .D(D2959_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D4235 ( .Q(D4235_Q), .D(D4170_Y), .RN(D4461_Y),     .CK(D5931_QN));
KC_DFFRNHQ_X1 D4136 ( .Q(D4136_Q), .D(D4229_Y), .RN(D4461_Y),     .CK(D5799_Y));
KC_DFFRNHQ_X1 D4122 ( .Q(D4122_Q), .D(D198_Y), .RN(D5683_Y),     .CK(D5679_QN));
KC_DFFRNHQ_X1 D4121 ( .Q(D4121_Q), .D(D5674_Y), .RN(D5683_Y),     .CK(D5679_QN));
KC_DFFRNHQ_X1 D4120 ( .Q(D4120_Q), .D(D5702_Y), .RN(D5683_Y),     .CK(D5679_QN));
KC_DFFRNHQ_X1 D4119 ( .Q(D4119_Q), .D(D184_Y), .RN(D5683_Y),     .CK(D5679_QN));
KC_DFFRNHQ_X1 D4118 ( .Q(D4118_Q), .D(D4107_Y), .RN(D5683_Y),     .CK(D5679_QN));
KC_DFFRNHQ_X1 D3700 ( .Q(D3700_Q), .D(D1461_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3648 ( .Q(D3648_Q), .D(D3617_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3647 ( .Q(D3647_Q), .D(D3619_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3646 ( .Q(D3646_Q), .D(D3615_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3645 ( .Q(D3645_Q), .D(D3608_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3644 ( .Q(D3644_Q), .D(D3606_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3643 ( .Q(D3643_Q), .D(D3612_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3642 ( .Q(D3642_Q), .D(D3601_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3641 ( .Q(D3641_Q), .D(D1462_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3640 ( .Q(D3640_Q), .D(D3613_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3639 ( .Q(D3639_Q), .D(D3605_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3638 ( .Q(D3638_Q), .D(D3621_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3637 ( .Q(D3637_Q), .D(D3620_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3636 ( .Q(D3636_Q), .D(D3616_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3635 ( .Q(D3635_Q), .D(D3614_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3580 ( .Q(D3580_Q), .D(D1534_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3579 ( .Q(D3579_Q), .D(D3623_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D3484 ( .Q(D3484_Q), .D(D3424_Y), .RN(D3542_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D3483 ( .Q(D3483_Q), .D(D3425_Y), .RN(D3542_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D3482 ( .Q(D3482_Q), .D(D3436_Y), .RN(D3542_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D3481 ( .Q(D3481_Q), .D(D3464_Y), .RN(D3542_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D3388 ( .Q(D3388_Q), .D(D3466_Y), .RN(D3542_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D3387 ( .Q(D3387_Q), .D(D3240_Y), .RN(D4827_Y),     .CK(D3271_QN));
KC_DFFRNHQ_X1 D3386 ( .Q(D3386_Q), .D(D3324_Y), .RN(D4827_Y),     .CK(D3271_QN));
KC_DFFRNHQ_X1 D3385 ( .Q(D3385_Q), .D(D412_Y), .RN(D4827_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D3384 ( .Q(D3384_Q), .D(D3316_Y), .RN(D4827_Y),     .CK(D3271_QN));
KC_DFFRNHQ_X1 D3383 ( .Q(D3383_Q), .D(D3358_Y), .RN(D4827_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D3382 ( .Q(D3382_Q), .D(D3328_Y), .RN(D4827_Y),     .CK(D3271_QN));
KC_DFFRNHQ_X1 D3283 ( .Q(D3283_Q), .D(D3236_Y), .RN(D4827_Y),     .CK(D3176_QN));
KC_DFFRNHQ_X1 D3282 ( .Q(D3282_Q), .D(D3233_Y), .RN(D4827_Y),     .CK(D3176_QN));
KC_DFFRNHQ_X1 D3281 ( .Q(D3281_Q), .D(D3254_Y), .RN(D4827_Y),     .CK(D3176_QN));
KC_DFFRNHQ_X1 D3280 ( .Q(D3280_Q), .D(D3216_Y), .RN(D4827_Y),     .CK(D3271_QN));
KC_DFFRNHQ_X1 D3190 ( .Q(D3190_Q), .D(D3115_Y), .RN(D4634_Y),     .CK(D3177_QN));
KC_DFFRNHQ_X1 D3189 ( .Q(D3189_Q), .D(D3160_Y), .RN(D4634_Y),     .CK(D3177_QN));
KC_DFFRNHQ_X1 D3188 ( .Q(D3188_Q), .D(D3109_Y), .RN(D4634_Y),     .CK(D3177_QN));
KC_DFFRNHQ_X1 D3187 ( .Q(D3187_Q), .D(D3168_Y), .RN(D4634_Y),     .CK(D3177_QN));
KC_DFFRNHQ_X1 D3186 ( .Q(D3186_Q), .D(D3101_Y), .RN(D4634_Y),     .CK(D3177_QN));
KC_DFFRNHQ_X1 D3185 ( .Q(D3185_Q), .D(D3099_Y), .RN(D4634_Y),     .CK(D3177_QN));
KC_DFFRNHQ_X1 D3184 ( .Q(D3184_Q), .D(D1420_Y), .RN(D4634_Y),     .CK(D3176_QN));
KC_DFFRNHQ_X1 D3093 ( .Q(D3093_Q), .D(D1470_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D3084 ( .Q(D3084_Q), .D(D3047_Y), .RN(D4634_Y),     .CK(D3179_QN));
KC_DFFRNHQ_X1 D3083 ( .Q(D3083_Q), .D(D3060_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D3082 ( .Q(D3082_Q), .D(D317_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D3081 ( .Q(D3081_Q), .D(D3058_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D3080 ( .Q(D3080_Q), .D(D3164_Y), .RN(D4634_Y),     .CK(D3179_QN));
KC_DFFRNHQ_X1 D3079 ( .Q(D3079_Q), .D(D49_Y), .RN(D4634_Y),     .CK(D3179_QN));
KC_DFFRNHQ_X1 D3078 ( .Q(D3078_Q), .D(D3173_Y), .RN(D4634_Y),     .CK(D3179_QN));
KC_DFFRNHQ_X1 D3077 ( .Q(D3077_Q), .D(D3059_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D3004 ( .Q(D3004_Q), .D(D3006_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D3003 ( .Q(D3003_Q), .D(D2974_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D3002 ( .Q(D3002_Q), .D(D2972_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D3001 ( .Q(D3001_Q), .D(D2963_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D3000 ( .Q(D3000_Q), .D(D2913_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D2999 ( .Q(D2999_Q), .D(D2912_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D2891 ( .Q(D2891_Q), .D(D2897_Y), .RN(D2882_Y),     .CK(D2864_Y));
KC_DFFRNHQ_X1 D2890 ( .Q(D2890_Q), .D(D2841_Y), .RN(D2882_Y),     .CK(D2864_Y));
KC_DFFRNHQ_X1 D2889 ( .Q(D2889_Q), .D(D2879_Y), .RN(D2882_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D2888 ( .Q(D2888_Q), .D(D2840_Y), .RN(D2882_Y),     .CK(D2864_Y));
KC_DFFRNHQ_X1 D2887 ( .Q(D2887_Q), .D(D2837_Y), .RN(D2882_Y),     .CK(D2864_Y));
KC_DFFRNHQ_X1 D2886 ( .Q(D2886_Q), .D(D2835_Y), .RN(D2882_Y),     .CK(D7962_Y));
KC_DFFRNHQ_X1 D2885 ( .Q(D2885_Q), .D(D2872_Y), .RN(D2882_Y),     .CK(D2864_Y));
KC_DFFRNHQ_X1 D2884 ( .Q(D2884_Q), .D(D2828_Y), .RN(D2882_Y),     .CK(D2864_Y));
KC_DFFRNHQ_X1 D2883 ( .Q(D2883_Q), .D(D2976_Y), .RN(D2882_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D2801 ( .Q(D2801_Q), .D(D2789_Y), .RN(D2882_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D2800 ( .Q(D2800_Q), .D(D2806_Y), .RN(D2882_Y),     .CK(D2864_Y));
KC_DFFRNHQ_X1 D2799 ( .Q(D2799_Q), .D(D2786_Y), .RN(D4483_Y),     .CK(D2790_QN));
KC_DFFRNHQ_X1 D2798 ( .Q(D2798_Q), .D(D2779_Y), .RN(D4483_Y),     .CK(D2790_QN));
KC_DFFRNHQ_X1 D2797 ( .Q(D2797_Q), .D(D2787_Y), .RN(D4483_Y),     .CK(D2790_QN));
KC_DFFRNHQ_X1 D2796 ( .Q(D2796_Q), .D(D2807_Y), .RN(D4483_Y),     .CK(D2790_QN));
KC_DFFRNHQ_X1 D2795 ( .Q(D2795_Q), .D(D2742_Y), .RN(D2882_Y),     .CK(D2790_QN));
KC_DFFRNHQ_X1 D2794 ( .Q(D2794_Q), .D(D2774_Y), .RN(D2882_Y),     .CK(D2790_QN));
KC_DFFRNHQ_X1 D2681 ( .Q(D2681_Q), .D(D2664_Y), .RN(D16383_Y),     .CK(D2513_QN));
KC_DFFRNHQ_X1 D2680 ( .Q(D2680_Q), .D(D16196_Y), .RN(D15652_Y),     .CK(D2568_Y));
KC_DFFRNHQ_X1 D2679 ( .Q(D2679_Q), .D(D2676_Y), .RN(D2677_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D2678 ( .Q(D2678_Q), .D(D16351_Y), .RN(D16352_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D2641 ( .Q(D2641_Q), .D(D15683_Y), .RN(D2677_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D2640 ( .Q(D2640_Q), .D(D15763_Y), .RN(D15790_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D2639 ( .Q(D2639_Q), .D(D15773_Y), .RN(D15790_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D2638 ( .Q(D2638_Q), .D(D15851_Y), .RN(D16352_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D2574 ( .Q(D2574_Q), .D(D14546_Y), .RN(D13185_Y),     .CK(D14579_Y));
KC_DFFRNHQ_X1 D2573 ( .Q(D2573_Q), .D(D2560_Y), .RN(D15790_Y),     .CK(D14162_QN));
KC_DFFRNHQ_X1 D2572 ( .Q(D2572_Q), .D(D2551_Y), .RN(D14291_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D2524 ( .Q(D2524_Q), .D(D2550_Y), .RN(D14288_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D2523 ( .Q(D2523_Q), .D(D1191_Y), .RN(D14288_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D2518 ( .Q(D2518_Q), .D(D14079_Y), .RN(D13265_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D2517 ( .Q(D2517_Q), .D(D14758_Y), .RN(D14163_Y),     .CK(D14112_QN));
KC_DFFRNHQ_X1 D2516 ( .Q(D2516_Q), .D(D2676_Y), .RN(D14296_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D2515 ( .Q(D2515_Q), .D(D14786_Y), .RN(D14296_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D2474 ( .Q(D2474_Q), .D(D762_Y), .RN(D13758_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D2469 ( .Q(D2469_Q), .D(D13164_Y), .RN(D12679_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X1 D2468 ( .Q(D2468_Q), .D(D13684_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D2393 ( .Q(D2393_Q), .D(D12868_Y), .RN(D12846_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D2392 ( .Q(D2392_Q), .D(D12906_Y), .RN(D12846_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D2391 ( .Q(D2391_Q), .D(D2425_Y), .RN(D12898_Y),     .CK(D12975_Y));
KC_DFFRNHQ_X1 D2390 ( .Q(D2390_Q), .D(D2365_Y), .RN(D12679_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D2355 ( .Q(D2355_Q), .D(D12331_Y), .RN(D12339_Y),     .CK(D12831_Y));
KC_DFFRNHQ_X1 D2175 ( .Q(D2175_Q), .D(D10305_Q), .RN(D10357_Y),     .CK(D10706_Y));
KC_DFFRNHQ_X1 D2168 ( .Q(D2168_Q), .D(D9566_Y), .RN(D9538_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D2167 ( .Q(D2167_Q), .D(D10139_Y), .RN(D9271_Y),     .CK(D9212_QN));
KC_DFFRNHQ_X1 D2166 ( .Q(D2166_Q), .D(D9998_Y), .RN(D8818_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D2094 ( .Q(D2094_Q), .D(D9251_Y), .RN(D7892_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D2093 ( .Q(D2093_Q), .D(D9204_Y), .RN(D9128_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D2092 ( .Q(D2092_Q), .D(D9196_Y), .RN(D7788_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D2091 ( .Q(D2091_Q), .D(D9138_Y), .RN(D9214_Y),     .CK(D9141_QN));
KC_DFFRNHQ_X1 D2090 ( .Q(D2090_Q), .D(D8868_Y), .RN(D8818_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D1944 ( .Q(D1944_Q), .D(D8266_Y), .RN(D8229_Y),     .CK(D9458_QN));
KC_DFFRNHQ_X1 D1943 ( .Q(D1943_Q), .D(D8342_Q), .RN(D8300_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D1942 ( .Q(D1942_Q), .D(D3379_Y), .RN(D7880_Y),     .CK(D4799_Y));
KC_DFFRNHQ_X1 D1941 ( .Q(D1941_Q), .D(D6457_Y), .RN(D7880_Y),     .CK(D6462_Y));
KC_DFFRNHQ_X1 D1940 ( .Q(D1940_Q), .D(D1902_Y), .RN(D7880_Y),     .CK(D503_QN));
KC_DFFRNHQ_X1 D1793 ( .Q(D1793_Q), .D(D6487_Y), .RN(D7786_Y),     .CK(D6462_Y));
KC_DFFRNHQ_X1 D1792 ( .Q(D1792_Q), .D(D1959_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D1791 ( .Q(D1791_Q), .D(D7798_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D1655 ( .Q(D1655_Q), .D(D4793_Y), .RN(D965_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D1654 ( .Q(D1654_Q), .D(D4791_Y), .RN(D965_Y),     .CK(D3367_QN));
KC_DFFRNHQ_X1 D1527 ( .Q(D1527_Q), .D(D3440_Y), .RN(D3542_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D1518 ( .Q(D1518_Q), .D(D1464_Y), .RN(D3577_Y),     .CK(D3668_Y));
KC_DFFRNHQ_X1 D1517 ( .Q(D1517_Q), .D(D3491_Y), .RN(D3542_Y),     .CK(D4957_QN));
KC_DFFRNHQ_X1 D1516 ( .Q(D1516_Q), .D(D54_Y), .RN(D4634_Y),     .CK(D3179_QN));
KC_DFFRNHQ_X1 D1515 ( .Q(D1515_Q), .D(D3147_Y), .RN(D4634_Y),     .CK(D3179_QN));
KC_DFFRNHQ_X1 D1514 ( .Q(D1514_Q), .D(D19_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D1401 ( .Q(D1401_Q), .D(D2500_Y), .RN(D14474_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D1400 ( .Q(D1400_Q), .D(D16625_Y), .RN(D16579_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D1396 ( .Q(D1396_Q), .D(D16626_Y), .RN(D16579_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D1395 ( .Q(D1395_Q), .D(D16673_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D1386 ( .Q(D1386_Q), .D(D15838_Y), .RN(D14489_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D1385 ( .Q(D1385_Q), .D(D16527_Y), .RN(D16376_Y),     .CK(D16515_QN));
KC_DFFRNHQ_X1 D1384 ( .Q(D1384_Q), .D(D15128_Y), .RN(D15990_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D1383 ( .Q(D1383_Q), .D(D14760_Y), .RN(D14489_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D1382 ( .Q(D1382_Q), .D(D15113_Y), .RN(D14489_Y),     .CK(D13745_Y));
KC_DFFRNHQ_X1 D1381 ( .Q(D1381_Q), .D(D16509_Y), .RN(D16376_Y),     .CK(D16515_QN));
KC_DFFRNHQ_X1 D1380 ( .Q(D1380_Q), .D(D15789_Y), .RN(D15990_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D1379 ( .Q(D1379_Q), .D(D14760_Y), .RN(D14489_Y),     .CK(D14469_Y));
KC_DFFRNHQ_X1 D1378 ( .Q(D1378_Q), .D(D16409_Y), .RN(D16376_Y),     .CK(D16476_Y));
KC_DFFRNHQ_X1 D1377 ( .Q(D1377_Q), .D(D1282_Y), .RN(D15990_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D1376 ( .Q(D1376_Q), .D(D15199_Y), .RN(D14489_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D1375 ( .Q(D1375_Q), .D(D15113_Y), .RN(D14474_Y),     .CK(D1345_Y));
KC_DFFRNHQ_X1 D1374 ( .Q(D1374_Q), .D(D16605_Y), .RN(D16579_Y),     .CK(D16581_Y));
KC_DFFRNHQ_X1 D1373 ( .Q(D1373_Q), .D(D16674_Y), .RN(D16610_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D1327 ( .Q(D1327_Q), .D(D95_Y), .RN(D14291_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D1326 ( .Q(D1326_Q), .D(D15972_Y), .RN(D15990_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D1325 ( .Q(D1325_Q), .D(D15204_Y), .RN(D14489_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D1324 ( .Q(D1324_Q), .D(D16447_Y), .RN(D16377_Y),     .CK(D16476_Y));
KC_DFFRNHQ_X1 D1323 ( .Q(D1323_Q), .D(D15188_Y), .RN(D14489_Y),     .CK(D15219_Y));
KC_DFFRNHQ_X1 D1322 ( .Q(D1322_Q), .D(D16450_Y), .RN(D16377_Y),     .CK(D16476_Y));
KC_DFFRNHQ_X1 D1321 ( .Q(D1321_Q), .D(D13796_Y), .RN(D14474_Y),     .CK(D13794_Y));
KC_DFFRNHQ_X1 D1320 ( .Q(D1320_Q), .D(D16622_Y), .RN(D16579_Y),     .CK(D1402_QN));
KC_DFFRNHQ_X1 D1236 ( .Q(D1236_Q), .D(D16381_Y), .RN(D16384_Y),     .CK(D14466_Y));
KC_DFFRNHQ_X1 D1235 ( .Q(D1235_Q), .D(D13682_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D1234 ( .Q(D1234_Q), .D(D15850_Y), .RN(D965_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D1233 ( .Q(D1233_Q), .D(D15928_Y), .RN(D16384_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D1232 ( .Q(D1232_Q), .D(D15117_Y), .RN(D14291_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D1231 ( .Q(D1231_Q), .D(D15927_Y), .RN(D16384_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D1230 ( .Q(D1230_Q), .D(D1189_Y), .RN(D14291_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D1229 ( .Q(D1229_Q), .D(D16381_Y), .RN(D16384_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D1228 ( .Q(D1228_Q), .D(D16381_Y), .RN(D16384_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D1163 ( .Q(D1163_Q), .D(D15053_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D1159 ( .Q(D1159_Q), .D(D13030_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D1158 ( .Q(D1158_Q), .D(D15056_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D1157 ( .Q(D1157_Q), .D(D15062_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D1156 ( .Q(D1156_Q), .D(D15848_Y), .RN(D16352_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D1155 ( .Q(D1155_Q), .D(D2676_Y), .RN(D14296_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D1154 ( .Q(D1154_Q), .D(D15688_Y), .RN(D14296_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D1153 ( .Q(D1153_Q), .D(D15050_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D1152 ( .Q(D1152_Q), .D(D13688_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D1151 ( .Q(D1151_Q), .D(D15059_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D1150 ( .Q(D1150_Q), .D(D13679_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D1149 ( .Q(D1149_Q), .D(D15844_Y), .RN(D16352_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D1148 ( .Q(D1148_Q), .D(D15846_Y), .RN(D16352_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D1147 ( .Q(D1147_Q), .D(D1164_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D1077 ( .Q(D1077_Q), .D(D2666_Y), .RN(D2677_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D1074 ( .Q(D1074_Q), .D(D2666_Y), .RN(D2627_Y),     .CK(D14983_Y));
KC_DFFRNHQ_X1 D1070 ( .Q(D1070_Q), .D(D15758_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D1066 ( .Q(D1066_Q), .D(D15765_Y), .RN(D14869_Y),     .CK(D14229_Y));
KC_DFFRNHQ_X1 D1065 ( .Q(D1065_Q), .D(D14972_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D1054 ( .Q(D1054_Q), .D(D15683_Y), .RN(D14869_Y),     .CK(D14987_Y));
KC_DFFRNHQ_X1 D1053 ( .Q(D1053_Q), .D(D996_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D1052 ( .Q(D1052_Q), .D(D14970_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D1051 ( .Q(D1051_Q), .D(D14961_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D1050 ( .Q(D1050_Q), .D(D15751_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D1048 ( .Q(D1048_Q), .D(D14963_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D956 ( .Q(D956_Q), .D(D2451_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D954 ( .Q(D954_Q), .D(D13427_Y), .RN(D14163_Y),     .CK(D13511_Y));
KC_DFFRNHQ_X1 D953 ( .Q(D953_Q), .D(D15683_Y), .RN(D14869_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D952 ( .Q(D952_Q), .D(D97_Y), .RN(D14869_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D951 ( .Q(D951_Q), .D(D9639_Q), .RN(D10357_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D934 ( .Q(D934_Q), .D(D10365_Q), .RN(D10357_Y),     .CK(D2176_Y));
KC_DFFRNHQ_X1 D933 ( .Q(D933_Q), .D(D9601_Y), .RN(D8319_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D932 ( .Q(D932_Q), .D(D12868_Y), .RN(D12900_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D931 ( .Q(D931_Q), .D(D12890_Y), .RN(D12900_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D930 ( .Q(D930_Q), .D(D13465_Y), .RN(D14163_Y),     .CK(D13511_Y));
KC_DFFRNHQ_X1 D929 ( .Q(D929_Q), .D(D2453_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D928 ( .Q(D928_Q), .D(D14131_Y), .RN(D14163_Y),     .CK(D13511_Y));
KC_DFFRNHQ_X1 D927 ( .Q(D927_Q), .D(D12868_Y), .RN(D12900_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D926 ( .Q(D926_Q), .D(D15583_Y), .RN(D14163_Y),     .CK(D14231_Y));
KC_DFFRNHQ_X1 D925 ( .Q(D925_Q), .D(D15587_Y), .RN(D2677_Y),     .CK(D2631_Y));
KC_DFFRNHQ_X1 D924 ( .Q(D924_Q), .D(D15769_Y), .RN(D15790_Y),     .CK(D14992_Y));
KC_DFFRNHQ_X1 D856 ( .Q(D856_Q), .D(D14051_Y), .RN(D14474_Y),     .CK(D13261_QN));
KC_DFFRNHQ_X1 D855 ( .Q(D855_Q), .D(D13413_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D853 ( .Q(D853_Q), .D(D14766_Y), .RN(D14163_Y),     .CK(D14080_QN));
KC_DFFRNHQ_X1 D852 ( .Q(D852_Q), .D(D13412_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D851 ( .Q(D851_Q), .D(D15609_Y), .RN(D15652_Y),     .CK(D2568_Y));
KC_DFFRNHQ_X1 D843 ( .Q(D843_Q), .D(D12821_Y), .RN(D10725_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D842 ( .Q(D842_Q), .D(D12890_Y), .RN(D12846_Y),     .CK(D12742_QN));
KC_DFFRNHQ_X1 D836 ( .Q(D836_Q), .D(D10316_Q), .RN(D10726_Y),     .CK(D11631_Y));
KC_DFFRNHQ_X1 D827 ( .Q(D827_Q), .D(D9515_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D826 ( .Q(D826_Q), .D(D8123_Y), .RN(D12838_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D825 ( .Q(D825_Q), .D(D10259_Y), .RN(D12838_Y),     .CK(D9569_QN));
KC_DFFRNHQ_X1 D824 ( .Q(D824_Q), .D(D9492_Y), .RN(D12838_Y),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D823 ( .Q(D823_Q), .D(D12806_Y), .RN(D10725_Y),     .CK(D780_QN));
KC_DFFRNHQ_X1 D822 ( .Q(D822_Q), .D(D12806_Y), .RN(D12258_Y),     .CK(D782_QN));
KC_DFFRNHQ_X1 D821 ( .Q(D821_Q), .D(D12806_Y), .RN(D12258_Y),     .CK(D12843_QN));
KC_DFFRNHQ_X1 D820 ( .Q(D820_Q), .D(D14803_Y), .RN(D13265_Y),     .CK(D13261_QN));
KC_DFFRNHQ_X1 D819 ( .Q(D819_Q), .D(D753_Y), .RN(D12846_Y),     .CK(D13251_Y));
KC_DFFRNHQ_X1 D818 ( .Q(D818_Q), .D(D14769_Y), .RN(D14163_Y),     .CK(D13261_QN));
KC_DFFRNHQ_X1 D817 ( .Q(D817_Q), .D(D14767_Y), .RN(D14163_Y),     .CK(D13261_QN));
KC_DFFRNHQ_X1 D816 ( .Q(D816_Q), .D(D16194_Y), .RN(D16383_Y),     .CK(D2568_Y));
KC_DFFRNHQ_X1 D815 ( .Q(D815_Q), .D(D14763_Y), .RN(D14163_Y),     .CK(D14080_QN));
KC_DFFRNHQ_X1 D814 ( .Q(D814_Q), .D(D13407_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D722 ( .Q(D722_Q), .D(D14611_Y), .RN(D13265_Y),     .CK(D13263_QN));
KC_DFFRNHQ_X1 D721 ( .Q(D721_Q), .D(D14613_Y), .RN(D13265_Y),     .CK(D13263_QN));
KC_DFFRNHQ_X1 D717 ( .Q(D717_Q), .D(D12726_Y), .RN(D12258_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D716 ( .Q(D716_Q), .D(D12730_Y), .RN(D12258_Y),     .CK(D12827_Y));
KC_DFFRNHQ_X1 D704 ( .Q(D704_Q), .D(D9438_Y), .RN(D9375_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D703 ( .Q(D703_Q), .D(D715_Y), .RN(D9381_Y),     .CK(D8142_QN));
KC_DFFRNHQ_X1 D702 ( .Q(D702_Q), .D(D10238_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D701 ( .Q(D701_Q), .D(D10202_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D700 ( .Q(D700_Q), .D(D9429_Y), .RN(D9381_Y),     .CK(D9570_QN));
KC_DFFRNHQ_X1 D699 ( .Q(D699_Q), .D(D77_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D698 ( .Q(D698_Q), .D(D10222_Q), .RN(D10726_Y),     .CK(D10707_Y));
KC_DFFRNHQ_X1 D697 ( .Q(D697_Q), .D(D14078_Y), .RN(D13266_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D696 ( .Q(D696_Q), .D(D13250_Y), .RN(D13266_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D695 ( .Q(D695_Q), .D(D13386_Y), .RN(D13266_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D694 ( .Q(D694_Q), .D(D13250_Y), .RN(D13266_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D693 ( .Q(D693_Q), .D(D14078_Y), .RN(D13266_Y),     .CK(D13214_QN));
KC_DFFRNHQ_X1 D692 ( .Q(D692_Q), .D(D13399_Y), .RN(D13266_Y),     .CK(D12745_QN));
KC_DFFRNHQ_X1 D691 ( .Q(D691_Q), .D(D13399_Y), .RN(D13266_Y),     .CK(D12677_QN));
KC_DFFRNHQ_X1 D619 ( .Q(D619_Q), .D(D12665_Y), .RN(D13194_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D618 ( .Q(D618_Q), .D(D12673_Y), .RN(D13194_Y),     .CK(D13193_QN));
KC_DFFRNHQ_X1 D609 ( .Q(D609_Q), .D(D581_Y), .RN(D9374_Y),     .CK(D9447_Y));
KC_DFFRNHQ_X1 D608 ( .Q(D608_Q), .D(D14568_Y), .RN(D13185_Y),     .CK(D14579_Y));
KC_DFFRNHQ_X1 D607 ( .Q(D607_Q), .D(D12672_Y), .RN(D13194_Y),     .CK(D13262_QN));
KC_DFFRNHQ_X1 D605 ( .Q(D605_Q), .D(D12215_Y), .RN(D12734_Y),     .CK(D11713_QN));
KC_DFFRNHQ_X1 D543 ( .Q(D543_Q), .D(D13852_Y), .RN(D13185_Y),     .CK(D506_QN));
KC_DFFRNHQ_X1 D533 ( .Q(D533_Q), .D(D472_Y), .RN(D9375_Y),     .CK(D503_QN));
KC_DFFRNHQ_X1 D532 ( .Q(D532_Q), .D(D7826_Y), .RN(D9375_Y),     .CK(D503_QN));
KC_DFFRNHQ_X1 D531 ( .Q(D531_Q), .D(D1851_Y), .RN(D9375_Y),     .CK(D503_QN));
KC_DFFRNHQ_X1 D530 ( .Q(D530_Q), .D(D12665_Y), .RN(D13194_Y),     .CK(D13193_QN));
KC_DFFRNHQ_X1 D529 ( .Q(D529_Q), .D(D13849_Y), .RN(D13185_Y),     .CK(D506_QN));
KC_DFFRNHQ_X1 D485 ( .Q(D485_Q), .D(D1697_Y), .RN(D6463_Y),     .CK(D6462_Y));
KC_DFFRNHQ_X1 D484 ( .Q(D484_Q), .D(D9293_Y), .RN(D7892_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D483 ( .Q(D483_Q), .D(D9312_Y), .RN(D7892_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D482 ( .Q(D482_Q), .D(D9314_Y), .RN(D7892_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D452 ( .Q(D452_Q), .D(D7813_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D451 ( .Q(D451_Q), .D(D9256_Y), .RN(D9271_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D450 ( .Q(D450_Q), .D(D7778_Y), .RN(D7786_Y),     .CK(D6332_QN));
KC_DFFRNHQ_X1 D449 ( .Q(D449_Q), .D(D10138_Y), .RN(D7892_Y),     .CK(D415_QN));
KC_DFFRNHQ_X1 D421 ( .Q(D421_Q), .D(D10104_Y), .RN(D9271_Y),     .CK(D9142_QN));
KC_DFFRNHQ_X1 D420 ( .Q(D420_Q), .D(D7713_Y), .RN(VDD), .CK(D7575_Y));
KC_DFFRNHQ_X1 D419 ( .Q(D419_Q), .D(D423_Y), .RN(D9214_Y),     .CK(D9139_QN));
KC_DFFRNHQ_X1 D418 ( .Q(D418_Q), .D(D6324_Y), .RN(D7893_Y),     .CK(D6321_Y));
KC_DFFRNHQ_X1 D387 ( .Q(D387_Q), .D(D9161_Y), .RN(D9214_Y),     .CK(D443_QN));
KC_DFFRNHQ_X1 D386 ( .Q(D386_Q), .D(D9126_Y), .RN(D9214_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D385 ( .Q(D385_Q), .D(D9127_Y), .RN(D9214_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D384 ( .Q(D384_Q), .D(D6216_Y), .RN(D7795_Y),     .CK(D6321_Y));
KC_DFFRNHQ_X1 D354 ( .Q(D354_Q), .D(D10053_Y), .RN(D9128_Y),     .CK(D443_QN));
KC_DFFRNHQ_X1 D353 ( .Q(D353_Q), .D(D2173_Y), .RN(D9128_Y),     .CK(D443_QN));
KC_DFFRNHQ_X1 D334 ( .Q(D334_Q), .D(D9026_Y), .RN(D4461_Y),     .CK(D7466_QN));
KC_DFFRNHQ_X1 D328 ( .Q(D328_Q), .D(D4626_Y), .RN(D1652_Y),     .CK(D4527_Y));
KC_DFFRNHQ_X1 D326 ( .Q(D326_Q), .D(D10040_Y), .RN(D324_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D325 ( .Q(D325_Q), .D(D4541_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D305 ( .Q(D305_Q), .D(D10024_Y), .RN(D8894_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D304 ( .Q(D304_Q), .D(D4477_Y), .RN(D1652_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D303 ( .Q(D303_Q), .D(D292_Y), .RN(D8894_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D302 ( .Q(D302_Q), .D(D3007_Y), .RN(D1934_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D301 ( .Q(D301_Q), .D(D3005_Y), .RN(D1934_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D300 ( .Q(D300_Q), .D(D2969_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D299 ( .Q(D299_Q), .D(D2965_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D298 ( .Q(D298_Q), .D(D2905_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D297 ( .Q(D297_Q), .D(D2949_Y), .RN(D4553_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D268 ( .Q(D268_Q), .D(D7405_Y), .RN(D4461_Y),     .CK(D7712_Y));
KC_DFFRNHQ_X1 D265 ( .Q(D265_Q), .D(D2865_Y), .RN(D2882_Y),     .CK(D4543_Y));
KC_DFFRNHQ_X1 D264 ( .Q(D264_Q), .D(D4367_Y), .RN(D4461_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D233 ( .Q(D233_Q), .D(D9974_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D232 ( .Q(D232_Q), .D(D4230_Y), .RN(D4461_Y),     .CK(D5799_Y));
KC_DFFRNHQ_X1 D231 ( .Q(D231_Q), .D(D9957_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D230 ( .Q(D230_Q), .D(D9979_Y), .RN(D8818_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D229 ( .Q(D229_Q), .D(D225_Y), .RN(D4461_Y),     .CK(D5799_Y));
KC_DFFRNHQ_X1 D228 ( .Q(D228_Q), .D(D4236_Y), .RN(D4461_Y),     .CK(D5931_QN));
KC_DFFRNHQ_X1 D227 ( .Q(D227_Q), .D(D9975_Y), .RN(D8779_Y),     .CK(D8813_QN));
KC_DFFRNHQ_X1 D195 ( .Q(D195_Q), .D(D7277_Y), .RN(D8818_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D194 ( .Q(D194_Q), .D(D1669_Y), .RN(D4461_Y),     .CK(D5799_Y));
KC_DFFRNHQ_X1 D193 ( .Q(D193_Q), .D(D7159_Y), .RN(D7795_Y),     .CK(D7138_QN));
KC_DFFRNHQ_X1 D192 ( .Q(D192_Q), .D(D7139_Y), .RN(D5683_Y),     .CK(D191_QN));
KC_DFFRNHQ_X1 D146 ( .Q(D146_Q), .D(D13366_Y), .RN(D12901_Y),     .CK(D13388_QN));
KC_DFFRNHQ_X1 D164 ( .Q(D164_Q), .D(D13674_Y), .RN(D13758_Y),     .CK(D13698_Y));
KC_DFFRNHQ_X1 D155 ( .Q(D155_Q), .D(D9356_Q), .RN(D12302_Y),     .CK(D10176_Y));
KC_DFFRNHQ_X1 D154 ( .Q(D154_Q), .D(D9244_Y), .RN(D7892_Y),     .CK(D416_QN));
KC_DFFRNHQ_X1 D153 ( .Q(D153_Q), .D(D1847_Y), .RN(D7786_Y),     .CK(D6462_Y));
KC_DFFRNHQ_X1 D152 ( .Q(D152_Q), .D(D7891_Y), .RN(D9375_Y),     .CK(D503_QN));
KC_DFFRNHQ_X1 D151 ( .Q(D151_Q), .D(D2141_Y), .RN(D324_Y),     .CK(D296_QN));
KC_DFFRNHQ_X1 D150 ( .Q(D150_Q), .D(D3065_Y), .RN(D4553_Y),     .CK(D2791_QN));
KC_DFFRNHQ_X1 D149 ( .Q(D149_Q), .D(D7403_Y), .RN(D8894_Y),     .CK(D9211_QN));
KC_DFFRNHQ_X1 D148 ( .Q(D148_Q), .D(D4386_Y), .RN(D1652_Y),     .CK(D4462_Y));
KC_DFFRNHQ_X1 D147 ( .Q(D147_Q), .D(D258_Y), .RN(D8818_Y),     .CK(D261_QN));
KC_DFFRNHQ_X1 D145 ( .Q(D145_Q), .D(D15587_Y), .RN(D2677_Y),     .CK(D16348_Y));
KC_DFFRNHQ_X1 D144 ( .Q(D144_Q), .D(D15849_Y), .RN(D2677_Y),     .CK(D15807_Y));
KC_DFFRNHQ_X1 D143 ( .Q(D143_Q), .D(D2554_Y), .RN(D14296_Y),     .CK(D15083_Y));
KC_DFFRNHQ_X1 D142 ( .Q(D142_Q), .D(D2619_Y), .RN(D16352_Y),     .CK(D15934_Y));
KC_DFFRNHQ_X1 D141 ( .Q(D141_Q), .D(D11619_Y), .RN(D11636_SN),     .CK(D12174_Y));
KC_AOI21B_X1 D15453 ( .AN(D641_Y), .B0(D15394_Y), .Y(D15453_Y),     .B1(D15334_Y));
KC_AOI21B_X1 D14684 ( .AN(D14746_Y), .B0(D2509_Y), .Y(D14684_Y),     .B1(D8997_Y));
KC_AOI21B_X1 D13133 ( .AN(D13136_Y), .B0(D13803_Q), .Y(D13133_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D13131 ( .AN(D13099_Y), .B0(D2300_Y), .Y(D13131_Y),     .B1(D13819_Q));
KC_AOI21B_X1 D13130 ( .AN(D13151_Y), .B0(D13798_Q), .Y(D13130_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D13129 ( .AN(D13100_Y), .B0(D2300_Y), .Y(D13129_Y),     .B1(D13800_Q));
KC_AOI21B_X1 D13128 ( .AN(D13134_Y), .B0(D1358_Q), .Y(D13128_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D13127 ( .AN(D13141_Y), .B0(D2300_Y), .Y(D13127_Y),     .B1(D13803_Q));
KC_AOI21B_X1 D13126 ( .AN(D13137_Y), .B0(D13819_Q), .Y(D13126_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D13125 ( .AN(D13138_Y), .B0(D13800_Q), .Y(D13125_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D13124 ( .AN(D13139_Y), .B0(D2300_Y), .Y(D13124_Y),     .B1(D13798_Q));
KC_AOI21B_X1 D13123 ( .AN(D13135_Y), .B0(D2300_Y), .Y(D13123_Y),     .B1(D1358_Q));
KC_AOI21B_X1 D13122 ( .AN(D13142_Y), .B0(D2300_Y), .Y(D13122_Y),     .B1(D1304_Q));
KC_AOI21B_X1 D13121 ( .AN(D13140_Y), .B0(D1304_Q), .Y(D13121_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D13049 ( .AN(D13023_Y), .B0(D13042_Q), .Y(D13049_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D13048 ( .AN(D13013_Y), .B0(D13037_Q), .Y(D13048_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D13047 ( .AN(D13012_Y), .B0(D11970_Y), .Y(D13047_Y),     .B1(D13037_Q));
KC_AOI21B_X1 D13046 ( .AN(D13014_Y), .B0(D11970_Y), .Y(D13046_Y),     .B1(D13042_Q));
KC_AOI21B_X1 D12990 ( .AN(D13017_Y), .B0(D11970_Y), .Y(D12990_Y),     .B1(D12981_Q));
KC_AOI21B_X1 D12989 ( .AN(D13022_Y), .B0(D12981_Q), .Y(D12989_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D12747 ( .AN(D12732_Y), .B0(D12729_Y), .Y(D12747_Y),     .B1(D16199_Y));
KC_AOI21B_X1 D12616 ( .AN(D12604_Y), .B0(D2300_Y), .Y(D12616_Y),     .B1(D1313_Q));
KC_AOI21B_X1 D12595 ( .AN(D12603_Y), .B0(D1313_Q), .Y(D12595_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12594 ( .AN(D12597_Y), .B0(D2300_Y), .Y(D12594_Y),     .B1(D12573_Q));
KC_AOI21B_X1 D12593 ( .AN(D12600_Y), .B0(D12572_Q), .Y(D12593_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12592 ( .AN(D12596_Y), .B0(D12573_Q), .Y(D12592_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12591 ( .AN(D12598_Y), .B0(D12614_Q), .Y(D12591_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12590 ( .AN(D1337_Y), .B0(D13150_Q), .Y(D12590_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12589 ( .AN(D12601_Y), .B0(D2300_Y), .Y(D12589_Y),     .B1(D12572_Q));
KC_AOI21B_X1 D12588 ( .AN(D12602_Y), .B0(D2300_Y), .Y(D12588_Y),     .B1(D12617_Q));
KC_AOI21B_X1 D12587 ( .AN(D12599_Y), .B0(D2300_Y), .Y(D12587_Y),     .B1(D12614_Q));
KC_AOI21B_X1 D12586 ( .AN(D12606_Y), .B0(D12617_Q), .Y(D12586_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12510 ( .AN(D13024_Y), .B0(D11970_Y), .Y(D12510_Y),     .B1(D13036_Q));
KC_AOI21B_X1 D12509 ( .AN(D12472_Y), .B0(D11970_Y), .Y(D12509_Y),     .B1(D12498_Q));
KC_AOI21B_X1 D12508 ( .AN(D12473_Y), .B0(D12498_Q), .Y(D12508_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D12471 ( .AN(D982_Y), .B0(D11970_Y), .Y(D12471_Y),     .B1(D1039_Q));
KC_AOI21B_X1 D12470 ( .AN(D12945_Y), .B0(D1036_Q), .Y(D12470_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D12469 ( .AN(D12435_Y), .B0(D11970_Y), .Y(D12469_Y),     .B1(D1036_Q));
KC_AOI21B_X1 D12413 ( .AN(D82_Y), .B0(D916_Q), .Y(D12413_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D12412 ( .AN(D12379_Y), .B0(D11970_Y), .Y(D12412_Y),     .B1(D916_Q));
KC_AOI21B_X1 D12411 ( .AN(D2324_Y), .B0(D11970_Y), .Y(D12411_Y),     .B1(D912_Q));
KC_AOI21B_X1 D12124 ( .AN(D12110_Y), .B0(D2300_Y), .Y(D12124_Y),     .B1(D12091_Q));
KC_AOI21B_X1 D12103 ( .AN(D12111_Y), .B0(D12127_Q), .Y(D12103_Y),     .B1(D2300_Y));
KC_AOI21B_X1 D12102 ( .AN(D12106_Y), .B0(D12127_Q), .Y(D12102_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12101 ( .AN(D12105_Y), .B0(D12618_Q), .Y(D12101_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12100 ( .AN(D12107_Y), .B0(D12091_Q), .Y(D12100_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12099 ( .AN(D12109_Y), .B0(D12086_Q), .Y(D12099_Y),     .B1(D12048_Y));
KC_AOI21B_X1 D12098 ( .AN(D12060_Y), .B0(D2300_Y), .Y(D12098_Y),     .B1(D12086_Q));
KC_AOI21B_X1 D12097 ( .AN(D12108_Y), .B0(D2300_Y), .Y(D12097_Y),     .B1(D12618_Q));
KC_AOI21B_X1 D11988 ( .AN(D11935_Y), .B0(D12499_Q), .Y(D11988_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D11987 ( .AN(D11939_Y), .B0(D11970_Y), .Y(D11987_Y),     .B1(D11974_Q));
KC_AOI21B_X1 D11986 ( .AN(D11938_Y), .B0(D11974_Q), .Y(D11986_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D11985 ( .AN(D11937_Y), .B0(D11970_Y), .Y(D11985_Y),     .B1(D11976_Q));
KC_AOI21B_X1 D11984 ( .AN(D11936_Y), .B0(D11976_Q), .Y(D11984_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D11983 ( .AN(D11934_Y), .B0(D11970_Y), .Y(D11983_Y),     .B1(D12499_Q));
KC_AOI21B_X1 D11928 ( .AN(D2275_Y), .B0(D11970_Y), .Y(D11928_Y),     .B1(D1044_Q));
KC_AOI21B_X1 D11927 ( .AN(D11813_Y), .B0(D1044_Q), .Y(D11927_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D11877 ( .AN(D11812_Y), .B0(D918_Q), .Y(D11877_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D11876 ( .AN(D11814_Y), .B0(D11866_Q), .Y(D11876_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D11875 ( .AN(D11901_Y), .B0(D11865_Q), .Y(D11875_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D11874 ( .AN(D2274_Y), .B0(D11865_Q), .Y(D11874_Y),     .B1(D11970_Y));
KC_AOI21B_X1 D11873 ( .AN(D11811_Y), .B0(D11970_Y), .Y(D11873_Y),     .B1(D918_Q));
KC_AOI21B_X1 D11872 ( .AN(D11902_Y), .B0(D11970_Y), .Y(D11872_Y),     .B1(D11866_Q));
KC_AOI21B_X1 D11810 ( .AN(D11679_Y), .B0(D10776_Y), .Y(D11810_Y),     .B1(D11716_Q));
KC_AOI21B_X1 D11809 ( .AN(D11772_Y), .B0(D11800_Q), .Y(D11809_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D11808 ( .AN(D11690_Y), .B0(D11716_Q), .Y(D11808_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D11807 ( .AN(D11774_Y), .B0(D10776_Y), .Y(D11807_Y),     .B1(D11800_Q));
KC_AOI21B_X1 D11806 ( .AN(D11764_Y), .B0(D11797_Q), .Y(D11806_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D11805 ( .AN(D11766_Y), .B0(D10776_Y), .Y(D11805_Y),     .B1(D11797_Q));
KC_AOI21B_X1 D11730 ( .AN(D559_Y), .B0(D10776_Y), .Y(D11730_Y),     .B1(D11658_Q));
KC_AOI21B_X1 D11729 ( .AN(D11706_Y), .B0(D10776_Y), .Y(D11729_Y),     .B1(D126_Q));
KC_AOI21B_X1 D11728 ( .AN(D11693_Y), .B0(D10776_Y), .Y(D11728_Y),     .B1(D11721_Q));
KC_AOI21B_X1 D11727 ( .AN(D11694_Y), .B0(D11721_Q), .Y(D11727_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D11664 ( .AN(D11644_Y), .B0(D11658_Q), .Y(D11664_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D11663 ( .AN(D585_Y), .B0(D11671_Y), .Y(D11663_Y),     .B1(D10181_Y));
KC_AOI21B_X1 D11406 ( .AN(D11361_Y), .B0(D11391_Q), .Y(D11406_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D11405 ( .AN(D11368_Y), .B0(D11393_Q), .Y(D11405_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D11404 ( .AN(D11355_Y), .B0(D11388_Q), .Y(D11404_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D11403 ( .AN(D11360_Y), .B0(D11388_Q), .Y(D11403_Y),     .B1(D2227_Y));
KC_AOI21B_X1 D11344 ( .AN(D11282_Y), .B0(D2227_Y), .Y(D11344_Y),     .B1(D908_Q));
KC_AOI21B_X1 D11343 ( .AN(D11280_Y), .B0(D11336_Q), .Y(D11343_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D11278 ( .AN(D11141_Y), .B0(D10776_Y), .Y(D11278_Y),     .B1(D11179_Q));
KC_AOI21B_X1 D11277 ( .AN(D11227_Y), .B0(D11179_Q), .Y(D11277_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D11132 ( .AN(D11118_Y), .B0(D10776_Y), .Y(D11132_Y),     .B1(D11128_Q));
KC_AOI21B_X1 D11131 ( .AN(D11119_Y), .B0(D11128_Q), .Y(D11131_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D11130 ( .AN(D557_Y), .B0(D10776_Y), .Y(D11130_Y),     .B1(D11127_Q));
KC_AOI21B_X1 D11129 ( .AN(D11120_Y), .B0(D10776_Y), .Y(D11129_Y),     .B1(D2246_Q));
KC_AOI21B_X1 D11111 ( .AN(D11092_Y), .B0(D11108_Q), .Y(D11111_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D11087 ( .AN(D2177_Y), .B0(D11004_Y), .Y(D11087_Y),     .B1(D11081_Q));
KC_AOI21B_X1 D11086 ( .AN(D11060_Y), .B0(D11081_Q), .Y(D11086_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D11008 ( .AN(D11018_Y), .B0(D11004_Y), .Y(D11008_Y),     .B1(D10992_Q));
KC_AOI21B_X1 D10961 ( .AN(D10928_Y), .B0(D2227_Y), .Y(D10961_Y),     .B1(D1033_Q));
KC_AOI21B_X1 D10960 ( .AN(D10923_Y), .B0(D2227_Y), .Y(D10960_Y),     .B1(D10945_Q));
KC_AOI21B_X1 D10959 ( .AN(D10924_Y), .B0(D10945_Q), .Y(D10959_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D10958 ( .AN(D11359_Y), .B0(D2227_Y), .Y(D10958_Y),     .B1(D11391_Q));
KC_AOI21B_X1 D10957 ( .AN(D11362_Y), .B0(D2227_Y), .Y(D10957_Y),     .B1(D11393_Q));
KC_AOI21B_X1 D10893 ( .AN(D11281_Y), .B0(D2227_Y), .Y(D10893_Y),     .B1(D11336_Q));
KC_AOI21B_X1 D10659 ( .AN(D554_Y), .B0(D10649_Q), .Y(D10659_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D10658 ( .AN(D2207_Y), .B0(D2214_Q), .Y(D10658_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D10657 ( .AN(D10638_Y), .B0(D10776_Y), .Y(D10657_Y),     .B1(D10649_Q));
KC_AOI21B_X1 D10656 ( .AN(D10636_Y), .B0(D10652_Q), .Y(D10656_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D10655 ( .AN(D10637_Y), .B0(D10776_Y), .Y(D10655_Y),     .B1(D2214_Q));
KC_AOI21B_X1 D10654 ( .AN(D10639_Y), .B0(D10776_Y), .Y(D10654_Y),     .B1(D10651_Q));
KC_AOI21B_X1 D10628 ( .AN(D11097_Y), .B0(D11107_Q), .Y(D10628_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D10627 ( .AN(D10604_Y), .B0(D11004_Y), .Y(D10627_Y),     .B1(D10618_Q));
KC_AOI21B_X1 D10626 ( .AN(D11095_Y), .B0(D11004_Y), .Y(D10626_Y),     .B1(D11107_Q));
KC_AOI21B_X1 D10625 ( .AN(D10605_Y), .B0(D11004_Y), .Y(D10625_Y),     .B1(D1368_Q));
KC_AOI21B_X1 D10624 ( .AN(D10608_Y), .B0(D10618_Q), .Y(D10624_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D10623 ( .AN(D11094_Y), .B0(D1368_Q), .Y(D10623_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D10622 ( .AN(D1334_Y), .B0(D11004_Y), .Y(D10622_Y),     .B1(D10616_Q));
KC_AOI21B_X1 D10621 ( .AN(D10606_Y), .B0(D10616_Q), .Y(D10621_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D10620 ( .AN(D10609_Y), .B0(D10614_Q), .Y(D10620_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D10619 ( .AN(D10607_Y), .B0(D11004_Y), .Y(D10619_Y),     .B1(D10614_Q));
KC_AOI21B_X1 D10557 ( .AN(D11017_Y), .B0(D11053_Q), .Y(D10557_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D10556 ( .AN(D11016_Y), .B0(D11004_Y), .Y(D10556_Y),     .B1(D11053_Q));
KC_AOI21B_X1 D10440 ( .AN(D10444_Y), .B0(D10421_Q), .Y(D10440_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D10439 ( .AN(D2133_Y), .B0(D10355_Q), .Y(D10439_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D10438 ( .AN(D10405_Y), .B0(D2227_Y), .Y(D10438_Y),     .B1(D10355_Q));
KC_AOI21B_X1 D10437 ( .AN(D10404_Y), .B0(D1042_Q), .Y(D10437_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D10436 ( .AN(D10406_Y), .B0(D2227_Y), .Y(D10436_Y),     .B1(D1042_Q));
KC_AOI21B_X1 D10435 ( .AN(D2191_Y), .B0(D2227_Y), .Y(D10435_Y),     .B1(D10953_Q));
KC_AOI21B_X1 D10434 ( .AN(D2172_Y), .B0(D2227_Y), .Y(D10434_Y),     .B1(D10349_Q));
KC_AOI21B_X1 D10433 ( .AN(D10387_Y), .B0(D10349_Q), .Y(D10433_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D10432 ( .AN(D2134_Y), .B0(D2227_Y), .Y(D10432_Y),     .B1(D10421_Q));
KC_AOI21B_X1 D10046 ( .AN(D8910_Y), .B0(D7313_Y), .Y(D10046_Y),     .B1(D10049_Q));
KC_AOI21B_X1 D10030 ( .AN(D8848_Y), .B0(D2070_Y), .Y(D10030_Y),     .B1(D2166_Q));
KC_AOI21B_X1 D10029 ( .AN(D8912_Y), .B0(D2070_Y), .Y(D10029_Y),     .B1(D10009_Q));
KC_AOI21B_X1 D9940 ( .AN(D216_Y), .B0(D8697_Y), .Y(D9940_Y),     .B1(D9933_Y));
KC_AOI21B_X1 D9912 ( .AN(D9896_Y), .B0(D11004_Y), .Y(D9912_Y),     .B1(D1357_Q));
KC_AOI21B_X1 D9911 ( .AN(D9898_Y), .B0(D11004_Y), .Y(D9911_Y),     .B1(D9906_Q));
KC_AOI21B_X1 D9910 ( .AN(D9897_Y), .B0(D9906_Q), .Y(D9910_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D9848 ( .AN(D9824_Y), .B0(D11004_Y), .Y(D9848_Y),     .B1(D9835_Q));
KC_AOI21B_X1 D9847 ( .AN(D9825_Y), .B0(D11004_Y), .Y(D9847_Y),     .B1(D9837_Q));
KC_AOI21B_X1 D9846 ( .AN(D9826_Y), .B0(D9837_Q), .Y(D9846_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D9845 ( .AN(D9828_Y), .B0(D11004_Y), .Y(D9845_Y),     .B1(D1201_Q));
KC_AOI21B_X1 D9844 ( .AN(D9827_Y), .B0(D1201_Q), .Y(D9844_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D9843 ( .AN(D9829_Y), .B0(D9835_Q), .Y(D9843_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D9619 ( .AN(D858_Y), .B0(D9609_Q), .Y(D9619_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D9618 ( .AN(D9596_Y), .B0(D2227_Y), .Y(D9618_Y),     .B1(D9609_Q));
KC_AOI21B_X1 D9092 ( .AN(D9063_Y), .B0(D7494_Y), .Y(D9092_Y),     .B1(D387_Q));
KC_AOI21B_X1 D8820 ( .AN(D8763_Y), .B0(D233_Q), .Y(D8820_Y),     .B1(D8823_Q));
KC_AOI21B_X1 D8708 ( .AN(D7113_Y), .B0(D8704_Y), .Y(D8708_Y),     .B1(D7113_Y));
KC_AOI21B_X1 D8335 ( .AN(D6762_Y), .B0(D8344_Y), .Y(D8335_Y),     .B1(D11058_Y));
KC_AOI21B_X1 D8334 ( .AN(D6761_Y), .B0(D8344_Y), .Y(D8334_Y),     .B1(D10530_Y));
KC_AOI21B_X1 D8333 ( .AN(D6769_Y), .B0(D8344_Y), .Y(D8333_Y),     .B1(D2132_Y));
KC_AOI21B_X1 D8332 ( .AN(D6770_Y), .B0(D8344_Y), .Y(D8332_Y),     .B1(D10471_Y));
KC_AOI21B_X1 D8241 ( .AN(D8256_Y), .B0(D8223_Y), .Y(D8241_Y),     .B1(D8223_Y));
KC_AOI21B_X1 D8057 ( .AN(D610_Y), .B0(D1848_Y), .Y(D8057_Y),     .B1(D8033_Y));
KC_AOI21B_X1 D7658 ( .AN(D7618_Y), .B0(D393_Y), .Y(D7658_Y),     .B1(D7701_Y));
KC_AOI21B_X1 D7091 ( .AN(D1336_Y), .B0(D7044_Q), .Y(D7091_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D7090 ( .AN(D7069_Y), .B0(D1651_Y), .Y(D7090_Y),     .B1(D7044_Q));
KC_AOI21B_X1 D7089 ( .AN(D7064_Y), .B0(D1651_Y), .Y(D7089_Y),     .B1(D7080_Q));
KC_AOI21B_X1 D7088 ( .AN(D1335_Y), .B0(D1651_Y), .Y(D7088_Y),     .B1(D7075_Q));
KC_AOI21B_X1 D7087 ( .AN(D1333_Y), .B0(D7080_Q), .Y(D7087_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D7086 ( .AN(D1332_Y), .B0(D7075_Q), .Y(D7086_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D7062 ( .AN(D7035_Y), .B0(D7050_Q), .Y(D7062_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D7061 ( .AN(D7029_Y), .B0(D1651_Y), .Y(D7061_Y),     .B1(D7050_Q));
KC_AOI21B_X1 D7060 ( .AN(D1251_Y), .B0(D7049_Q), .Y(D7060_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D7059 ( .AN(D1253_Y), .B0(D1651_Y), .Y(D7059_Y),     .B1(D7049_Q));
KC_AOI21B_X1 D7058 ( .AN(D1250_Y), .B0(D7084_Q), .Y(D7058_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D7057 ( .AN(D7024_Y), .B0(D1651_Y), .Y(D7057_Y),     .B1(D7084_Q));
KC_AOI21B_X1 D6908 ( .AN(D6876_Y), .B0(D5454_Y), .Y(D6908_Y),     .B1(D6819_Q));
KC_AOI21B_X1 D6907 ( .AN(D6874_Y), .B0(D6903_Q), .Y(D6907_Y),     .B1(D5454_Y));
KC_AOI21B_X1 D6906 ( .AN(D6763_Y), .B0(D6903_Q), .Y(D6906_Y),     .B1(D6883_Y));
KC_AOI21B_X1 D6905 ( .AN(D977_Y), .B0(D6900_Q), .Y(D6905_Y),     .B1(D6883_Y));
KC_AOI21B_X1 D6904 ( .AN(D5447_Y), .B0(D5454_Y), .Y(D6904_Y),     .B1(D6900_Q));
KC_AOI21B_X1 D6343 ( .AN(D6312_Y), .B0(D428_Y), .Y(D6343_Y),     .B1(D6340_Y));
KC_AOI21B_X1 D6341 ( .AN(D6320_Y), .B0(D6176_Y), .Y(D6341_Y),     .B1(D6176_Y));
KC_AOI21B_X1 D6119 ( .AN(D6109_Y), .B0(D48_Y), .Y(D6119_Y),     .B1(D6116_Y));
KC_AOI21B_X1 D5934 ( .AN(D5933_Y), .B0(D5933_Y), .Y(D5934_Y),     .B1(D5933_Y));
KC_AOI21B_X1 D5639 ( .AN(D4075_Y), .B0(D1403_Q), .Y(D5639_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5638 ( .AN(D5620_Y), .B0(D1651_Y), .Y(D5638_Y),     .B1(D1403_Q));
KC_AOI21B_X1 D5637 ( .AN(D4074_Y), .B0(D1651_Y), .Y(D5637_Y),     .B1(D1355_Q));
KC_AOI21B_X1 D5636 ( .AN(D1331_Y), .B0(D1355_Q), .Y(D5636_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5635 ( .AN(D5616_Y), .B0(D1651_Y), .Y(D5635_Y),     .B1(D5628_Q));
KC_AOI21B_X1 D5634 ( .AN(D5617_Y), .B0(D5628_Q), .Y(D5634_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5614 ( .AN(D5595_Y), .B0(D1651_Y), .Y(D5614_Y),     .B1(D4051_Q));
KC_AOI21B_X1 D5613 ( .AN(D5598_Y), .B0(D1651_Y), .Y(D5613_Y),     .B1(D5610_Q));
KC_AOI21B_X1 D5612 ( .AN(D5594_Y), .B0(D4051_Q), .Y(D5612_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5611 ( .AN(D5591_Y), .B0(D5610_Q), .Y(D5611_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5541 ( .AN(D5503_Y), .B0(D1633_Q), .Y(D5541_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5539 ( .AN(D1083_Y), .B0(D1651_Y), .Y(D5539_Y),     .B1(D5533_Q));
KC_AOI21B_X1 D5538 ( .AN(D5504_Y), .B0(D1651_Y), .Y(D5538_Y),     .B1(D5532_Q));
KC_AOI21B_X1 D5537 ( .AN(D5517_Y), .B0(D5532_Q), .Y(D5537_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5536 ( .AN(D5505_Y), .B0(D1651_Y), .Y(D5536_Y),     .B1(D1633_Q));
KC_AOI21B_X1 D5535 ( .AN(D1081_Y), .B0(D5533_Q), .Y(D5535_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D5330 ( .AN(D5200_Y), .B0(D5323_Y), .Y(D5330_Y),     .B1(D663_Q));
KC_AOI21B_X1 D5329 ( .AN(D5287_Y), .B0(D663_Q), .Y(D5329_Y),     .B1(D921_Y));
KC_AOI21B_X1 D5328 ( .AN(D5284_Y), .B0(D794_Q), .Y(D5328_Y),     .B1(D5323_Y));
KC_AOI21B_X1 D5327 ( .AN(D5278_Y), .B0(D794_Q), .Y(D5327_Y),     .B1(D921_Y));
KC_AOI21B_X1 D5326 ( .AN(D5273_Y), .B0(D5323_Y), .Y(D5326_Y),     .B1(D791_Q));
KC_AOI21B_X1 D5325 ( .AN(D5270_Y), .B0(D791_Q), .Y(D5325_Y),     .B1(D921_Y));
KC_AOI21B_X1 D5324 ( .AN(D5262_Y), .B0(D5323_Y), .Y(D5324_Y),     .B1(D788_Q));
KC_AOI21B_X1 D5254 ( .AN(D5203_Y), .B0(D666_Q), .Y(D5254_Y),     .B1(D921_Y));
KC_AOI21B_X1 D5247 ( .AN(D5212_Y), .B0(D5240_Q), .Y(D5247_Y),     .B1(D921_Y));
KC_AOI21B_X1 D5246 ( .AN(D5211_Y), .B0(D5323_Y), .Y(D5246_Y),     .B1(D5240_Q));
KC_AOI21B_X1 D5245 ( .AN(D5209_Y), .B0(D5323_Y), .Y(D5245_Y),     .B1(D668_Q));
KC_AOI21B_X1 D5244 ( .AN(D5210_Y), .B0(D668_Q), .Y(D5244_Y),     .B1(D921_Y));
KC_AOI21B_X1 D5243 ( .AN(D5201_Y), .B0(D5323_Y), .Y(D5243_Y),     .B1(D666_Q));
KC_AOI21B_X1 D5242 ( .AN(D5205_Y), .B0(D5323_Y), .Y(D5242_Y),     .B1(D5235_Q));
KC_AOI21B_X1 D5241 ( .AN(D5204_Y), .B0(D5235_Q), .Y(D5241_Y),     .B1(D921_Y));
KC_AOI21B_X1 D4484 ( .AN(D7312_Y), .B0(D4434_Y), .Y(D4484_Y),     .B1(D4445_Y));
KC_AOI21B_X1 D4394 ( .AN(D4377_Y), .B0(D4391_Y), .Y(D4394_Y),     .B1(D4324_Y));
KC_AOI21B_X1 D4393 ( .AN(D7394_Y), .B0(D243_Y), .Y(D4393_Y),     .B1(D5876_Y));
KC_AOI21B_X1 D3979 ( .AN(D3957_Y), .B0(D3968_Q), .Y(D3979_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3978 ( .AN(D3956_Y), .B0(D5406_Y), .Y(D3978_Y),     .B1(D3975_Q));
KC_AOI21B_X1 D3977 ( .AN(D3952_Y), .B0(D3975_Q), .Y(D3977_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3976 ( .AN(D3953_Y), .B0(D3966_Q), .Y(D3976_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3950 ( .AN(D3919_Y), .B0(D3940_Q), .Y(D3950_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3949 ( .AN(D3920_Y), .B0(D5406_Y), .Y(D3949_Y),     .B1(D3940_Q));
KC_AOI21B_X1 D3948 ( .AN(D3913_Y), .B0(D5406_Y), .Y(D3948_Y),     .B1(D3939_Q));
KC_AOI21B_X1 D3947 ( .AN(D3914_Y), .B0(D3939_Q), .Y(D3947_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3946 ( .AN(D3899_Y), .B0(D3932_Q), .Y(D3946_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3945 ( .AN(D3894_Y), .B0(D5406_Y), .Y(D3945_Y),     .B1(D3932_Q));
KC_AOI21B_X1 D3885 ( .AN(D3886_Y), .B0(D3878_Q), .Y(D3885_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3884 ( .AN(D3845_Y), .B0(D5406_Y), .Y(D3884_Y),     .B1(D3878_Q));
KC_AOI21B_X1 D3883 ( .AN(D3840_Y), .B0(D5406_Y), .Y(D3883_Y),     .B1(D3876_Q));
KC_AOI21B_X1 D3882 ( .AN(D3834_Y), .B0(D3876_Q), .Y(D3882_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3828 ( .AN(D3785_Y), .B0(D3728_Q), .Y(D3828_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3827 ( .AN(D3778_Y), .B0(D5406_Y), .Y(D3827_Y),     .B1(D3796_Y));
KC_AOI21B_X1 D3826 ( .AN(D3791_Y), .B0(D5406_Y), .Y(D3826_Y),     .B1(D3814_Q));
KC_AOI21B_X1 D3825 ( .AN(D3784_Y), .B0(D3814_Q), .Y(D3825_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3824 ( .AN(D3781_Y), .B0(D3796_Y), .Y(D3824_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3823 ( .AN(D3768_Y), .B0(D5406_Y), .Y(D3823_Y),     .B1(D1498_Q));
KC_AOI21B_X1 D3822 ( .AN(D3774_Y), .B0(D5406_Y), .Y(D3822_Y),     .B1(D3803_Q));
KC_AOI21B_X1 D3821 ( .AN(D3775_Y), .B0(D3803_Q), .Y(D3821_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3820 ( .AN(D3766_Y), .B0(D1498_Q), .Y(D3820_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3749 ( .AN(D3712_Y), .B0(D5323_Y), .Y(D3749_Y),     .B1(D3737_Q));
KC_AOI21B_X1 D3748 ( .AN(D3705_Y), .B0(D3738_Q), .Y(D3748_Y),     .B1(D5406_Y));
KC_AOI21B_X1 D3747 ( .AN(D3706_Y), .B0(D3738_Q), .Y(D3747_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3746 ( .AN(D3704_Y), .B0(D3733_Q), .Y(D3746_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D3745 ( .AN(D3702_Y), .B0(D5406_Y), .Y(D3745_Y),     .B1(D3728_Q));
KC_AOI21B_X1 D3744 ( .AN(D3703_Y), .B0(D5406_Y), .Y(D3744_Y),     .B1(D3733_Q));
KC_AOI21B_X1 D3699 ( .AN(D3666_Y), .B0(D5323_Y), .Y(D3699_Y),     .B1(D1503_Q));
KC_AOI21B_X1 D3698 ( .AN(D3665_Y), .B0(D5323_Y), .Y(D3698_Y),     .B1(D3625_Q));
KC_AOI21B_X1 D3697 ( .AN(D3660_Y), .B0(D5323_Y), .Y(D3697_Y),     .B1(D3686_Q));
KC_AOI21B_X1 D3696 ( .AN(D3664_Y), .B0(D5323_Y), .Y(D3696_Y),     .B1(D3673_Q));
KC_AOI21B_X1 D3695 ( .AN(D3661_Y), .B0(D3686_Q), .Y(D3695_Y),     .B1(D921_Y));
KC_AOI21B_X1 D3694 ( .AN(D3663_Y), .B0(D3625_Q), .Y(D3694_Y),     .B1(D921_Y));
KC_AOI21B_X1 D3693 ( .AN(D3651_Y), .B0(D5323_Y), .Y(D3693_Y),     .B1(D3681_Q));
KC_AOI21B_X1 D3692 ( .AN(D3650_Y), .B0(D3681_Q), .Y(D3692_Y),     .B1(D921_Y));
KC_AOI21B_X1 D3691 ( .AN(D3659_Y), .B0(D3677_Q), .Y(D3691_Y),     .B1(D921_Y));
KC_AOI21B_X1 D3690 ( .AN(D3653_Y), .B0(D5323_Y), .Y(D3690_Y),     .B1(D3677_Q));
KC_AOI21B_X1 D3689 ( .AN(D3649_Y), .B0(D1503_Q), .Y(D3689_Y),     .B1(D921_Y));
KC_AOI21B_X1 D3688 ( .AN(D3652_Y), .B0(D5323_Y), .Y(D3688_Y),     .B1(D3675_Q));
KC_AOI21B_X1 D3687 ( .AN(D3654_Y), .B0(D3675_Q), .Y(D3687_Y),     .B1(D921_Y));
KC_AOI21B_X1 D3578 ( .AN(D4875_Y), .B0(D3067_Y), .Y(D3578_Y),     .B1(D3446_Y));
KC_AOI21B_X1 D3076 ( .AN(D2951_Y), .B0(D3070_Y), .Y(D3076_Y),     .B1(D1513_Y));
KC_AOI21B_X1 D3075 ( .AN(D4506_Y), .B0(D3046_Y), .Y(D3075_Y),     .B1(D3029_Y));
KC_AOI21B_X1 D2998 ( .AN(D2991_Y), .B0(D2989_Y), .Y(D2998_Y),     .B1(D2982_Y));
KC_AOI21B_X1 D2354 ( .AN(D12957_Y), .B0(D912_Q), .Y(D2354_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D2305 ( .AN(D2264_Y), .B0(D126_Q), .Y(D2305_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D2299 ( .AN(D11647_Y), .B0(D599_Q), .Y(D2299_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D2298 ( .AN(D11643_Y), .B0(D599_Q), .Y(D2298_Y),     .B1(D10776_Y));
KC_AOI21B_X1 D2226 ( .AN(D11019_Y), .B0(D2218_Q), .Y(D2226_Y),     .B1(D11004_Y));
KC_AOI21B_X1 D2225 ( .AN(D10635_Y), .B0(D10776_Y), .Y(D2225_Y),     .B1(D10653_Q));
KC_AOI21B_X1 D2224 ( .AN(D611_Y), .B0(D10653_Q), .Y(D2224_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D2165 ( .AN(D11020_Y), .B0(D11004_Y), .Y(D2165_Y),     .B1(D1314_Q));
KC_AOI21B_X1 D2164 ( .AN(D2178_Y), .B0(D1314_Q), .Y(D2164_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D2163 ( .AN(D8849_Y), .B0(D2070_Y), .Y(D2163_Y),     .B1(D9983_Q));
KC_AOI21B_X1 D2089 ( .AN(D2115_Y), .B0(D2227_Y), .Y(D2089_Y),     .B1(D9615_Q));
KC_AOI21B_X1 D2088 ( .AN(D2114_Y), .B0(D9615_Q), .Y(D2088_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D2087 ( .AN(D10317_Y), .B0(D2227_Y), .Y(D2087_Y),     .B1(D1024_Q));
KC_AOI21B_X1 D1938 ( .AN(D7639_Y), .B0(D7628_Y), .Y(D1938_Y),     .B1(D7572_Y));
KC_AOI21B_X1 D1790 ( .AN(D6246_Y), .B0(D6234_Y), .Y(D1790_Y),     .B1(D1765_Y));
KC_AOI21B_X1 D1789 ( .AN(D1686_Y), .B0(D1778_Q), .Y(D1789_Y),     .B1(D6883_Y));
KC_AOI21B_X1 D1788 ( .AN(D1687_Y), .B0(D6819_Q), .Y(D1788_Y),     .B1(D6883_Y));
KC_AOI21B_X1 D1650 ( .AN(D1079_Y), .B0(D5563_Q), .Y(D1650_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D1649 ( .AN(D5500_Y), .B0(D5563_Q), .Y(D1649_Y),     .B1(D1651_Y));
KC_AOI21B_X1 D1512 ( .AN(D3537_Y), .B0(D4916_Y), .Y(D1512_Y),     .B1(D4960_Y));
KC_AOI21B_X1 D1511 ( .AN(D3711_Y), .B0(D3737_Q), .Y(D1511_Y),     .B1(D921_Y));
KC_AOI21B_X1 D1510 ( .AN(D1409_Y), .B0(D5406_Y), .Y(D1510_Y),     .B1(D3968_Q));
KC_AOI21B_X1 D1509 ( .AN(D1408_Y), .B0(D3928_Q), .Y(D1509_Y),     .B1(D5409_Y));
KC_AOI21B_X1 D1508 ( .AN(D3955_Y), .B0(D5406_Y), .Y(D1508_Y),     .B1(D3928_Q));
KC_AOI21B_X1 D1507 ( .AN(D3954_Y), .B0(D5406_Y), .Y(D1507_Y),     .B1(D3966_Q));
KC_AOI21B_X1 D1372 ( .AN(D12605_Y), .B0(D2300_Y), .Y(D1372_Y),     .B1(D13150_Q));
KC_AOI21B_X1 D1371 ( .AN(D11093_Y), .B0(D11004_Y), .Y(D1371_Y),     .B1(D11108_Q));
KC_AOI21B_X1 D1370 ( .AN(D9895_Y), .B0(D1357_Q), .Y(D1370_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D1319 ( .AN(D1256_Y), .B0(D7055_Q), .Y(D1319_Y),     .B1(D6971_Y));
KC_AOI21B_X1 D1318 ( .AN(D1259_Y), .B0(D1651_Y), .Y(D1318_Y),     .B1(D7055_Q));
KC_AOI21B_X1 D1146 ( .AN(D2179_Y), .B0(D10992_Q), .Y(D1146_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D1145 ( .AN(D1088_Y), .B0(D13036_Q), .Y(D1145_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D1047 ( .AN(D12958_Y), .B0(D1039_Q), .Y(D1047_Y),     .B1(D11982_Y));
KC_AOI21B_X1 D1046 ( .AN(D2193_Y), .B0(D10953_Q), .Y(D1046_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D1045 ( .AN(D11367_Y), .B0(D1033_Q), .Y(D1045_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D923 ( .AN(D11283_Y), .B0(D908_Q), .Y(D923_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D922 ( .AN(D11370_Y), .B0(D11402_Q), .Y(D922_Y),     .B1(D11007_Y));
KC_AOI21B_X1 D811 ( .AN(D5261_Y), .B0(D788_Q), .Y(D811_Y),     .B1(D921_Y));
KC_AOI21B_X1 D604 ( .AN(D555_Y), .B0(D11127_Q), .Y(D604_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D603 ( .AN(D556_Y), .B0(D10651_Q), .Y(D603_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D602 ( .AN(D10640_Y), .B0(D10776_Y), .Y(D602_Y),     .B1(D10652_Q));
KC_AOI21B_X1 D601 ( .AN(D11121_Y), .B0(D2246_Q), .Y(D601_Y),     .B1(D10806_Y));
KC_AOI21B_X1 D600 ( .AN(D3662_Y), .B0(D3673_Q), .Y(D600_Y),     .B1(D921_Y));
KC_AOI21B_X1 D140 ( .AN(D11371_Y), .B0(D2227_Y), .Y(D140_Y),     .B1(D11402_Q));
KC_AOI21B_X1 D139 ( .AN(D11021_Y), .B0(D2218_Q), .Y(D139_Y),     .B1(D10516_Y));
KC_AOI21B_X1 D138 ( .AN(D9595_Y), .B0(D1024_Q), .Y(D138_Y),     .B1(D11007_Y));
KC_DFFHQ_X1 D13820 ( .Q(D13820_Q), .D(D2303_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D13819 ( .Q(D13819_Q), .D(D2303_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D13803 ( .Q(D13803_Q), .D(D12057_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D13802 ( .Q(D13802_Q), .D(D2303_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D13801 ( .Q(D13801_Q), .D(D12057_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D13800 ( .Q(D13800_Q), .D(D2302_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D13799 ( .Q(D13799_Q), .D(D12054_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D13798 ( .Q(D13798_Q), .D(D12054_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D13756 ( .Q(D13756_Q), .D(D12054_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D13150 ( .Q(D13150_Q), .D(D11586_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D13149 ( .Q(D13149_Q), .D(D12055_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D13148 ( .Q(D13148_Q), .D(D12054_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D13147 ( .Q(D13147_Q), .D(D11993_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D13146 ( .Q(D13146_Q), .D(D11993_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D13145 ( .Q(D13145_Q), .D(D11586_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D13144 ( .Q(D13144_Q), .D(D12055_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D13143 ( .Q(D13143_Q), .D(D12054_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D13120 ( .Q(D13120_Q), .D(D12055_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D13119 ( .Q(D13119_Q), .D(D2302_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D13118 ( .Q(D13118_Q), .D(D2302_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D13117 ( .Q(D13117_Q), .D(D2302_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D13116 ( .Q(D13116_Q), .D(D12055_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D13115 ( .Q(D13115_Q), .D(D12055_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D13114 ( .Q(D13114_Q), .D(D12055_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D16097 ( .Q(D16097_Q), .D(D12054_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D13096 ( .Q(D13096_Q), .D(D12057_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D13095 ( .Q(D13095_Q), .D(D12057_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D13088 ( .Q(D13088_Q), .D(D11993_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D13087 ( .Q(D13087_Q), .D(D12054_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D13086 ( .Q(D13086_Q), .D(D12054_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D13083 ( .Q(D13083_Q), .D(D2303_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D13082 ( .Q(D13082_Q), .D(D2303_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D13081 ( .Q(D13081_Q), .D(D11993_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D13080 ( .Q(D13080_Q), .D(D12057_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D13045 ( .Q(D13045_Q), .D(D11993_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D13044 ( .Q(D13044_Q), .D(D11993_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D13043 ( .Q(D13043_Q), .D(D2303_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D13042 ( .Q(D13042_Q), .D(D11995_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D13041 ( .Q(D13041_Q), .D(D11995_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D13040 ( .Q(D13040_Q), .D(D11384_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D13039 ( .Q(D13039_Q), .D(D11453_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D13038 ( .Q(D13038_Q), .D(D11384_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D13037 ( .Q(D13037_Q), .D(D1161_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D13036 ( .Q(D13036_Q), .D(D11453_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D13035 ( .Q(D13035_Q), .D(D11995_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D13034 ( .Q(D13034_Q), .D(D11453_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D13033 ( .Q(D13033_Q), .D(D1161_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D13032 ( .Q(D13032_Q), .D(D11453_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D13031 ( .Q(D13031_Q), .D(D1161_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D12987 ( .Q(D12987_Q), .D(D11851_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D12986 ( .Q(D12986_Q), .D(D11852_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D12985 ( .Q(D12985_Q), .D(D11852_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D12984 ( .Q(D12984_Q), .D(D11847_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D12983 ( .Q(D12983_Q), .D(D11847_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D12982 ( .Q(D12982_Q), .D(D11384_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D12981 ( .Q(D12981_Q), .D(D11384_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D12980 ( .Q(D12980_Q), .D(D11384_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D12979 ( .Q(D12979_Q), .D(D11995_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D12978 ( .Q(D12978_Q), .D(D11995_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D12977 ( .Q(D12977_Q), .D(D11384_Y), .CK(D112_QN));
KC_DFFHQ_X1 D12976 ( .Q(D12976_Q), .D(D1161_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D12913 ( .Q(D12913_Q), .D(D11846_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D12912 ( .Q(D12912_Q), .D(D11846_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D12620 ( .Q(D12620_Q), .D(D11968_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D12619 ( .Q(D12619_Q), .D(D12053_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D12618 ( .Q(D12618_Q), .D(D11968_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D12617 ( .Q(D12617_Q), .D(D11992_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D12615 ( .Q(D12615_Q), .D(D11966_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D12614 ( .Q(D12614_Q), .D(D12056_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D12613 ( .Q(D12613_Q), .D(D12056_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D12612 ( .Q(D12612_Q), .D(D11966_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D12611 ( .Q(D12611_Q), .D(D12056_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D12610 ( .Q(D12610_Q), .D(D11992_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D12609 ( .Q(D12609_Q), .D(D12053_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D12608 ( .Q(D12608_Q), .D(D11968_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D12607 ( .Q(D12607_Q), .D(D11992_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D12585 ( .Q(D12585_Q), .D(D11968_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D12584 ( .Q(D12584_Q), .D(D12056_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D12583 ( .Q(D12583_Q), .D(D12056_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D12582 ( .Q(D12582_Q), .D(D11968_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D12581 ( .Q(D12581_Q), .D(D11586_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D12580 ( .Q(D12580_Q), .D(D11968_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D12579 ( .Q(D12579_Q), .D(D12056_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D12578 ( .Q(D12578_Q), .D(D11968_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D12577 ( .Q(D12577_Q), .D(D11586_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D12576 ( .Q(D12576_Q), .D(D12056_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D12575 ( .Q(D12575_Q), .D(D11586_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D12574 ( .Q(D12574_Q), .D(D11586_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D12573 ( .Q(D12573_Q), .D(D11966_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D12572 ( .Q(D12572_Q), .D(D12053_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D12551 ( .Q(D12551_Q), .D(D12053_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D12550 ( .Q(D12550_Q), .D(D11992_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D12546 ( .Q(D12546_Q), .D(D11992_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D12545 ( .Q(D12545_Q), .D(D11994_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D12544 ( .Q(D12544_Q), .D(D11992_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D12543 ( .Q(D12543_Q), .D(D11994_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D12542 ( .Q(D12542_Q), .D(D12053_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D12541 ( .Q(D12541_Q), .D(D11966_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D12540 ( .Q(D12540_Q), .D(D11966_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D12539 ( .Q(D12539_Q), .D(D12053_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D12507 ( .Q(D12507_Q), .D(D11994_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D12506 ( .Q(D12506_Q), .D(D1161_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D12505 ( .Q(D12505_Q), .D(D11453_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D12504 ( .Q(D12504_Q), .D(D1004_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D12503 ( .Q(D12503_Q), .D(D1004_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D12502 ( .Q(D12502_Q), .D(D11995_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D12501 ( .Q(D12501_Q), .D(D1004_Y), .CK(D112_QN));
KC_DFFHQ_X1 D12500 ( .Q(D12500_Q), .D(D1161_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D12499 ( .Q(D12499_Q), .D(D11454_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D12498 ( .Q(D12498_Q), .D(D1004_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D12497 ( .Q(D12497_Q), .D(D11453_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D12496 ( .Q(D12496_Q), .D(D1161_Y), .CK(D112_QN));
KC_DFFHQ_X1 D12495 ( .Q(D12495_Q), .D(D1004_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D12494 ( .Q(D12494_Q), .D(D1004_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D12468 ( .Q(D12468_Q), .D(D11852_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D12467 ( .Q(D12467_Q), .D(D11852_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D12466 ( .Q(D12466_Q), .D(D11852_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D12465 ( .Q(D12465_Q), .D(D11852_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D12464 ( .Q(D12464_Q), .D(D11847_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D12463 ( .Q(D12463_Q), .D(D11847_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D12462 ( .Q(D12462_Q), .D(D11847_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D12461 ( .Q(D12461_Q), .D(D11847_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D12460 ( .Q(D12460_Q), .D(D11847_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D12459 ( .Q(D12459_Q), .D(D11847_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D12458 ( .Q(D12458_Q), .D(D1004_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D12457 ( .Q(D12457_Q), .D(D11384_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D12456 ( .Q(D12456_Q), .D(D11384_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D12455 ( .Q(D12455_Q), .D(D11454_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D12454 ( .Q(D12454_Q), .D(D11454_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D12453 ( .Q(D12453_Q), .D(D11995_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D12452 ( .Q(D12452_Q), .D(D1004_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D12451 ( .Q(D12451_Q), .D(D1161_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D12450 ( .Q(D12450_Q), .D(D11995_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D12449 ( .Q(D12449_Q), .D(D1004_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D12410 ( .Q(D12410_Q), .D(D11846_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D12409 ( .Q(D12409_Q), .D(D11846_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D12408 ( .Q(D12408_Q), .D(D11846_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D12407 ( .Q(D12407_Q), .D(D11852_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D12406 ( .Q(D12406_Q), .D(D11852_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D12405 ( .Q(D12405_Q), .D(D11846_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D12404 ( .Q(D12404_Q), .D(D11851_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D12403 ( .Q(D12403_Q), .D(D11851_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D12402 ( .Q(D12402_Q), .D(D11854_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D12401 ( .Q(D12401_Q), .D(D11846_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D12400 ( .Q(D12400_Q), .D(D11854_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D12399 ( .Q(D12399_Q), .D(D11846_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D12398 ( .Q(D12398_Q), .D(D11851_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D12397 ( .Q(D12397_Q), .D(D11851_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D12337 ( .Q(D12337_Q), .D(D11778_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D12336 ( .Q(D12336_Q), .D(D11778_Y), .CK(D660_QN));
KC_DFFHQ_X1 D12306 ( .Q(D12306_Q), .D(D11786_Y), .CK(D660_QN));
KC_DFFHQ_X1 D12270 ( .Q(D12270_Q), .D(D11785_Y), .CK(D660_QN));
KC_DFFHQ_X1 D12127 ( .Q(D12127_Q), .D(D11477_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D12122 ( .Q(D12122_Q), .D(D11967_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D12121 ( .Q(D12121_Q), .D(D11967_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D12120 ( .Q(D12120_Q), .D(D11534_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D12119 ( .Q(D12119_Q), .D(D11477_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D12117 ( .Q(D12117_Q), .D(D11477_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D12116 ( .Q(D12116_Q), .D(D11534_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D12096 ( .Q(D12096_Q), .D(D11967_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D12095 ( .Q(D12095_Q), .D(D11967_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D12094 ( .Q(D12094_Q), .D(D11967_Y), .CK(D12085_QN));
KC_DFFHQ_X1 D12093 ( .Q(D12093_Q), .D(D11967_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D12092 ( .Q(D12092_Q), .D(D11477_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D12091 ( .Q(D12091_Q), .D(D11534_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D12090 ( .Q(D12090_Q), .D(D11534_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D12089 ( .Q(D12089_Q), .D(D11534_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D12088 ( .Q(D12088_Q), .D(D11967_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D12087 ( .Q(D12087_Q), .D(D11967_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D12086 ( .Q(D12086_Q), .D(D11967_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D12058 ( .Q(D12058_Q), .D(D12053_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D12046 ( .Q(D12046_Q), .D(D11477_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D12045 ( .Q(D12045_Q), .D(D12056_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D12044 ( .Q(D12044_Q), .D(D11992_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D12043 ( .Q(D12043_Q), .D(D12005_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D12042 ( .Q(D12042_Q), .D(D12029_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D11980 ( .Q(D11980_Q), .D(D11383_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D11979 ( .Q(D11979_Q), .D(D11382_Y), .CK(D112_QN));
KC_DFFHQ_X1 D11978 ( .Q(D11978_Q), .D(D11383_Y), .CK(D112_QN));
KC_DFFHQ_X1 D11977 ( .Q(D11977_Q), .D(D11382_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D11976 ( .Q(D11976_Q), .D(D11383_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D11975 ( .Q(D11975_Q), .D(D11382_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D11974 ( .Q(D11974_Q), .D(D11382_Y), .CK(D1118_QN));
KC_DFFHQ_X1 D11973 ( .Q(D11973_Q), .D(D11383_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D11972 ( .Q(D11972_Q), .D(D11383_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D11971 ( .Q(D11971_Q), .D(D11382_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D11926 ( .Q(D11926_Q), .D(D11848_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D11925 ( .Q(D11925_Q), .D(D11849_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D11924 ( .Q(D11924_Q), .D(D11849_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D11923 ( .Q(D11923_Q), .D(D11383_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D11922 ( .Q(D11922_Q), .D(D11382_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D11921 ( .Q(D11921_Q), .D(D11382_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D11920 ( .Q(D11920_Q), .D(D11383_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D11919 ( .Q(D11919_Q), .D(D11382_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D11918 ( .Q(D11918_Q), .D(D11383_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D11917 ( .Q(D11917_Q), .D(D11382_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D11871 ( .Q(D11871_Q), .D(D11848_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D11870 ( .Q(D11870_Q), .D(D11908_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D11869 ( .Q(D11869_Q), .D(D11848_Y), .CK(D11912_QN));
KC_DFFHQ_X1 D11868 ( .Q(D11868_Q), .D(D11908_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D11867 ( .Q(D11867_Q), .D(D11848_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D11866 ( .Q(D11866_Q), .D(D11908_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D11865 ( .Q(D11865_Q), .D(D11848_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D11864 ( .Q(D11864_Q), .D(D11908_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D11863 ( .Q(D11863_Q), .D(D11848_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D11862 ( .Q(D11862_Q), .D(D11908_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D11861 ( .Q(D11861_Q), .D(D11848_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D11860 ( .Q(D11860_Q), .D(D11908_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D11859 ( .Q(D11859_Q), .D(D11300_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11858 ( .Q(D11858_Q), .D(D11908_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D11857 ( .Q(D11857_Q), .D(D11848_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D11856 ( .Q(D11856_Q), .D(D11908_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D11855 ( .Q(D11855_Q), .D(D11848_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D11804 ( .Q(D11804_Q), .D(D11783_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D11803 ( .Q(D11803_Q), .D(D11785_Y), .CK(D718_QN));
KC_DFFHQ_X1 D11802 ( .Q(D11802_Q), .D(D2283_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D11801 ( .Q(D11801_Q), .D(D11783_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D11800 ( .Q(D11800_Q), .D(D2283_Y), .CK(D661_QN));
KC_DFFHQ_X1 D11799 ( .Q(D11799_Q), .D(D11783_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D11798 ( .Q(D11798_Q), .D(D11783_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D11797 ( .Q(D11797_Q), .D(D11778_Y), .CK(D661_QN));
KC_DFFHQ_X1 D11796 ( .Q(D11796_Q), .D(D11783_Y), .CK(D718_QN));
KC_DFFHQ_X1 D11795 ( .Q(D11795_Q), .D(D2283_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D11794 ( .Q(D11794_Q), .D(D2283_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D11793 ( .Q(D11793_Q), .D(D2283_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D11792 ( .Q(D11792_Q), .D(D11779_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D11791 ( .Q(D11791_Q), .D(D2283_Y), .CK(D718_QN));
KC_DFFHQ_X1 D11790 ( .Q(D11790_Q), .D(D11778_Y), .CK(D718_QN));
KC_DFFHQ_X1 D11789 ( .Q(D11789_Q), .D(D11779_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D11788 ( .Q(D11788_Q), .D(D11779_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D11735 ( .Q(D11735_Q), .D(D11787_Y), .CK(D718_QN));
KC_DFFHQ_X1 D11734 ( .Q(D11734_Q), .D(D11787_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D11733 ( .Q(D11733_Q), .D(D11786_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D11732 ( .Q(D11732_Q), .D(D11785_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D11731 ( .Q(D11731_Q), .D(D11785_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D11726 ( .Q(D11726_Q), .D(D11786_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D11725 ( .Q(D11725_Q), .D(D11786_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D11724 ( .Q(D11724_Q), .D(D11787_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D11723 ( .Q(D11723_Q), .D(D11787_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D11722 ( .Q(D11722_Q), .D(D11787_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D11721 ( .Q(D11721_Q), .D(D11785_Y), .CK(D661_QN));
KC_DFFHQ_X1 D11720 ( .Q(D11720_Q), .D(D11786_Y), .CK(D718_QN));
KC_DFFHQ_X1 D11719 ( .Q(D11719_Q), .D(D11783_Y), .CK(D660_QN));
KC_DFFHQ_X1 D11718 ( .Q(D11718_Q), .D(D11785_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D11717 ( .Q(D11717_Q), .D(D11784_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D11716 ( .Q(D11716_Q), .D(D11783_Y), .CK(D661_QN));
KC_DFFHQ_X1 D11715 ( .Q(D11715_Q), .D(D11785_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D11662 ( .Q(D11662_Q), .D(D11779_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D11661 ( .Q(D11661_Q), .D(D11787_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D11659 ( .Q(D11659_Q), .D(D11779_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D11658 ( .Q(D11658_Q), .D(D11787_Y), .CK(D661_QN));
KC_DFFHQ_X1 D11656 ( .Q(D11656_Q), .D(D11787_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D11585 ( .Q(D11585_Q), .D(D11534_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D11584 ( .Q(D11584_Q), .D(D11534_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D11543 ( .Q(D11543_Q), .D(D11508_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D11542 ( .Q(D11542_Q), .D(D11487_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D11541 ( .Q(D11541_Q), .D(D11507_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D11539 ( .Q(D11539_Q), .D(D1176_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D11538 ( .Q(D11538_Q), .D(D11512_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D11537 ( .Q(D11537_Q), .D(D11511_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D11475 ( .Q(D11475_Q), .D(D11437_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D11474 ( .Q(D11474_Q), .D(D10503_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D11473 ( .Q(D11473_Q), .D(D1003_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D11472 ( .Q(D11472_Q), .D(D1003_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D11471 ( .Q(D11471_Q), .D(D1003_Y), .CK(D899_QN));
KC_DFFHQ_X1 D11470 ( .Q(D11470_Q), .D(D10503_Y), .CK(D901_QN));
KC_DFFHQ_X1 D11469 ( .Q(D11469_Q), .D(D11430_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D11468 ( .Q(D11468_Q), .D(D11420_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D11467 ( .Q(D11467_Q), .D(D1003_Y), .CK(D901_QN));
KC_DFFHQ_X1 D11466 ( .Q(D11466_Q), .D(D11424_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D11402 ( .Q(D11402_Q), .D(D10415_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D11401 ( .Q(D11401_Q), .D(D10415_Y), .CK(D897_QN));
KC_DFFHQ_X1 D11400 ( .Q(D11400_Q), .D(D10414_Y), .CK(D897_QN));
KC_DFFHQ_X1 D11399 ( .Q(D11399_Q), .D(D10503_Y), .CK(D897_QN));
KC_DFFHQ_X1 D11398 ( .Q(D11398_Q), .D(D10503_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D11397 ( .Q(D11397_Q), .D(D10502_Y), .CK(D897_QN));
KC_DFFHQ_X1 D11396 ( .Q(D11396_Q), .D(D1003_Y), .CK(D897_QN));
KC_DFFHQ_X1 D11395 ( .Q(D11395_Q), .D(D10502_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D11394 ( .Q(D11394_Q), .D(D1003_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D11393 ( .Q(D11393_Q), .D(D10503_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D11392 ( .Q(D11392_Q), .D(D11357_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D11391 ( .Q(D11391_Q), .D(D10502_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D11390 ( .Q(D11390_Q), .D(D11373_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D11389 ( .Q(D11389_Q), .D(D11435_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D11388 ( .Q(D11388_Q), .D(D1003_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D11342 ( .Q(D11342_Q), .D(D11299_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11341 ( .Q(D11341_Q), .D(D11294_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11340 ( .Q(D11340_Q), .D(D11286_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11339 ( .Q(D11339_Q), .D(D1113_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D11338 ( .Q(D11338_Q), .D(D1113_Y), .CK(D897_QN));
KC_DFFHQ_X1 D11337 ( .Q(D11337_Q), .D(D1007_Y), .CK(D897_QN));
KC_DFFHQ_X1 D11336 ( .Q(D11336_Q), .D(D1007_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D11335 ( .Q(D11335_Q), .D(D1007_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D11330 ( .Q(D11330_Q), .D(D10415_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D11329 ( .Q(D11329_Q), .D(D868_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11328 ( .Q(D11328_Q), .D(D2233_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11327 ( .Q(D11327_Q), .D(D11188_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D11326 ( .Q(D11326_Q), .D(D11292_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11325 ( .Q(D11325_Q), .D(D11285_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11275 ( .Q(D11275_Q), .D(D11252_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D11274 ( .Q(D11274_Q), .D(D11246_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D11273 ( .Q(D11273_Q), .D(D11246_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D11272 ( .Q(D11272_Q), .D(D11252_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D11271 ( .Q(D11271_Q), .D(D11254_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D11270 ( .Q(D11270_Q), .D(D11252_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D11269 ( .Q(D11269_Q), .D(D11246_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D11268 ( .Q(D11268_Q), .D(D11784_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D11267 ( .Q(D11267_Q), .D(D11252_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D11266 ( .Q(D11266_Q), .D(D11246_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D11265 ( .Q(D11265_Q), .D(D11202_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11264 ( .Q(D11264_Q), .D(D11230_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11263 ( .Q(D11263_Q), .D(D11199_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D11262 ( .Q(D11262_Q), .D(D11201_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11261 ( .Q(D11261_Q), .D(D11197_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11260 ( .Q(D11260_Q), .D(D11233_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D11187 ( .Q(D11187_Q), .D(D11253_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D11182 ( .Q(D11182_Q), .D(D11253_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D11181 ( .Q(D11181_Q), .D(D11253_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D11180 ( .Q(D11180_Q), .D(D11253_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D11179 ( .Q(D11179_Q), .D(D11784_Y), .CK(D661_QN));
KC_DFFHQ_X1 D11178 ( .Q(D11178_Q), .D(D11246_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D11177 ( .Q(D11177_Q), .D(D11252_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D11176 ( .Q(D11176_Q), .D(D11246_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D11175 ( .Q(D11175_Q), .D(D11784_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D11128 ( .Q(D11128_Q), .D(D11246_Y), .CK(D588_QN));
KC_DFFHQ_X1 D11127 ( .Q(D11127_Q), .D(D11252_Y), .CK(D588_QN));
KC_DFFHQ_X1 D11126 ( .Q(D11126_Q), .D(D11246_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D11125 ( .Q(D11125_Q), .D(D11246_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D11110 ( .Q(D11110_Q), .D(D10563_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D11109 ( .Q(D11109_Q), .D(D10563_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D11108 ( .Q(D11108_Q), .D(D10562_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D11107 ( .Q(D11107_Q), .D(D10563_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D11106 ( .Q(D11106_Q), .D(D10562_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D11105 ( .Q(D11105_Q), .D(D10562_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D11104 ( .Q(D11104_Q), .D(D1955_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D11085 ( .Q(D11085_Q), .D(D10563_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D11084 ( .Q(D11084_Q), .D(D10562_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D11083 ( .Q(D11083_Q), .D(D10563_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D11082 ( .Q(D11082_Q), .D(D10562_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D11081 ( .Q(D11081_Q), .D(D9780_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D11080 ( .Q(D11080_Q), .D(D9780_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D11079 ( .Q(D11079_Q), .D(D9780_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D11078 ( .Q(D11078_Q), .D(D9780_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D11077 ( .Q(D11077_Q), .D(D9780_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D11076 ( .Q(D11076_Q), .D(D10562_Y), .CK(D111_QN));
KC_DFFHQ_X1 D11075 ( .Q(D11075_Q), .D(D10563_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D11074 ( .Q(D11074_Q), .D(D10563_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D11073 ( .Q(D11073_Q), .D(D10563_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D11056 ( .Q(D11056_Q), .D(D10496_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D11053 ( .Q(D11053_Q), .D(D10496_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D11035 ( .Q(D11035_Q), .D(D10492_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D11034 ( .Q(D11034_Q), .D(D10542_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D11033 ( .Q(D11033_Q), .D(D10542_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D11031 ( .Q(D11031_Q), .D(D10498_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D11030 ( .Q(D11030_Q), .D(D10492_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D11027 ( .Q(D11027_Q), .D(D10496_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D11026 ( .Q(D11026_Q), .D(D10496_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D11002 ( .Q(D11002_Q), .D(D10502_Y), .CK(D899_QN));
KC_DFFHQ_X1 D11001 ( .Q(D11001_Q), .D(D10507_Y), .CK(D899_QN));
KC_DFFHQ_X1 D11000 ( .Q(D11000_Q), .D(D10502_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10999 ( .Q(D10999_Q), .D(D10503_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10998 ( .Q(D10998_Q), .D(D10507_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10997 ( .Q(D10997_Q), .D(D10507_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D10996 ( .Q(D10996_Q), .D(D10502_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D10995 ( .Q(D10995_Q), .D(D10502_Y), .CK(D901_QN));
KC_DFFHQ_X1 D10994 ( .Q(D10994_Q), .D(D10981_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D10993 ( .Q(D10993_Q), .D(D1003_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10992 ( .Q(D10992_Q), .D(D10498_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D10991 ( .Q(D10991_Q), .D(D10492_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D10956 ( .Q(D10956_Q), .D(D9777_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D10955 ( .Q(D10955_Q), .D(D10414_Y), .CK(D899_QN));
KC_DFFHQ_X1 D10954 ( .Q(D10954_Q), .D(D1113_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D10953 ( .Q(D10953_Q), .D(D9777_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D10952 ( .Q(D10952_Q), .D(D10507_Y), .CK(D897_QN));
KC_DFFHQ_X1 D10951 ( .Q(D10951_Q), .D(D1113_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D10950 ( .Q(D10950_Q), .D(D10414_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10949 ( .Q(D10949_Q), .D(D9777_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D10948 ( .Q(D10948_Q), .D(D10414_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D10947 ( .Q(D10947_Q), .D(D10507_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D10946 ( .Q(D10946_Q), .D(D9795_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D10945 ( .Q(D10945_Q), .D(D10507_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D10944 ( .Q(D10944_Q), .D(D10414_Y), .CK(D901_QN));
KC_DFFHQ_X1 D10943 ( .Q(D10943_Q), .D(D10507_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D10942 ( .Q(D10942_Q), .D(D10414_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D10941 ( .Q(D10941_Q), .D(D10507_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D10940 ( .Q(D10940_Q), .D(D10502_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D10892 ( .Q(D10892_Q), .D(D1113_Y), .CK(D899_QN));
KC_DFFHQ_X1 D10891 ( .Q(D10891_Q), .D(D1113_Y), .CK(D901_QN));
KC_DFFHQ_X1 D10890 ( .Q(D10890_Q), .D(D10415_Y), .CK(D899_QN));
KC_DFFHQ_X1 D10889 ( .Q(D10889_Q), .D(D10415_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D10888 ( .Q(D10888_Q), .D(D10415_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D10887 ( .Q(D10887_Q), .D(D1007_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D10886 ( .Q(D10886_Q), .D(D1007_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10885 ( .Q(D10885_Q), .D(D10873_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D10884 ( .Q(D10884_Q), .D(D1007_Y), .CK(D899_QN));
KC_DFFHQ_X1 D10883 ( .Q(D10883_Q), .D(D1113_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D10882 ( .Q(D10882_Q), .D(D10415_Y), .CK(D901_QN));
KC_DFFHQ_X1 D10881 ( .Q(D10881_Q), .D(D1113_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10880 ( .Q(D10880_Q), .D(D10415_Y), .CK(D10877_QN));
KC_DFFHQ_X1 D10802 ( .Q(D10802_Q), .D(D10823_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D10801 ( .Q(D10801_Q), .D(D10823_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D10800 ( .Q(D10800_Q), .D(D10823_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D10793 ( .Q(D10793_Q), .D(D10739_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D10792 ( .Q(D10792_Q), .D(D11193_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D10791 ( .Q(D10791_Q), .D(D10731_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D10790 ( .Q(D10790_Q), .D(D2203_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D10789 ( .Q(D10789_Q), .D(D10740_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D10724 ( .Q(D10724_Q), .D(D10783_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D10723 ( .Q(D10723_Q), .D(D10824_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D10722 ( .Q(D10722_Q), .D(D10783_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D10721 ( .Q(D10721_Q), .D(D10783_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D10720 ( .Q(D10720_Q), .D(D10824_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D10719 ( .Q(D10719_Q), .D(D10824_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D10718 ( .Q(D10718_Q), .D(D10783_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D10717 ( .Q(D10717_Q), .D(D10783_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D10716 ( .Q(D10716_Q), .D(D10824_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D10715 ( .Q(D10715_Q), .D(D11254_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D10714 ( .Q(D10714_Q), .D(D10824_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D10713 ( .Q(D10713_Q), .D(D834_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D10712 ( .Q(D10712_Q), .D(D834_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D10711 ( .Q(D10711_Q), .D(D10823_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D10710 ( .Q(D10710_Q), .D(D10823_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D10709 ( .Q(D10709_Q), .D(D834_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D10708 ( .Q(D10708_Q), .D(D834_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D10653 ( .Q(D10653_Q), .D(D10783_Y), .CK(D588_QN));
KC_DFFHQ_X1 D10652 ( .Q(D10652_Q), .D(D11254_Y), .CK(D588_QN));
KC_DFFHQ_X1 D10651 ( .Q(D10651_Q), .D(D10824_Y), .CK(D588_QN));
KC_DFFHQ_X1 D10650 ( .Q(D10650_Q), .D(D11254_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D10649 ( .Q(D10649_Q), .D(D10823_Y), .CK(D588_QN));
KC_DFFHQ_X1 D10632 ( .Q(D10632_Q), .D(D11252_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D10631 ( .Q(D10631_Q), .D(D834_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D10630 ( .Q(D10630_Q), .D(D834_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D10618 ( .Q(D10618_Q), .D(D9832_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D10617 ( .Q(D10617_Q), .D(D8628_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D10616 ( .Q(D10616_Q), .D(D8628_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D10615 ( .Q(D10615_Q), .D(D9832_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D10614 ( .Q(D10614_Q), .D(D8626_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D10613 ( .Q(D10613_Q), .D(D8628_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D10612 ( .Q(D10612_Q), .D(D8626_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D10611 ( .Q(D10611_Q), .D(D9832_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D10610 ( .Q(D10610_Q), .D(D8628_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D10603 ( .Q(D10603_Q), .D(D1955_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D10602 ( .Q(D10602_Q), .D(D10562_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D10601 ( .Q(D10601_Q), .D(D1955_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D10600 ( .Q(D10600_Q), .D(D1955_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D10599 ( .Q(D10599_Q), .D(D1955_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D10598 ( .Q(D10598_Q), .D(D1955_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D10597 ( .Q(D10597_Q), .D(D1955_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D10596 ( .Q(D10596_Q), .D(D8626_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D10595 ( .Q(D10595_Q), .D(D8626_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D10594 ( .Q(D10594_Q), .D(D8626_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D10555 ( .Q(D10555_Q), .D(D10496_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D10554 ( .Q(D10554_Q), .D(D9780_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D10553 ( .Q(D10553_Q), .D(D10498_Y), .CK(D111_QN));
KC_DFFHQ_X1 D10552 ( .Q(D10552_Q), .D(D10496_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D10551 ( .Q(D10551_Q), .D(D9780_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D10550 ( .Q(D10550_Q), .D(D10496_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D10549 ( .Q(D10549_Q), .D(D10542_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D10548 ( .Q(D10548_Q), .D(D10542_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D10547 ( .Q(D10547_Q), .D(D10492_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D10546 ( .Q(D10546_Q), .D(D10498_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D10545 ( .Q(D10545_Q), .D(D10492_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D10544 ( .Q(D10544_Q), .D(D10542_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D10515 ( .Q(D10515_Q), .D(D10517_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D10513 ( .Q(D10513_Q), .D(D10491_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D10512 ( .Q(D10512_Q), .D(D10492_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D10511 ( .Q(D10511_Q), .D(D10498_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D10510 ( .Q(D10510_Q), .D(D10498_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D10509 ( .Q(D10509_Q), .D(D10490_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D10508 ( .Q(D10508_Q), .D(D10482_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D10431 ( .Q(D10431_Q), .D(D9795_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D10430 ( .Q(D10430_Q), .D(D9795_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D10429 ( .Q(D10429_Q), .D(D10873_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D10428 ( .Q(D10428_Q), .D(D10873_Y), .CK(D900_QN));
KC_DFFHQ_X1 D10427 ( .Q(D10427_Q), .D(D9696_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D10426 ( .Q(D10426_Q), .D(D9696_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D10425 ( .Q(D10425_Q), .D(D9696_Y), .CK(D900_QN));
KC_DFFHQ_X1 D10424 ( .Q(D10424_Q), .D(D9777_Y), .CK(D900_QN));
KC_DFFHQ_X1 D10423 ( .Q(D10423_Q), .D(D9795_Y), .CK(D900_QN));
KC_DFFHQ_X1 D10422 ( .Q(D10422_Q), .D(D9777_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D10421 ( .Q(D10421_Q), .D(D9795_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D10420 ( .Q(D10420_Q), .D(D10873_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D10419 ( .Q(D10419_Q), .D(D9696_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D10418 ( .Q(D10418_Q), .D(D9777_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D10417 ( .Q(D10417_Q), .D(D9795_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D10355 ( .Q(D10355_Q), .D(D10873_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D10354 ( .Q(D10354_Q), .D(D9698_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D10353 ( .Q(D10353_Q), .D(D9698_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D10352 ( .Q(D10352_Q), .D(D10873_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D10351 ( .Q(D10351_Q), .D(D9702_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D10350 ( .Q(D10350_Q), .D(D9697_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D10349 ( .Q(D10349_Q), .D(D9698_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D10348 ( .Q(D10348_Q), .D(D9702_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D10347 ( .Q(D10347_Q), .D(D9697_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D10234 ( .Q(D10234_Q), .D(D10783_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D10185 ( .Q(D10185_Q), .D(D10783_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D10184 ( .Q(D10184_Q), .D(D10824_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D10183 ( .Q(D10183_Q), .D(D10783_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D9909 ( .Q(D9909_Q), .D(D8583_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D9908 ( .Q(D9908_Q), .D(D8585_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D9906 ( .Q(D9906_Q), .D(D8583_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D9905 ( .Q(D9905_Q), .D(D8583_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D9903 ( .Q(D9903_Q), .D(D8583_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D9892 ( .Q(D9892_Q), .D(D9833_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D9890 ( .Q(D9890_Q), .D(D8572_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D9889 ( .Q(D9889_Q), .D(D8572_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D9888 ( .Q(D9888_Q), .D(D9832_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D9887 ( .Q(D9887_Q), .D(D8628_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D9886 ( .Q(D9886_Q), .D(D9832_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D9885 ( .Q(D9885_Q), .D(D8628_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D9884 ( .Q(D9884_Q), .D(D8626_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D9883 ( .Q(D9883_Q), .D(D8628_Y), .CK(D111_QN));
KC_DFFHQ_X1 D9882 ( .Q(D9882_Q), .D(D9832_Y), .CK(D111_QN));
KC_DFFHQ_X1 D9881 ( .Q(D9881_Q), .D(D9832_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D9880 ( .Q(D9880_Q), .D(D8628_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D9879 ( .Q(D9879_Q), .D(D9832_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D9878 ( .Q(D9878_Q), .D(D9832_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D9877 ( .Q(D9877_Q), .D(D8628_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D9876 ( .Q(D9876_Q), .D(D8585_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D9842 ( .Q(D9842_Q), .D(D8573_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D9841 ( .Q(D9841_Q), .D(D9833_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D9840 ( .Q(D9840_Q), .D(D9833_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D9839 ( .Q(D9839_Q), .D(D2031_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D9838 ( .Q(D9838_Q), .D(D8572_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D9837 ( .Q(D9837_Q), .D(D8573_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D9836 ( .Q(D9836_Q), .D(D8572_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D9835 ( .Q(D9835_Q), .D(D8572_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D9834 ( .Q(D9834_Q), .D(D9833_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D9793 ( .Q(D9793_Q), .D(D9757_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D9792 ( .Q(D9792_Q), .D(D9763_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D9791 ( .Q(D9791_Q), .D(D9796_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D9790 ( .Q(D9790_Q), .D(D9762_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D9789 ( .Q(D9789_Q), .D(D1097_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D9788 ( .Q(D9788_Q), .D(D2037_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D9787 ( .Q(D9787_Q), .D(D2034_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D9786 ( .Q(D9786_Q), .D(D9685_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D9785 ( .Q(D9785_Q), .D(D1100_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D9784 ( .Q(D9784_Q), .D(D1099_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D9717 ( .Q(D9717_Q), .D(D9697_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D9714 ( .Q(D9714_Q), .D(D9697_Y), .CK(D900_QN));
KC_DFFHQ_X1 D9712 ( .Q(D9712_Q), .D(D9702_Y), .CK(D900_QN));
KC_DFFHQ_X1 D9711 ( .Q(D9711_Q), .D(D9695_Y), .CK(D900_QN));
KC_DFFHQ_X1 D9710 ( .Q(D9710_Q), .D(D9698_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D9709 ( .Q(D9709_Q), .D(D9698_Y), .CK(D898_QN));
KC_DFFHQ_X1 D9708 ( .Q(D9708_Q), .D(D9697_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D9707 ( .Q(D9707_Q), .D(D9696_Y), .CK(D898_QN));
KC_DFFHQ_X1 D9706 ( .Q(D9706_Q), .D(D9695_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D9705 ( .Q(D9705_Q), .D(D9697_Y), .CK(D898_QN));
KC_DFFHQ_X1 D9704 ( .Q(D9704_Q), .D(D9723_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D9703 ( .Q(D9703_Q), .D(D9695_Y), .CK(D898_QN));
KC_DFFHQ_X1 D9615 ( .Q(D9615_Q), .D(D9702_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D9614 ( .Q(D9614_Q), .D(D9695_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D9613 ( .Q(D9613_Q), .D(D9702_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D9612 ( .Q(D9612_Q), .D(D9702_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D9611 ( .Q(D9611_Q), .D(D9698_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D9610 ( .Q(D9610_Q), .D(D9697_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D9609 ( .Q(D9609_Q), .D(D9695_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D9608 ( .Q(D9608_Q), .D(D9695_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D9607 ( .Q(D9607_Q), .D(D9697_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D9606 ( .Q(D9606_Q), .D(D9698_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D8658 ( .Q(D8658_Q), .D(D8584_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D8657 ( .Q(D8657_Q), .D(D8629_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D8656 ( .Q(D8656_Q), .D(D8583_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D8655 ( .Q(D8655_Q), .D(D8627_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D8654 ( .Q(D8654_Q), .D(D8627_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D8653 ( .Q(D8653_Q), .D(D8581_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D8652 ( .Q(D8652_Q), .D(D8629_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D8651 ( .Q(D8651_Q), .D(D8629_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D8650 ( .Q(D8650_Q), .D(D8627_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D8643 ( .Q(D8643_Q), .D(D8585_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D8642 ( .Q(D8642_Q), .D(D8581_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D8641 ( .Q(D8641_Q), .D(D8584_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D8640 ( .Q(D8640_Q), .D(D8585_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D8639 ( .Q(D8639_Q), .D(D8583_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D8638 ( .Q(D8638_Q), .D(D8629_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D8637 ( .Q(D8637_Q), .D(D8585_Y), .CK(D111_QN));
KC_DFFHQ_X1 D8636 ( .Q(D8636_Q), .D(D8629_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D8635 ( .Q(D8635_Q), .D(D8583_Y), .CK(D111_QN));
KC_DFFHQ_X1 D8634 ( .Q(D8634_Q), .D(D8584_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D8633 ( .Q(D8633_Q), .D(D8627_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D8632 ( .Q(D8632_Q), .D(D8583_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D8631 ( .Q(D8631_Q), .D(D8581_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D8630 ( .Q(D8630_Q), .D(D8627_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D8595 ( .Q(D8595_Q), .D(D8566_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D8594 ( .Q(D8594_Q), .D(D8565_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8593 ( .Q(D8593_Q), .D(D8573_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D8591 ( .Q(D8591_Q), .D(D8573_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D8589 ( .Q(D8589_Q), .D(D8557_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8588 ( .Q(D8588_Q), .D(D8573_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D8549 ( .Q(D8549_Q), .D(D1096_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D8548 ( .Q(D8548_Q), .D(D1098_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8547 ( .Q(D8547_Q), .D(D8509_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8546 ( .Q(D8546_Q), .D(D8552_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8545 ( .Q(D8545_Q), .D(D8516_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8544 ( .Q(D8544_Q), .D(D1103_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8543 ( .Q(D8543_Q), .D(D8514_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8541 ( .Q(D8541_Q), .D(D8511_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8539 ( .Q(D8539_Q), .D(D8506_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8538 ( .Q(D8538_Q), .D(D8507_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8463 ( .Q(D8463_Q), .D(D8402_Y), .CK(D884_Y));
KC_DFFHQ_X1 D8460 ( .Q(D8460_Q), .D(D8426_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8459 ( .Q(D8459_Q), .D(D8425_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8458 ( .Q(D8458_Q), .D(D9686_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D8330 ( .Q(D8330_Q), .D(D8316_Y), .CK(D884_Y));
KC_DFFHQ_X1 D8329 ( .Q(D8329_Q), .D(D8255_Y), .CK(D884_Y));
KC_DFFHQ_X1 D8328 ( .Q(D8328_Q), .D(D8314_Y), .CK(D884_Y));
KC_DFFHQ_X1 D8238 ( .Q(D8238_Q), .D(D8205_Y), .CK(D884_Y));
KC_DFFHQ_X1 D8145 ( .Q(D8145_Q), .D(D8021_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D8055 ( .Q(D8055_Q), .D(D1898_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D8054 ( .Q(D8054_Q), .D(D7998_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D8053 ( .Q(D8053_Q), .D(D8014_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D8052 ( .Q(D8052_Q), .D(D7997_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D8051 ( .Q(D8051_Q), .D(D8022_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D7971 ( .Q(D7971_Q), .D(D6492_Y), .CK(D7964_QN));
KC_DFFHQ_X1 D7970 ( .Q(D7970_Q), .D(D6453_Y), .CK(D7964_QN));
KC_DFFHQ_X1 D7969 ( .Q(D7969_Q), .D(D7868_Y), .CK(D7964_QN));
KC_DFFHQ_X1 D7968 ( .Q(D7968_Q), .D(D7981_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D7967 ( .Q(D7967_Q), .D(D487_Y), .CK(D7964_QN));
KC_DFFHQ_X1 D7966 ( .Q(D7966_Q), .D(D7982_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D7890 ( .Q(D7890_Q), .D(D7847_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7889 ( .Q(D7889_Q), .D(D7853_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7888 ( .Q(D7888_Q), .D(D7876_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7887 ( .Q(D7887_Q), .D(D7871_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7886 ( .Q(D7886_Q), .D(D7873_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7885 ( .Q(D7885_Q), .D(D7870_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7884 ( .Q(D7884_Q), .D(D7897_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7883 ( .Q(D7883_Q), .D(D7900_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D7085 ( .Q(D7085_Q), .D(D8581_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D7084 ( .Q(D7084_Q), .D(D8581_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D7083 ( .Q(D7083_Q), .D(D8581_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D7082 ( .Q(D7082_Q), .D(D8581_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D7081 ( .Q(D7081_Q), .D(D8584_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D7080 ( .Q(D7080_Q), .D(D8584_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D7079 ( .Q(D7079_Q), .D(D8584_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D7078 ( .Q(D7078_Q), .D(D8584_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D7077 ( .Q(D7077_Q), .D(D8629_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D7076 ( .Q(D7076_Q), .D(D8629_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D7075 ( .Q(D7075_Q), .D(D8629_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D7056 ( .Q(D7056_Q), .D(D8570_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D7055 ( .Q(D7055_Q), .D(D8571_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D7054 ( .Q(D7054_Q), .D(D8570_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D7053 ( .Q(D7053_Q), .D(D8571_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D7052 ( .Q(D7052_Q), .D(D8571_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D7051 ( .Q(D7051_Q), .D(D8570_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D7050 ( .Q(D7050_Q), .D(D8570_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D7049 ( .Q(D7049_Q), .D(D8580_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D7048 ( .Q(D7048_Q), .D(D8580_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D7047 ( .Q(D7047_Q), .D(D8570_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D7046 ( .Q(D7046_Q), .D(D8580_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D7045 ( .Q(D7045_Q), .D(D8580_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D7044 ( .Q(D7044_Q), .D(D8627_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D7043 ( .Q(D7043_Q), .D(D8627_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D7042 ( .Q(D7042_Q), .D(D8627_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D7014 ( .Q(D7014_Q), .D(D8570_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D7013 ( .Q(D7013_Q), .D(D8571_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D7012 ( .Q(D7012_Q), .D(D8570_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D7011 ( .Q(D7011_Q), .D(D8571_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D7010 ( .Q(D7010_Q), .D(D8570_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D7009 ( .Q(D7009_Q), .D(D6957_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D7008 ( .Q(D7008_Q), .D(D6995_Y), .CK(D6954_Y));
KC_DFFHQ_X1 D7007 ( .Q(D7007_Q), .D(D6957_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D7006 ( .Q(D7006_Q), .D(D6957_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D7005 ( .Q(D7005_Q), .D(D6993_Y), .CK(D6954_Y));
KC_DFFHQ_X1 D7004 ( .Q(D7004_Q), .D(D8571_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D6970 ( .Q(D6970_Q), .D(D6946_Y), .CK(D6954_Y));
KC_DFFHQ_X1 D6969 ( .Q(D6969_Q), .D(D6890_Y), .CK(D1009_QN));
KC_DFFHQ_X1 D6968 ( .Q(D6968_Q), .D(D1002_Y), .CK(D5462_QN));
KC_DFFHQ_X1 D6967 ( .Q(D6967_Q), .D(D6890_Y), .CK(D893_QN));
KC_DFFHQ_X1 D6966 ( .Q(D6966_Q), .D(D1002_Y), .CK(D1009_QN));
KC_DFFHQ_X1 D6965 ( .Q(D6965_Q), .D(D6939_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D6964 ( .Q(D6964_Q), .D(D1002_Y), .CK(D893_QN));
KC_DFFHQ_X1 D6963 ( .Q(D6963_Q), .D(D6941_Y), .CK(D6954_Y));
KC_DFFHQ_X1 D6962 ( .Q(D6962_Q), .D(D6940_Y), .CK(D6954_Y));
KC_DFFHQ_X1 D6912 ( .Q(D6912_Q), .D(D6891_Y), .CK(D6815_QN));
KC_DFFHQ_X1 D6911 ( .Q(D6911_Q), .D(D6891_Y), .CK(D6814_QN));
KC_DFFHQ_X1 D6903 ( .Q(D6903_Q), .D(D6891_Y), .CK(D6811_QN));
KC_DFFHQ_X1 D6902 ( .Q(D6902_Q), .D(D6890_Y), .CK(D6814_QN));
KC_DFFHQ_X1 D6901 ( .Q(D6901_Q), .D(D6890_Y), .CK(D6815_QN));
KC_DFFHQ_X1 D6900 ( .Q(D6900_Q), .D(D1002_Y), .CK(D6811_QN));
KC_DFFHQ_X1 D6899 ( .Q(D6899_Q), .D(D6797_Y), .CK(D6814_QN));
KC_DFFHQ_X1 D6898 ( .Q(D6898_Q), .D(D1002_Y), .CK(D6815_QN));
KC_DFFHQ_X1 D6897 ( .Q(D6897_Q), .D(D1002_Y), .CK(D6814_QN));
KC_DFFHQ_X1 D6896 ( .Q(D6896_Q), .D(D6891_Y), .CK(D6810_QN));
KC_DFFHQ_X1 D6895 ( .Q(D6895_Q), .D(D6797_Y), .CK(D6815_QN));
KC_DFFHQ_X1 D6894 ( .Q(D6894_Q), .D(D1002_Y), .CK(D6810_QN));
KC_DFFHQ_X1 D6893 ( .Q(D6893_Q), .D(D6891_Y), .CK(D1009_QN));
KC_DFFHQ_X1 D6892 ( .Q(D6892_Q), .D(D6797_Y), .CK(D6810_QN));
KC_DFFHQ_X1 D6830 ( .Q(D6830_Q), .D(D1759_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D6829 ( .Q(D6829_Q), .D(D960_Y), .CK(D884_Y));
KC_DFFHQ_X1 D6828 ( .Q(D6828_Q), .D(D1759_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D6827 ( .Q(D6827_Q), .D(D1759_Y), .CK(D657_QN));
KC_DFFHQ_X1 D6826 ( .Q(D6826_Q), .D(D869_Y), .CK(D884_Y));
KC_DFFHQ_X1 D6825 ( .Q(D6825_Q), .D(D6771_Y), .CK(D884_Y));
KC_DFFHQ_X1 D6824 ( .Q(D6824_Q), .D(D6797_Y), .CK(D6817_QN));
KC_DFFHQ_X1 D6823 ( .Q(D6823_Q), .D(D6797_Y), .CK(D6816_QN));
KC_DFFHQ_X1 D6822 ( .Q(D6822_Q), .D(D6891_Y), .CK(D6816_QN));
KC_DFFHQ_X1 D6821 ( .Q(D6821_Q), .D(D6890_Y), .CK(D6816_QN));
KC_DFFHQ_X1 D6820 ( .Q(D6820_Q), .D(D6890_Y), .CK(D6817_QN));
KC_DFFHQ_X1 D6819 ( .Q(D6819_Q), .D(D6797_Y), .CK(D6811_QN));
KC_DFFHQ_X1 D6818 ( .Q(D6818_Q), .D(D6891_Y), .CK(D6817_QN));
KC_DFFHQ_X1 D6758 ( .Q(D6758_Q), .D(D6718_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D6757 ( .Q(D6757_Q), .D(D6742_Y), .CK(D655_QN));
KC_DFFHQ_X1 D6756 ( .Q(D6756_Q), .D(D6742_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D6755 ( .Q(D6755_Q), .D(D6731_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D6754 ( .Q(D6754_Q), .D(D8203_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D6753 ( .Q(D6753_Q), .D(D6731_Y), .CK(D657_QN));
KC_DFFHQ_X1 D6752 ( .Q(D6752_Q), .D(D6731_Y), .CK(D655_QN));
KC_DFFHQ_X1 D6751 ( .Q(D6751_Q), .D(D6731_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6750 ( .Q(D6750_Q), .D(D8179_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D6749 ( .Q(D6749_Q), .D(D6731_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D6748 ( .Q(D6748_Q), .D(D6805_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D6747 ( .Q(D6747_Q), .D(D6805_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6746 ( .Q(D6746_Q), .D(D1759_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D6745 ( .Q(D6745_Q), .D(D1759_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6744 ( .Q(D6744_Q), .D(D6713_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D6743 ( .Q(D6743_Q), .D(D6805_Y), .CK(D655_QN));
KC_DFFHQ_X1 D6675 ( .Q(D6675_Q), .D(D1760_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D6674 ( .Q(D6674_Q), .D(D1760_Y), .CK(D657_QN));
KC_DFFHQ_X1 D6673 ( .Q(D6673_Q), .D(D6649_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D6672 ( .Q(D6672_Q), .D(D6649_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6671 ( .Q(D6671_Q), .D(D6649_Y), .CK(D655_QN));
KC_DFFHQ_X1 D6670 ( .Q(D6670_Q), .D(D6649_Y), .CK(D657_QN));
KC_DFFHQ_X1 D6669 ( .Q(D6669_Q), .D(D1760_Y), .CK(D655_QN));
KC_DFFHQ_X1 D6668 ( .Q(D6668_Q), .D(D1760_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D6667 ( .Q(D6667_Q), .D(D1760_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6666 ( .Q(D6666_Q), .D(D576_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6663 ( .Q(D6663_Q), .D(D6645_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D6662 ( .Q(D6662_Q), .D(D6645_Y), .CK(D655_QN));
KC_DFFHQ_X1 D6661 ( .Q(D6661_Q), .D(D6645_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D6660 ( .Q(D6660_Q), .D(D6645_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D6659 ( .Q(D6659_Q), .D(D6645_Y), .CK(D657_QN));
KC_DFFHQ_X1 D6658 ( .Q(D6658_Q), .D(D6645_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6657 ( .Q(D6657_Q), .D(D6742_Y), .CK(D657_QN));
KC_DFFHQ_X1 D6656 ( .Q(D6656_Q), .D(D6742_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D6655 ( .Q(D6655_Q), .D(D6742_Y), .CK(D5217_QN));
KC_DFFHQ_X1 D6652 ( .Q(D6652_Q), .D(D6649_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D6612 ( .Q(D6612_Q), .D(D8038_Y), .CK(D586_QN));
KC_DFFHQ_X1 D6611 ( .Q(D6611_Q), .D(D8038_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D6610 ( .Q(D6610_Q), .D(D8038_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D6609 ( .Q(D6609_Q), .D(D8038_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D6608 ( .Q(D6608_Q), .D(D8038_Y), .CK(D587_QN));
KC_DFFHQ_X1 D6607 ( .Q(D6607_Q), .D(D577_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D6606 ( .Q(D6606_Q), .D(D577_Y), .CK(D586_QN));
KC_DFFHQ_X1 D6605 ( .Q(D6605_Q), .D(D100_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D6604 ( .Q(D6604_Q), .D(D100_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D6603 ( .Q(D6603_Q), .D(D100_Y), .CK(D586_QN));
KC_DFFHQ_X1 D6602 ( .Q(D6602_Q), .D(D577_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D6601 ( .Q(D6601_Q), .D(D100_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D6600 ( .Q(D6600_Q), .D(D577_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D6599 ( .Q(D6599_Q), .D(D577_Y), .CK(D587_QN));
KC_DFFHQ_X1 D6598 ( .Q(D6598_Q), .D(D577_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D6597 ( .Q(D6597_Q), .D(D8038_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D6596 ( .Q(D6596_Q), .D(D6614_Y), .CK(D586_QN));
KC_DFFHQ_X1 D6595 ( .Q(D6595_Q), .D(D100_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D6594 ( .Q(D6594_Q), .D(D100_Y), .CK(D587_QN));
KC_DFFHQ_X1 D6555 ( .Q(D6555_Q), .D(D6510_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D6554 ( .Q(D6554_Q), .D(D6515_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D6553 ( .Q(D6553_Q), .D(D6537_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D6552 ( .Q(D6552_Q), .D(D10144_Y), .CK(D6538_QN));
KC_DFFHQ_X1 D6551 ( .Q(D6551_Q), .D(D6529_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D6550 ( .Q(D6550_Q), .D(D6530_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D6549 ( .Q(D6549_Q), .D(D6535_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D6548 ( .Q(D6548_Q), .D(D6536_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D6547 ( .Q(D6547_Q), .D(D6533_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D6546 ( .Q(D6546_Q), .D(D6531_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D6544 ( .Q(D6544_Q), .D(D6527_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D6540 ( .Q(D6540_Q), .D(D7956_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D6539 ( .Q(D6539_Q), .D(D6523_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D6476 ( .Q(D6476_Q), .D(D1666_Y), .CK(D6466_QN));
KC_DFFHQ_X1 D6475 ( .Q(D6475_Q), .D(D6459_Y), .CK(D6466_QN));
KC_DFFHQ_X1 D6474 ( .Q(D6474_Q), .D(D5086_Y), .CK(D6466_QN));
KC_DFFHQ_X1 D6473 ( .Q(D6473_Q), .D(D1809_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D6472 ( .Q(D6472_Q), .D(D5063_Y), .CK(D6466_QN));
KC_DFFHQ_X1 D6376 ( .Q(D6376_Q), .D(D439_Y), .CK(D6374_QN));
KC_DFFHQ_X1 D6375 ( .Q(D6375_Q), .D(D6404_Y), .CK(D6374_QN));
KC_DFFHQ_X1 D5633 ( .Q(D5633_Q), .D(D7003_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D5632 ( .Q(D5632_Q), .D(D7018_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D5631 ( .Q(D5631_Q), .D(D7018_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D5630 ( .Q(D5630_Q), .D(D7018_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D5629 ( .Q(D5629_Q), .D(D7003_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D5628 ( .Q(D5628_Q), .D(D7003_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D5627 ( .Q(D5627_Q), .D(D7018_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D5626 ( .Q(D5626_Q), .D(D7003_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D5625 ( .Q(D5625_Q), .D(D7003_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D5624 ( .Q(D5624_Q), .D(D7003_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D5610 ( .Q(D5610_Q), .D(D7002_Y), .CK(D4042_QN));
KC_DFFHQ_X1 D5609 ( .Q(D5609_Q), .D(D7002_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D5608 ( .Q(D5608_Q), .D(D7002_Y), .CK(D4040_QN));
KC_DFFHQ_X1 D5607 ( .Q(D5607_Q), .D(D7018_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D5606 ( .Q(D5606_Q), .D(D7018_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D5605 ( .Q(D5605_Q), .D(D7003_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D5604 ( .Q(D5604_Q), .D(D7003_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D5603 ( .Q(D5603_Q), .D(D5640_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D5574 ( .Q(D5574_Q), .D(D6909_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D5573 ( .Q(D5573_Q), .D(D6957_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D5571 ( .Q(D5571_Q), .D(D6956_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D5570 ( .Q(D5570_Q), .D(D6952_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D5569 ( .Q(D5569_Q), .D(D7002_Y), .CK(D4008_QN));
KC_DFFHQ_X1 D5568 ( .Q(D5568_Q), .D(D7002_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D5567 ( .Q(D5567_Q), .D(D7002_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D5566 ( .Q(D5566_Q), .D(D7002_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D5565 ( .Q(D5565_Q), .D(D6956_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D5564 ( .Q(D5564_Q), .D(D6909_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D5563 ( .Q(D5563_Q), .D(D6956_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D5562 ( .Q(D5562_Q), .D(D6909_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D5561 ( .Q(D5561_Q), .D(D6956_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D5560 ( .Q(D5560_Q), .D(D6956_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D5534 ( .Q(D5534_Q), .D(D6957_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D5533 ( .Q(D5533_Q), .D(D6957_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D5532 ( .Q(D5532_Q), .D(D6952_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D5531 ( .Q(D5531_Q), .D(D6956_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D5530 ( .Q(D5530_Q), .D(D5458_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D5529 ( .Q(D5529_Q), .D(D5455_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D5528 ( .Q(D5528_Q), .D(D6909_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D5527 ( .Q(D5527_Q), .D(D5458_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D5526 ( .Q(D5526_Q), .D(D5456_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D5525 ( .Q(D5525_Q), .D(D6952_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D5524 ( .Q(D5524_Q), .D(D6909_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D5492 ( .Q(D5492_Q), .D(D1619_Y), .CK(D891_QN));
KC_DFFHQ_X1 D5491 ( .Q(D5491_Q), .D(D1619_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D5476 ( .Q(D5476_Q), .D(D1619_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D5474 ( .Q(D5474_Q), .D(D1619_Y), .CK(D892_QN));
KC_DFFHQ_X1 D5472 ( .Q(D5472_Q), .D(D5457_Y), .CK(D892_QN));
KC_DFFHQ_X1 D5471 ( .Q(D5471_Q), .D(D6273_Y), .CK(D892_QN));
KC_DFFHQ_X1 D5470 ( .Q(D5470_Q), .D(D5455_Y), .CK(D891_QN));
KC_DFFHQ_X1 D5469 ( .Q(D5469_Q), .D(D5458_Y), .CK(D892_QN));
KC_DFFHQ_X1 D5468 ( .Q(D5468_Q), .D(D5455_Y), .CK(D892_QN));
KC_DFFHQ_X1 D5467 ( .Q(D5467_Q), .D(D5458_Y), .CK(D891_QN));
KC_DFFHQ_X1 D5466 ( .Q(D5466_Q), .D(D5456_Y), .CK(D891_QN));
KC_DFFHQ_X1 D5465 ( .Q(D5465_Q), .D(D6797_Y), .CK(D5462_QN));
KC_DFFHQ_X1 D5464 ( .Q(D5464_Q), .D(D5456_Y), .CK(D892_QN));
KC_DFFHQ_X1 D5463 ( .Q(D5463_Q), .D(D5456_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D5402 ( .Q(D5402_Q), .D(D5386_Y), .CK(D894_QN));
KC_DFFHQ_X1 D5401 ( .Q(D5401_Q), .D(D5386_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D5400 ( .Q(D5400_Q), .D(D5386_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D5399 ( .Q(D5399_Q), .D(D5379_Y), .CK(D891_QN));
KC_DFFHQ_X1 D5398 ( .Q(D5398_Q), .D(D5379_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D5397 ( .Q(D5397_Q), .D(D5379_Y), .CK(D892_QN));
KC_DFFHQ_X1 D5396 ( .Q(D5396_Q), .D(D5379_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D5395 ( .Q(D5395_Q), .D(D5379_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D5394 ( .Q(D5394_Q), .D(D5379_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D5321 ( .Q(D5321_Q), .D(D6742_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5320 ( .Q(D5320_Q), .D(D5297_Y), .CK(D894_QN));
KC_DFFHQ_X1 D5319 ( .Q(D5319_Q), .D(D5297_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D5318 ( .Q(D5318_Q), .D(D6731_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5317 ( .Q(D5317_Q), .D(D5296_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D5316 ( .Q(D5316_Q), .D(D5296_Y), .CK(D894_QN));
KC_DFFHQ_X1 D5315 ( .Q(D5315_Q), .D(D6731_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5314 ( .Q(D5314_Q), .D(D5297_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D5313 ( .Q(D5313_Q), .D(D6805_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5312 ( .Q(D5312_Q), .D(D6805_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5311 ( .Q(D5311_Q), .D(D5298_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D5310 ( .Q(D5310_Q), .D(D5297_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D5309 ( .Q(D5309_Q), .D(D5296_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D5308 ( .Q(D5308_Q), .D(D1759_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5307 ( .Q(D5307_Q), .D(D1759_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5306 ( .Q(D5306_Q), .D(D5296_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D5305 ( .Q(D5305_Q), .D(D5382_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D5304 ( .Q(D5304_Q), .D(D5382_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D5303 ( .Q(D5303_Q), .D(D5382_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D5302 ( .Q(D5302_Q), .D(D5382_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D5240 ( .Q(D5240_Q), .D(D576_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D5239 ( .Q(D5239_Q), .D(D576_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D5238 ( .Q(D5238_Q), .D(D576_Y), .CK(D657_QN));
KC_DFFHQ_X1 D5237 ( .Q(D5237_Q), .D(D576_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5236 ( .Q(D5236_Q), .D(D576_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5235 ( .Q(D5235_Q), .D(D1760_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D5234 ( .Q(D5234_Q), .D(D1760_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5233 ( .Q(D5233_Q), .D(D576_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D5232 ( .Q(D5232_Q), .D(D6649_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5231 ( .Q(D5231_Q), .D(D1760_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5230 ( .Q(D5230_Q), .D(D5298_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D5229 ( .Q(D5229_Q), .D(D5297_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D5228 ( .Q(D5228_Q), .D(D6649_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5227 ( .Q(D5227_Q), .D(D6645_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5226 ( .Q(D5226_Q), .D(D5298_Y), .CK(D894_QN));
KC_DFFHQ_X1 D5225 ( .Q(D5225_Q), .D(D5296_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D5224 ( .Q(D5224_Q), .D(D6742_Y), .CK(D656_QN));
KC_DFFHQ_X1 D5223 ( .Q(D5223_Q), .D(D6645_Y), .CK(D5218_QN));
KC_DFFHQ_X1 D5222 ( .Q(D5222_Q), .D(D5297_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D5221 ( .Q(D5221_Q), .D(D5296_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D5198 ( .Q(D5198_Q), .D(D8059_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D5197 ( .Q(D5197_Q), .D(D580_Y), .CK(D586_QN));
KC_DFFHQ_X1 D5196 ( .Q(D5196_Q), .D(D8059_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D5195 ( .Q(D5195_Q), .D(D8059_Y), .CK(D586_QN));
KC_DFFHQ_X1 D5194 ( .Q(D5194_Q), .D(D6613_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D5193 ( .Q(D5193_Q), .D(D579_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D5192 ( .Q(D5192_Q), .D(D579_Y), .CK(D587_QN));
KC_DFFHQ_X1 D5191 ( .Q(D5191_Q), .D(D6613_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D5190 ( .Q(D5190_Q), .D(D579_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D5189 ( .Q(D5189_Q), .D(D6613_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D5188 ( .Q(D5188_Q), .D(D579_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D5187 ( .Q(D5187_Q), .D(D579_Y), .CK(D586_QN));
KC_DFFHQ_X1 D5186 ( .Q(D5186_Q), .D(D6614_Y), .CK(D587_QN));
KC_DFFHQ_X1 D5185 ( .Q(D5185_Q), .D(D8059_Y), .CK(D587_QN));
KC_DFFHQ_X1 D5142 ( .Q(D5142_Q), .D(D4990_Y), .CK(D478_QN));
KC_DFFHQ_X1 D5141 ( .Q(D5141_Q), .D(D5049_Y), .CK(D478_QN));
KC_DFFHQ_X1 D5140 ( .Q(D5140_Q), .D(D1621_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D5139 ( .Q(D5139_Q), .D(D5120_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D5138 ( .Q(D5138_Q), .D(D5087_Y), .CK(D6538_QN));
KC_DFFHQ_X1 D5137 ( .Q(D5137_Q), .D(D5121_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D5136 ( .Q(D5136_Q), .D(D5117_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D5135 ( .Q(D5135_Q), .D(D5118_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D5134 ( .Q(D5134_Q), .D(D5115_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D5133 ( .Q(D5133_Q), .D(D5107_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D5132 ( .Q(D5132_Q), .D(D5111_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D5131 ( .Q(D5131_Q), .D(D6528_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D5130 ( .Q(D5130_Q), .D(D5113_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D5129 ( .Q(D5129_Q), .D(D5112_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D5128 ( .Q(D5128_Q), .D(D5105_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D5127 ( .Q(D5127_Q), .D(D580_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D5126 ( .Q(D5126_Q), .D(D580_Y), .CK(D587_QN));
KC_DFFHQ_X1 D5125 ( .Q(D5125_Q), .D(D5099_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D5124 ( .Q(D5124_Q), .D(D5106_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D5123 ( .Q(D5123_Q), .D(D5108_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D5078 ( .Q(D5078_Q), .D(D5075_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D4083 ( .Q(D4083_Q), .D(D5640_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D4082 ( .Q(D4082_Q), .D(D5640_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D4081 ( .Q(D4081_Q), .D(D7018_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D4080 ( .Q(D4080_Q), .D(D7018_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D4051 ( .Q(D4051_Q), .D(D5555_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D4050 ( .Q(D4050_Q), .D(D5555_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D4049 ( .Q(D4049_Q), .D(D5555_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D4048 ( .Q(D4048_Q), .D(D5555_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D4047 ( .Q(D4047_Q), .D(D5555_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D4045 ( .Q(D4045_Q), .D(D5640_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D3985 ( .Q(D3985_Q), .D(D5455_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3975 ( .Q(D3975_Q), .D(D5456_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3974 ( .Q(D3974_Q), .D(D5458_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3973 ( .Q(D3973_Q), .D(D6909_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D3972 ( .Q(D3972_Q), .D(D6952_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D3969 ( .Q(D3969_Q), .D(D5458_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D3968 ( .Q(D3968_Q), .D(D5458_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3967 ( .Q(D3967_Q), .D(D5457_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3966 ( .Q(D3966_Q), .D(D5455_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3965 ( .Q(D3965_Q), .D(D5456_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D3964 ( .Q(D3964_Q), .D(D5455_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3963 ( .Q(D3963_Q), .D(D5458_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3962 ( .Q(D3962_Q), .D(D5456_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3961 ( .Q(D3961_Q), .D(D6952_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D3960 ( .Q(D3960_Q), .D(D5457_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3959 ( .Q(D3959_Q), .D(D5456_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3944 ( .Q(D3944_Q), .D(D1618_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3943 ( .Q(D3943_Q), .D(D1618_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3942 ( .Q(D3942_Q), .D(D1618_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D3941 ( .Q(D3941_Q), .D(D1618_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D3940 ( .Q(D3940_Q), .D(D1618_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3939 ( .Q(D3939_Q), .D(D1619_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3938 ( .Q(D3938_Q), .D(D1619_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3937 ( .Q(D3937_Q), .D(D5457_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D3936 ( .Q(D3936_Q), .D(D5457_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D3935 ( .Q(D3935_Q), .D(D1619_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3934 ( .Q(D3934_Q), .D(D5457_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D3933 ( .Q(D3933_Q), .D(D5457_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D3932 ( .Q(D3932_Q), .D(D6273_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3931 ( .Q(D3931_Q), .D(D6273_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3930 ( .Q(D3930_Q), .D(D6273_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D3929 ( .Q(D3929_Q), .D(D6273_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D3928 ( .Q(D3928_Q), .D(D5457_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3927 ( .Q(D3927_Q), .D(D6273_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3926 ( .Q(D3926_Q), .D(D6273_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D3925 ( .Q(D3925_Q), .D(D6273_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D3880 ( .Q(D3880_Q), .D(D5386_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3879 ( .Q(D3879_Q), .D(D5386_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D3878 ( .Q(D3878_Q), .D(D5386_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D3877 ( .Q(D3877_Q), .D(D5379_Y), .CK(D3866_QN));
KC_DFFHQ_X1 D3876 ( .Q(D3876_Q), .D(D5379_Y), .CK(D3865_QN));
KC_DFFHQ_X1 D3875 ( .Q(D3875_Q), .D(D5379_Y), .CK(D1484_QN));
KC_DFFHQ_X1 D3874 ( .Q(D3874_Q), .D(D1618_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D3819 ( .Q(D3819_Q), .D(D5299_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3818 ( .Q(D3818_Q), .D(D5300_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D3817 ( .Q(D3817_Q), .D(D5299_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D3816 ( .Q(D3816_Q), .D(D5299_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D3815 ( .Q(D3815_Q), .D(D5300_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3814 ( .Q(D3814_Q), .D(D5299_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D3813 ( .Q(D3813_Q), .D(D5299_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D3812 ( .Q(D3812_Q), .D(D5300_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D3811 ( .Q(D3811_Q), .D(D5299_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D3810 ( .Q(D3810_Q), .D(D5300_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D3809 ( .Q(D3809_Q), .D(D5300_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D3808 ( .Q(D3808_Q), .D(D5299_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D3807 ( .Q(D3807_Q), .D(D5381_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3806 ( .Q(D3806_Q), .D(D5299_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D3805 ( .Q(D3805_Q), .D(D5381_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D3804 ( .Q(D3804_Q), .D(D5381_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D3803 ( .Q(D3803_Q), .D(D5381_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D3802 ( .Q(D3802_Q), .D(D5382_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3801 ( .Q(D3801_Q), .D(D5381_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D3800 ( .Q(D3800_Q), .D(D5381_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D3799 ( .Q(D3799_Q), .D(D5381_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D3743 ( .Q(D3743_Q), .D(D5298_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D3742 ( .Q(D3742_Q), .D(D5298_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3741 ( .Q(D3741_Q), .D(D5297_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D3740 ( .Q(D3740_Q), .D(D5297_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3739 ( .Q(D3739_Q), .D(D5296_Y), .CK(D3870_QN));
KC_DFFHQ_X1 D3738 ( .Q(D3738_Q), .D(D5296_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D3737 ( .Q(D3737_Q), .D(D100_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D3736 ( .Q(D3736_Q), .D(D100_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D3735 ( .Q(D3735_Q), .D(D100_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D3734 ( .Q(D3734_Q), .D(D5296_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D3733 ( .Q(D3733_Q), .D(D5298_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D3728 ( .Q(D3728_Q), .D(D5297_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D3727 ( .Q(D3727_Q), .D(D5298_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D3726 ( .Q(D3726_Q), .D(D5300_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D3725 ( .Q(D3725_Q), .D(D5299_Y), .CK(D894_QN));
KC_DFFHQ_X1 D3686 ( .Q(D3686_Q), .D(D8059_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D3685 ( .Q(D3685_Q), .D(D8059_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D3684 ( .Q(D3684_Q), .D(D8059_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D3683 ( .Q(D3683_Q), .D(D6614_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D3682 ( .Q(D3682_Q), .D(D577_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D3681 ( .Q(D3681_Q), .D(D577_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D3680 ( .Q(D3680_Q), .D(D579_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D3679 ( .Q(D3679_Q), .D(D579_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D3678 ( .Q(D3678_Q), .D(D6613_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D3677 ( .Q(D3677_Q), .D(D6613_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D3676 ( .Q(D3676_Q), .D(D577_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D3675 ( .Q(D3675_Q), .D(D579_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D3674 ( .Q(D3674_Q), .D(D6614_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D3673 ( .Q(D3673_Q), .D(D6614_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D3672 ( .Q(D3672_Q), .D(D6613_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D3632 ( .Q(D3632_Q), .D(D3622_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D3631 ( .Q(D3631_Q), .D(D3618_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D3630 ( .Q(D3630_Q), .D(D3610_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D3629 ( .Q(D3629_Q), .D(D3611_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D3628 ( .Q(D3628_Q), .D(D3604_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D3627 ( .Q(D3627_Q), .D(D580_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D3626 ( .Q(D3626_Q), .D(D8038_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D3625 ( .Q(D3625_Q), .D(D8038_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D3624 ( .Q(D3624_Q), .D(D3607_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D3576 ( .Q(D3576_Q), .D(D1463_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D3575 ( .Q(D3575_Q), .D(D3558_Y), .CK(D4957_QN));
KC_DFFHQ_X1 D3376 ( .Q(D3376_Q), .D(D3354_Y), .CK(D4958_QN));
KC_DFFHQ_X1 D3375 ( .Q(D3375_Q), .D(D408_Y), .CK(D4958_QN));
KC_DFFHQ_X1 D3374 ( .Q(D3374_Q), .D(D3395_Y), .CK(D4958_QN));
KC_DFFHQ_X1 D3373 ( .Q(D3373_Q), .D(D1416_Y), .CK(D4958_QN));
KC_DFFHQ_X1 D3372 ( .Q(D3372_Q), .D(D4782_Y), .CK(D4958_QN));
KC_DFFHQ_X1 D2467 ( .Q(D2467_Q), .D(D2303_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D2389 ( .Q(D2389_Q), .D(D11851_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D2388 ( .Q(D2388_Q), .D(D11453_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D2387 ( .Q(D2387_Q), .D(D1161_Y), .CK(D11916_QN));
KC_DFFHQ_X1 D2385 ( .Q(D2385_Q), .D(D2303_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D2384 ( .Q(D2384_Q), .D(D2302_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D2352 ( .Q(D2352_Q), .D(D11851_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D2351 ( .Q(D2351_Q), .D(D11851_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D2350 ( .Q(D2350_Q), .D(D11849_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D2349 ( .Q(D2349_Q), .D(D11453_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D2348 ( .Q(D2348_Q), .D(D11994_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D2347 ( .Q(D2347_Q), .D(D11966_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D2346 ( .Q(D2346_Q), .D(D12053_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D2345 ( .Q(D2345_Q), .D(D12056_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D2344 ( .Q(D2344_Q), .D(D11992_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D2297 ( .Q(D2297_Q), .D(D11778_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D2296 ( .Q(D2296_Q), .D(D11779_Y), .CK(D718_QN));
KC_DFFHQ_X1 D2295 ( .Q(D2295_Q), .D(D11778_Y), .CK(D11171_QN));
KC_DFFHQ_X1 D2294 ( .Q(D2294_Q), .D(D11908_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D2293 ( .Q(D2293_Q), .D(D11849_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D2292 ( .Q(D2292_Q), .D(D11992_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D2291 ( .Q(D2291_Q), .D(D11968_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D2290 ( .Q(D2290_Q), .D(D11477_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D2289 ( .Q(D2289_Q), .D(D11968_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D2288 ( .Q(D2288_Q), .D(D11786_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D2256 ( .Q(D2256_Q), .D(D11196_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D2255 ( .Q(D2255_Q), .D(D1007_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D2254 ( .Q(D2254_Q), .D(D10415_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D2253 ( .Q(D2253_Q), .D(D11352_Y), .CK(D10412_Y));
KC_DFFHQ_X1 D2252 ( .Q(D2252_Q), .D(D10503_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D2251 ( .Q(D2251_Q), .D(D11509_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D2250 ( .Q(D2250_Q), .D(D78_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D2249 ( .Q(D2249_Q), .D(D11502_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D2248 ( .Q(D2248_Q), .D(D11477_Y), .CK(D12041_QN));
KC_DFFHQ_X1 D2247 ( .Q(D2247_Q), .D(D11253_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D2246 ( .Q(D2246_Q), .D(D11253_Y), .CK(D588_QN));
KC_DFFHQ_X1 D2245 ( .Q(D2245_Q), .D(D11253_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D2221 ( .Q(D2221_Q), .D(D8320_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D2220 ( .Q(D2220_Q), .D(D9777_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D2219 ( .Q(D2219_Q), .D(D10507_Y), .CK(D901_QN));
KC_DFFHQ_X1 D2218 ( .Q(D2218_Q), .D(D10492_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D2217 ( .Q(D2217_Q), .D(D10498_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D2216 ( .Q(D2216_Q), .D(D9780_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D2215 ( .Q(D2215_Q), .D(D9780_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D2214 ( .Q(D2214_Q), .D(D834_Y), .CK(D588_QN));
KC_DFFHQ_X1 D2213 ( .Q(D2213_Q), .D(D10823_Y), .CK(D11134_QN));
KC_DFFHQ_X1 D2161 ( .Q(D2161_Q), .D(D9795_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D2159 ( .Q(D2159_Q), .D(D10542_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D2157 ( .Q(D2157_Q), .D(D10477_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D2156 ( .Q(D2156_Q), .D(D10498_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D2085 ( .Q(D2085_Q), .D(D8573_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D2084 ( .Q(D2084_Q), .D(D8573_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D2083 ( .Q(D2083_Q), .D(D9833_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D2082 ( .Q(D2082_Q), .D(D9833_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D2081 ( .Q(D2081_Q), .D(D9695_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D2080 ( .Q(D2080_Q), .D(D9702_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D2079 ( .Q(D2079_Q), .D(D90_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D2078 ( .Q(D2078_Q), .D(D8573_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D1933 ( .Q(D1933_Q), .D(D8580_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D1931 ( .Q(D1931_Q), .D(D8169_Y), .CK(D884_Y));
KC_DFFHQ_X1 D1930 ( .Q(D1930_Q), .D(D8411_Y), .CK(D884_Y));
KC_DFFHQ_X1 D1929 ( .Q(D1929_Q), .D(D1078_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D1928 ( .Q(D1928_Q), .D(D1890_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D1927 ( .Q(D1927_Q), .D(D8505_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D1786 ( .Q(D1786_Q), .D(D6516_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D1785 ( .Q(D1785_Q), .D(D4995_Y), .CK(D478_QN));
KC_DFFHQ_X1 D1784 ( .Q(D1784_Q), .D(D8571_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D1783 ( .Q(D1783_Q), .D(D8571_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D1782 ( .Q(D1782_Q), .D(D1759_Y), .CK(D655_QN));
KC_DFFHQ_X1 D1781 ( .Q(D1781_Q), .D(D6805_Y), .CK(D657_QN));
KC_DFFHQ_X1 D1780 ( .Q(D1780_Q), .D(D6805_Y), .CK(D5216_QN));
KC_DFFHQ_X1 D1779 ( .Q(D1779_Q), .D(D983_Y), .CK(D884_Y));
KC_DFFHQ_X1 D1778 ( .Q(D1778_Q), .D(D6890_Y), .CK(D6811_QN));
KC_DFFHQ_X1 D1777 ( .Q(D1777_Q), .D(D6890_Y), .CK(D6810_QN));
KC_DFFHQ_X1 D1776 ( .Q(D1776_Q), .D(D6797_Y), .CK(D1009_QN));
KC_DFFHQ_X1 D1775 ( .Q(D1775_Q), .D(D6891_Y), .CK(D5462_QN));
KC_DFFHQ_X1 D1774 ( .Q(D1774_Q), .D(D1742_Y), .CK(D6954_Y));
KC_DFFHQ_X1 D1773 ( .Q(D1773_Q), .D(D6957_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D1645 ( .Q(D1645_Q), .D(D1601_Y), .CK(D478_QN));
KC_DFFHQ_X1 D1644 ( .Q(D1644_Q), .D(D5119_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D1643 ( .Q(D1643_Q), .D(D6614_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D1642 ( .Q(D1642_Q), .D(D580_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D1641 ( .Q(D1641_Q), .D(D5101_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D1640 ( .Q(D1640_Q), .D(D580_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D1639 ( .Q(D1639_Q), .D(D7002_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D1638 ( .Q(D1638_Q), .D(D5386_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D1637 ( .Q(D1637_Q), .D(D5386_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D1636 ( .Q(D1636_Q), .D(D5382_Y), .CK(D894_QN));
KC_DFFHQ_X1 D1635 ( .Q(D1635_Q), .D(D1619_Y), .CK(D3864_QN));
KC_DFFHQ_X1 D1634 ( .Q(D1634_Q), .D(D5455_Y), .CK(D3868_QN));
KC_DFFHQ_X1 D1633 ( .Q(D1633_Q), .D(D6909_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D1503 ( .Q(D1503_Q), .D(D580_Y), .CK(D3671_QN));
KC_DFFHQ_X1 D1502 ( .Q(D1502_Q), .D(D8038_Y), .CK(D3722_QN));
KC_DFFHQ_X1 D1501 ( .Q(D1501_Q), .D(D580_Y), .CK(D3724_QN));
KC_DFFHQ_X1 D1500 ( .Q(D1500_Q), .D(D5555_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D1499 ( .Q(D1499_Q), .D(D5555_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D1498 ( .Q(D1498_Q), .D(D5382_Y), .CK(D3797_QN));
KC_DFFHQ_X1 D1497 ( .Q(D1497_Q), .D(D5382_Y), .CK(D3798_QN));
KC_DFFHQ_X1 D1496 ( .Q(D1496_Q), .D(D1618_Y), .CK(D892_QN));
KC_DFFHQ_X1 D1495 ( .Q(D1495_Q), .D(D1618_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D1494 ( .Q(D1494_Q), .D(D5455_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D1493 ( .Q(D1493_Q), .D(D5455_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D1403 ( .Q(D1403_Q), .D(D5640_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D1369 ( .Q(D1369_Q), .D(D11586_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D1368 ( .Q(D1368_Q), .D(D1955_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D1367 ( .Q(D1367_Q), .D(D11994_Y), .CK(D12114_QN));
KC_DFFHQ_X1 D1366 ( .Q(D1366_Q), .D(D1955_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D1365 ( .Q(D1365_Q), .D(D11994_Y), .CK(D12113_QN));
KC_DFFHQ_X1 D1364 ( .Q(D1364_Q), .D(D10562_Y), .CK(D11103_QN));
KC_DFFHQ_X1 D1363 ( .Q(D1363_Q), .D(D8626_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D1362 ( .Q(D1362_Q), .D(D12057_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D1361 ( .Q(D1361_Q), .D(D2302_Y), .CK(D12115_QN));
KC_DFFHQ_X1 D1360 ( .Q(D1360_Q), .D(D12057_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D1359 ( .Q(D1359_Q), .D(D2302_Y), .CK(D1347_QN));
KC_DFFHQ_X1 D1358 ( .Q(D1358_Q), .D(D12055_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D1357 ( .Q(D1357_Q), .D(D8585_Y), .CK(D11066_QN));
KC_DFFHQ_X1 D1356 ( .Q(D1356_Q), .D(D8581_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D1355 ( .Q(D1355_Q), .D(D7018_Y), .CK(D4007_QN));
KC_DFFHQ_X1 D1354 ( .Q(D1354_Q), .D(D8585_Y), .CK(D2153_QN));
KC_DFFHQ_X1 D1353 ( .Q(D1353_Q), .D(D8584_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D1352 ( .Q(D1352_Q), .D(D8584_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D1351 ( .Q(D1351_Q), .D(D8585_Y), .CK(D11067_QN));
KC_DFFHQ_X1 D1350 ( .Q(D1350_Q), .D(D8627_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D1349 ( .Q(D1349_Q), .D(D8629_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D1348 ( .Q(D1348_Q), .D(D7003_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D1317 ( .Q(D1317_Q), .D(D11534_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D1316 ( .Q(D1316_Q), .D(D11534_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D1315 ( .Q(D1315_Q), .D(D10562_Y), .CK(D9783_QN));
KC_DFFHQ_X1 D1314 ( .Q(D1314_Q), .D(D10542_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D1313 ( .Q(D1313_Q), .D(D11994_Y), .CK(D1287_QN));
KC_DFFHQ_X1 D1312 ( .Q(D1312_Q), .D(D11477_Y), .CK(D11579_QN));
KC_DFFHQ_X1 D1311 ( .Q(D1311_Q), .D(D11586_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D1310 ( .Q(D1310_Q), .D(D11586_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D1309 ( .Q(D1309_Q), .D(D10563_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D1308 ( .Q(D1308_Q), .D(D11993_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D1307 ( .Q(D1307_Q), .D(D2302_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D1306 ( .Q(D1306_Q), .D(D2302_Y), .CK(D11577_QN));
KC_DFFHQ_X1 D1305 ( .Q(D1305_Q), .D(D12055_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D1304 ( .Q(D1304_Q), .D(D11993_Y), .CK(D11595_QN));
KC_DFFHQ_X1 D1303 ( .Q(D1303_Q), .D(D10542_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D1302 ( .Q(D1302_Q), .D(D10542_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D1301 ( .Q(D1301_Q), .D(D8572_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D1300 ( .Q(D1300_Q), .D(D8580_Y), .CK(D4028_QN));
KC_DFFHQ_X1 D1299 ( .Q(D1299_Q), .D(D7002_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D1298 ( .Q(D1298_Q), .D(D8580_Y), .CK(D4009_QN));
KC_DFFHQ_X1 D1297 ( .Q(D1297_Q), .D(D8626_Y), .CK(D1198_QN));
KC_DFFHQ_X1 D1296 ( .Q(D1296_Q), .D(D8583_Y), .CK(D10543_QN));
KC_DFFHQ_X1 D1295 ( .Q(D1295_Q), .D(D8581_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D1294 ( .Q(D1294_Q), .D(D5640_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D1293 ( .Q(D1293_Q), .D(D5640_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D1292 ( .Q(D1292_Q), .D(D8580_Y), .CK(D4041_QN));
KC_DFFHQ_X1 D1291 ( .Q(D1291_Q), .D(D5640_Y), .CK(D4011_QN));
KC_DFFHQ_X1 D1290 ( .Q(D1290_Q), .D(D8626_Y), .CK(D10593_QN));
KC_DFFHQ_X1 D1289 ( .Q(D1289_Q), .D(D8585_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D1288 ( .Q(D1288_Q), .D(D5640_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D1247 ( .Q(D1247_Q), .D(D12053_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D1246 ( .Q(D1246_Q), .D(D11510_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D1227 ( .Q(D1227_Q), .D(D11966_Y), .CK(D11578_QN));
KC_DFFHQ_X1 D1226 ( .Q(D1226_Q), .D(D10496_Y), .CK(D11102_QN));
KC_DFFHQ_X1 D1225 ( .Q(D1225_Q), .D(D11994_Y), .CK(D11581_QN));
KC_DFFHQ_X1 D1224 ( .Q(D1224_Q), .D(D11999_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D1223 ( .Q(D1223_Q), .D(D10496_Y), .CK(D111_QN));
KC_DFFHQ_X1 D1222 ( .Q(D1222_Q), .D(D11966_Y), .CK(D11580_QN));
KC_DFFHQ_X1 D1221 ( .Q(D1221_Q), .D(D10498_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D1220 ( .Q(D1220_Q), .D(D10492_Y), .CK(D1197_QN));
KC_DFFHQ_X1 D1219 ( .Q(D1219_Q), .D(D11486_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D1218 ( .Q(D1218_Q), .D(D11506_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D1217 ( .Q(D1217_Q), .D(D12057_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D1216 ( .Q(D1216_Q), .D(D12054_Y), .CK(D11070_QN));
KC_DFFHQ_X1 D1215 ( .Q(D1215_Q), .D(D10492_Y), .CK(D111_QN));
KC_DFFHQ_X1 D1214 ( .Q(D1214_Q), .D(D2303_Y), .CK(D11582_QN));
KC_DFFHQ_X1 D1213 ( .Q(D1213_Q), .D(D12057_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D1212 ( .Q(D1212_Q), .D(D1187_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D1211 ( .Q(D1211_Q), .D(D8571_Y), .CK(D5559_QN));
KC_DFFHQ_X1 D1210 ( .Q(D1210_Q), .D(D6909_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D1209 ( .Q(D1209_Q), .D(D8572_Y), .CK(D2071_QN));
KC_DFFHQ_X1 D1208 ( .Q(D1208_Q), .D(D8572_Y), .CK(D11068_QN));
KC_DFFHQ_X1 D1207 ( .Q(D1207_Q), .D(D8570_Y), .CK(D4016_QN));
KC_DFFHQ_X1 D1206 ( .Q(D1206_Q), .D(D5555_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D1205 ( .Q(D1205_Q), .D(D9833_Y), .CK(D9782_QN));
KC_DFFHQ_X1 D1204 ( .Q(D1204_Q), .D(D9833_Y), .CK(D11072_QN));
KC_DFFHQ_X1 D1203 ( .Q(D1203_Q), .D(D6952_Y), .CK(D4027_QN));
KC_DFFHQ_X1 D1202 ( .Q(D1202_Q), .D(D6956_Y), .CK(D4010_QN));
KC_DFFHQ_X1 D1201 ( .Q(D1201_Q), .D(D9833_Y), .CK(D10592_QN));
KC_DFFHQ_X1 D1200 ( .Q(D1200_Q), .D(D6952_Y), .CK(D4012_QN));
KC_DFFHQ_X1 D1199 ( .Q(D1199_Q), .D(D8572_Y), .CK(D11071_QN));
KC_DFFHQ_X1 D1142 ( .Q(D1142_Q), .D(D11994_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D1141 ( .Q(D1141_Q), .D(D10503_Y), .CK(D899_QN));
KC_DFFHQ_X1 D1140 ( .Q(D1140_Q), .D(D11995_Y), .CK(D112_QN));
KC_DFFHQ_X1 D1139 ( .Q(D1139_Q), .D(D11454_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D1138 ( .Q(D1138_Q), .D(D11454_Y), .CK(D112_QN));
KC_DFFHQ_X1 D1137 ( .Q(D1137_Q), .D(D10503_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D1136 ( .Q(D1136_Q), .D(D11453_Y), .CK(D112_QN));
KC_DFFHQ_X1 D1135 ( .Q(D1135_Q), .D(D11454_Y), .CK(D2286_QN));
KC_DFFHQ_X1 D1134 ( .Q(D1134_Q), .D(D11454_Y), .CK(D1120_QN));
KC_DFFHQ_X1 D1133 ( .Q(D1133_Q), .D(D1003_Y), .CK(D10876_QN));
KC_DFFHQ_X1 D1132 ( .Q(D1132_Q), .D(D6952_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D1131 ( .Q(D1131_Q), .D(D9767_Y), .CK(D2059_Y));
KC_DFFHQ_X1 D1130 ( .Q(D1130_Q), .D(D6957_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D1129 ( .Q(D1129_Q), .D(D6890_Y), .CK(D5462_QN));
KC_DFFHQ_X1 D1128 ( .Q(D1128_Q), .D(D5458_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D1127 ( .Q(D1127_Q), .D(D10480_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D1126 ( .Q(D1126_Q), .D(D1102_Y), .CK(D8441_Y));
KC_DFFHQ_X1 D1125 ( .Q(D1125_Q), .D(D6909_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D1124 ( .Q(D1124_Q), .D(D5456_Y), .CK(D1483_QN));
KC_DFFHQ_X1 D1123 ( .Q(D1123_Q), .D(D1101_Y), .CK(D10494_Y));
KC_DFFHQ_X1 D1122 ( .Q(D1122_Q), .D(D6956_Y), .CK(D4014_QN));
KC_DFFHQ_X1 D1121 ( .Q(D1121_Q), .D(D6956_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D1044 ( .Q(D1044_Q), .D(D11849_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D1043 ( .Q(D1043_Q), .D(D1007_Y), .CK(D10939_QN));
KC_DFFHQ_X1 D1042 ( .Q(D1042_Q), .D(D9696_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D1041 ( .Q(D1041_Q), .D(D11849_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D1040 ( .Q(D1040_Q), .D(D10414_Y), .CK(D11324_QN));
KC_DFFHQ_X1 D1039 ( .Q(D1039_Q), .D(D11852_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D1038 ( .Q(D1038_Q), .D(D11849_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D1037 ( .Q(D1037_Q), .D(D9696_Y), .CK(D2154_QN));
KC_DFFHQ_X1 D1036 ( .Q(D1036_Q), .D(D11847_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D1035 ( .Q(D1035_Q), .D(D11849_Y), .CK(D11910_QN));
KC_DFFHQ_X1 D1034 ( .Q(D1034_Q), .D(D11849_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D1033 ( .Q(D1033_Q), .D(D10414_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D1032 ( .Q(D1032_Q), .D(D9777_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D1031 ( .Q(D1031_Q), .D(D11384_Y), .CK(D1119_QN));
KC_DFFHQ_X1 D1030 ( .Q(D1030_Q), .D(D11383_Y), .CK(D11387_QN));
KC_DFFHQ_X1 D1029 ( .Q(D1029_Q), .D(D10414_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D1028 ( .Q(D1028_Q), .D(D9795_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D1027 ( .Q(D1027_Q), .D(D11454_Y), .CK(D11909_QN));
KC_DFFHQ_X1 D1026 ( .Q(D1026_Q), .D(D11454_Y), .CK(D1010_QN));
KC_DFFHQ_X1 D1025 ( .Q(D1025_Q), .D(D10502_Y), .CK(D1011_QN));
KC_DFFHQ_X1 D1024 ( .Q(D1024_Q), .D(D9697_Y), .CK(D10875_QN));
KC_DFFHQ_X1 D1023 ( .Q(D1023_Q), .D(D1618_Y), .CK(D891_QN));
KC_DFFHQ_X1 D1022 ( .Q(D1022_Q), .D(D9698_Y), .CK(D2150_QN));
KC_DFFHQ_X1 D1021 ( .Q(D1021_Q), .D(D10873_Y), .CK(D898_QN));
KC_DFFHQ_X1 D1020 ( .Q(D1020_Q), .D(D9698_Y), .CK(D900_QN));
KC_DFFHQ_X1 D1019 ( .Q(D1019_Q), .D(D1619_Y), .CK(D3867_QN));
KC_DFFHQ_X1 D1018 ( .Q(D1018_Q), .D(D9702_Y), .CK(D898_QN));
KC_DFFHQ_X1 D1017 ( .Q(D1017_Q), .D(D5457_Y), .CK(D891_QN));
KC_DFFHQ_X1 D1016 ( .Q(D1016_Q), .D(D9777_Y), .CK(D898_QN));
KC_DFFHQ_X1 D1015 ( .Q(D1015_Q), .D(D9702_Y), .CK(D10416_QN));
KC_DFFHQ_X1 D1014 ( .Q(D1014_Q), .D(D6273_Y), .CK(D891_QN));
KC_DFFHQ_X1 D1013 ( .Q(D1013_Q), .D(D9795_Y), .CK(D898_QN));
KC_DFFHQ_X1 D1012 ( .Q(D1012_Q), .D(D6891_Y), .CK(D893_QN));
KC_DFFHQ_X1 D920 ( .Q(D920_Q), .D(D11854_Y), .CK(D11913_QN));
KC_DFFHQ_X1 D919 ( .Q(D919_Q), .D(D11854_Y), .CK(D11911_QN));
KC_DFFHQ_X1 D918 ( .Q(D918_Q), .D(D11854_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D917 ( .Q(D917_Q), .D(D10873_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D916 ( .Q(D916_Q), .D(D11846_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D915 ( .Q(D915_Q), .D(D11854_Y), .CK(D12448_QN));
KC_DFFHQ_X1 D914 ( .Q(D914_Q), .D(D1007_Y), .CK(D901_QN));
KC_DFFHQ_X1 D913 ( .Q(D913_Q), .D(D10873_Y), .CK(D10878_QN));
KC_DFFHQ_X1 D912 ( .Q(D912_Q), .D(D11851_Y), .CK(D2287_QN));
KC_DFFHQ_X1 D911 ( .Q(D911_Q), .D(D9696_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D910 ( .Q(D910_Q), .D(D11854_Y), .CK(D11914_QN));
KC_DFFHQ_X1 D909 ( .Q(D909_Q), .D(D11854_Y), .CK(D11915_QN));
KC_DFFHQ_X1 D908 ( .Q(D908_Q), .D(D1113_Y), .CK(D11323_QN));
KC_DFFHQ_X1 D907 ( .Q(D907_Q), .D(D6805_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D906 ( .Q(D906_Q), .D(D5386_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D905 ( .Q(D905_Q), .D(D9695_Y), .CK(D10879_QN));
KC_DFFHQ_X1 D904 ( .Q(D904_Q), .D(D9695_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D903 ( .Q(D903_Q), .D(D6764_Y), .CK(D884_Y));
KC_DFFHQ_X1 D902 ( .Q(D902_Q), .D(D1002_Y), .CK(D6816_QN));
KC_DFFHQ_X1 D810 ( .Q(D810_Q), .D(D2283_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D809 ( .Q(D809_Q), .D(D11784_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D808 ( .Q(D808_Q), .D(D11254_Y), .CK(D11166_QN));
KC_DFFHQ_X1 D807 ( .Q(D807_Q), .D(D11778_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D806 ( .Q(D806_Q), .D(D11784_Y), .CK(D11167_QN));
KC_DFFHQ_X1 D805 ( .Q(D805_Q), .D(D11254_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D804 ( .Q(D804_Q), .D(D11778_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D803 ( .Q(D803_Q), .D(D11784_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D802 ( .Q(D802_Q), .D(D11779_Y), .CK(D660_QN));
KC_DFFHQ_X1 D801 ( .Q(D801_Q), .D(D11254_Y), .CK(D11174_QN));
KC_DFFHQ_X1 D800 ( .Q(D800_Q), .D(D11779_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D799 ( .Q(D799_Q), .D(D2283_Y), .CK(D660_QN));
KC_DFFHQ_X1 D798 ( .Q(D798_Q), .D(D2283_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D797 ( .Q(D797_Q), .D(D11229_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D796 ( .Q(D796_Q), .D(D738_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D795 ( .Q(D795_Q), .D(D6742_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D794 ( .Q(D794_Q), .D(D6731_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D793 ( .Q(D793_Q), .D(D6731_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D792 ( .Q(D792_Q), .D(D5298_Y), .CK(D3872_QN));
KC_DFFHQ_X1 D791 ( .Q(D791_Q), .D(D6805_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D790 ( .Q(D790_Q), .D(D5300_Y), .CK(D3871_QN));
KC_DFFHQ_X1 D789 ( .Q(D789_Q), .D(D8178_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D788 ( .Q(D788_Q), .D(D1759_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D787 ( .Q(D787_Q), .D(D5381_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D786 ( .Q(D786_Q), .D(D5382_Y), .CK(D3873_QN));
KC_DFFHQ_X1 D785 ( .Q(D785_Q), .D(D8208_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D784 ( .Q(D784_Q), .D(D8206_Y), .CK(D884_Y));
KC_DFFHQ_X1 D730 ( .Q(D730_Q), .D(D11253_Y), .CK(D11164_QN));
KC_DFFHQ_X1 D729 ( .Q(D729_Q), .D(D11785_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D728 ( .Q(D728_Q), .D(D11786_Y), .CK(D11165_QN));
KC_DFFHQ_X1 D690 ( .Q(D690_Q), .D(D11786_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D689 ( .Q(D689_Q), .D(D11253_Y), .CK(D11168_QN));
KC_DFFHQ_X1 D688 ( .Q(D688_Q), .D(D10824_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D687 ( .Q(D687_Q), .D(D11787_Y), .CK(D660_QN));
KC_DFFHQ_X1 D686 ( .Q(D686_Q), .D(D834_Y), .CK(D11170_QN));
KC_DFFHQ_X1 D685 ( .Q(D685_Q), .D(D834_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D684 ( .Q(D684_Q), .D(D11785_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D683 ( .Q(D683_Q), .D(D11784_Y), .CK(D718_QN));
KC_DFFHQ_X1 D682 ( .Q(D682_Q), .D(D11252_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D681 ( .Q(D681_Q), .D(D11783_Y), .CK(D11714_QN));
KC_DFFHQ_X1 D680 ( .Q(D680_Q), .D(D11254_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D679 ( .Q(D679_Q), .D(D10823_Y), .CK(D11169_QN));
KC_DFFHQ_X1 D678 ( .Q(D678_Q), .D(D11783_Y), .CK(D11173_QN));
KC_DFFHQ_X1 D677 ( .Q(D677_Q), .D(D11784_Y), .CK(D660_QN));
KC_DFFHQ_X1 D676 ( .Q(D676_Q), .D(D8129_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D675 ( .Q(D675_Q), .D(D576_Y), .CK(D655_QN));
KC_DFFHQ_X1 D674 ( .Q(D674_Q), .D(D8114_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D673 ( .Q(D673_Q), .D(D576_Y), .CK(D5220_QN));
KC_DFFHQ_X1 D672 ( .Q(D672_Q), .D(D8126_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D671 ( .Q(D671_Q), .D(D1760_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D670 ( .Q(D670_Q), .D(D6649_Y), .CK(D3723_QN));
KC_DFFHQ_X1 D669 ( .Q(D669_Q), .D(D8122_Y), .CK(D9448_Y));
KC_DFFHQ_X1 D668 ( .Q(D668_Q), .D(D6649_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D667 ( .Q(D667_Q), .D(D5298_Y), .CK(D1486_QN));
KC_DFFHQ_X1 D666 ( .Q(D666_Q), .D(D6645_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D665 ( .Q(D665_Q), .D(D5300_Y), .CK(D1485_QN));
KC_DFFHQ_X1 D664 ( .Q(D664_Q), .D(D8132_Y), .CK(D6735_Y));
KC_DFFHQ_X1 D663 ( .Q(D663_Q), .D(D6742_Y), .CK(D5219_QN));
KC_DFFHQ_X1 D662 ( .Q(D662_Q), .D(D5300_Y), .CK(D894_QN));
KC_DFFHQ_X1 D599 ( .Q(D599_Q), .D(D11779_Y), .CK(D661_QN));
KC_DFFHQ_X1 D598 ( .Q(D598_Q), .D(D6614_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D597 ( .Q(D597_Q), .D(D6614_Y), .CK(D5183_QN));
KC_DFFHQ_X1 D596 ( .Q(D596_Q), .D(D580_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D595 ( .Q(D595_Q), .D(D8059_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D594 ( .Q(D594_Q), .D(D6613_Y), .CK(D587_QN));
KC_DFFHQ_X1 D593 ( .Q(D593_Q), .D(D6613_Y), .CK(D586_QN));
KC_DFFHQ_X1 D592 ( .Q(D592_Q), .D(D579_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D591 ( .Q(D591_Q), .D(D6614_Y), .CK(D3669_QN));
KC_DFFHQ_X1 D590 ( .Q(D590_Q), .D(D8059_Y), .CK(D5184_QN));
KC_DFFHQ_X1 D589 ( .Q(D589_Q), .D(D6613_Y), .CK(D3670_QN));
KC_DFFHQ_X1 D527 ( .Q(D527_Q), .D(D11254_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D526 ( .Q(D526_Q), .D(D11252_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D525 ( .Q(D525_Q), .D(D10823_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D524 ( .Q(D524_Q), .D(D537_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D523 ( .Q(D523_Q), .D(D489_Y), .CK(D6538_QN));
KC_DFFHQ_X1 D522 ( .Q(D522_Q), .D(D5116_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D521 ( .Q(D521_Q), .D(D7976_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D520 ( .Q(D520_Q), .D(D5114_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D519 ( .Q(D519_Q), .D(D6532_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D518 ( .Q(D518_Q), .D(D3609_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D517 ( .Q(D517_Q), .D(D7977_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D516 ( .Q(D516_Q), .D(D5110_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D515 ( .Q(D515_Q), .D(D6526_Y), .CK(D6534_Y));
KC_DFFHQ_X1 D514 ( .Q(D514_Q), .D(D5103_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D513 ( .Q(D513_Q), .D(D498_Y), .CK(D6525_Y));
KC_DFFHQ_X1 D512 ( .Q(D512_Q), .D(D5109_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D480 ( .Q(D480_Q), .D(D7844_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D479 ( .Q(D479_Q), .D(D7879_Y), .CK(D6471_QN));
KC_DFFHQ_X1 D446 ( .Q(D446_Q), .D(D6366_Y), .CK(D6374_QN));
KC_DFFHQ_X1 D445 ( .Q(D445_Q), .D(D6364_Y), .CK(D6374_QN));
KC_DFFHQ_X1 D444 ( .Q(D444_Q), .D(D6403_Y), .CK(D6374_QN));
KC_DFFHQ_X1 D137 ( .Q(D137_Q), .D(D11778_Y), .CK(D11712_QN));
KC_DFFHQ_X1 D136 ( .Q(D136_Q), .D(D11190_Y), .CK(D10938_Y));
KC_DFFHQ_X1 D135 ( .Q(D135_Q), .D(D743_Y), .CK(D2211_Y));
KC_DFFHQ_X1 D134 ( .Q(D134_Q), .D(D11854_Y), .CK(D12447_QN));
KC_DFFHQ_X1 D133 ( .Q(D133_Q), .D(D9696_Y), .CK(D10345_QN));
KC_DFFHQ_X1 D132 ( .Q(D132_Q), .D(D11966_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D131 ( .Q(D131_Q), .D(D11503_Y), .CK(D10411_Y));
KC_DFFHQ_X1 D130 ( .Q(D130_Q), .D(D12055_Y), .CK(D11576_QN));
KC_DFFHQ_X1 D129 ( .Q(D129_Q), .D(D11477_Y), .CK(D11583_QN));
KC_DFFHQ_X1 D128 ( .Q(D128_Q), .D(D11993_Y), .CK(D12571_QN));
KC_DFFHQ_X1 D127 ( .Q(D127_Q), .D(D10824_Y), .CK(D11115_QN));
KC_DFFHQ_X1 D126 ( .Q(D126_Q), .D(D11786_Y), .CK(D661_QN));
KC_DFFHQ_X1 D125 ( .Q(D125_Q), .D(D1810_Y), .CK(D6538_QN));
KC_DFFHQ_X1 D124 ( .Q(D124_Q), .D(D5122_Y), .CK(D6468_QN));
KC_DFFHQ_X1 D123 ( .Q(D123_Q), .D(D5100_Y), .CK(D1631_QN));
KC_DFFHQ_X1 D122 ( .Q(D122_Q), .D(D8573_Y), .CK(D11069_QN));
KC_DFFHQ_X1 D121 ( .Q(D121_Q), .D(D8580_Y), .CK(D4013_QN));
KC_DFFHQ_X1 D120 ( .Q(D120_Q), .D(D5555_Y), .CK(D1196_QN));
KC_DFFHQ_X1 D119 ( .Q(D119_Q), .D(D5381_Y), .CK(D894_QN));
KC_DFFHQ_X1 D118 ( .Q(D118_Q), .D(D1002_Y), .CK(D6817_QN));
KC_DFFHQ_X1 D117 ( .Q(D117_Q), .D(D6797_Y), .CK(D893_QN));
KC_DFFHQ_X1 D115 ( .Q(D115_Q), .D(D6994_Y), .CK(D6954_Y));
KC_DFFHQ_X1 D114 ( .Q(D114_Q), .D(D6952_Y), .CK(D1487_QN));
KC_DFFHQ_X1 D113 ( .Q(D113_Q), .D(D6957_Y), .CK(D4015_QN));
KC_DFFHQ_X1 D116 ( .Q(D116_Q), .D(D10472_Y), .CK(D10494_Y));
KC_MXI2_X2 D16456 ( .Y(D16456_Y), .A(D16431_Y), .B(D16424_Y),     .S0(D16443_Y));
KC_MXI2_X2 D16221 ( .Y(D16221_Y), .A(D10126_Y), .B(D16401_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16220 ( .Y(D16220_Y), .A(D2171_Y), .B(D959_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16219 ( .Y(D16219_Y), .A(D10166_Y), .B(D2685_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16218 ( .Y(D16218_Y), .A(D10171_Y), .B(D16243_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16217 ( .Y(D16217_Y), .A(D10189_Y), .B(D776_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16216 ( .Y(D16216_Y), .A(D10634_Y), .B(D16371_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16215 ( .Y(D16215_Y), .A(D10175_Y), .B(D963_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16213 ( .Y(D16213_Y), .A(D14512_Y), .B(D964_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16212 ( .Y(D16212_Y), .A(D14508_Y), .B(D16344_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16211 ( .Y(D16211_Y), .A(D10112_Y), .B(D2686_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16210 ( .Y(D16210_Y), .A(D10188_Y), .B(D15957_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16209 ( .Y(D16209_Y), .A(D502_Y), .B(D16402_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16208 ( .Y(D16208_Y), .A(D15249_Y), .B(D16302_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16207 ( .Y(D16207_Y), .A(D14511_Y), .B(D16343_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16206 ( .Y(D16206_Y), .A(D10172_Y), .B(D16244_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16205 ( .Y(D16205_Y), .A(D10150_Y), .B(D16339_Y),     .S0(D13186_Y));
KC_MXI2_X2 D16204 ( .Y(D16204_Y), .A(D16224_Y), .B(D16193_Y),     .S0(D16242_Q));
KC_MXI2_X2 D16163 ( .Y(D16163_Y), .A(D16115_Y), .B(D16161_Y),     .S0(D14573_Y));
KC_MXI2_X2 D16162 ( .Y(D16162_Y), .A(D14510_Y), .B(D16367_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16161 ( .Y(D16161_Y), .A(D10167_Y), .B(D16335_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16160 ( .Y(D16160_Y), .A(D16103_Y), .B(D16148_Y),     .S0(D15447_Y));
KC_MXI2_X2 D16159 ( .Y(D16159_Y), .A(D10173_Y), .B(D16301_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16158 ( .Y(D16158_Y), .A(D10190_Y), .B(D2684_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16157 ( .Y(D16157_Y), .A(D10169_Y), .B(D16304_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16155 ( .Y(D16155_Y), .A(D16037_Y), .B(D2591_Y),     .S0(D16102_Y));
KC_MXI2_X2 D16153 ( .Y(D16153_Y), .A(D12141_Y), .B(D16303_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16152 ( .Y(D16152_Y), .A(D10110_Y), .B(D16300_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16151 ( .Y(D16151_Y), .A(D10113_Y), .B(D1249_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16150 ( .Y(D16150_Y), .A(D10114_Y), .B(D16368_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16149 ( .Y(D16149_Y), .A(D14509_Y), .B(D16370_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16148 ( .Y(D16148_Y), .A(D10170_Y), .B(D16366_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16146 ( .Y(D16146_Y), .A(D10168_Y), .B(D2687_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16145 ( .Y(D16145_Y), .A(D10174_Y), .B(D16338_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16144 ( .Y(D16144_Y), .A(D10165_Y), .B(D15956_Y),     .S0(D16195_Y));
KC_MXI2_X2 D16142 ( .Y(D16142_Y), .A(D16161_Y), .B(D16115_Y),     .S0(D15434_Y));
KC_MXI2_X2 D16141 ( .Y(D16141_Y), .A(D16103_Y), .B(D16148_Y),     .S0(D16157_Y));
KC_MXI2_X2 D16099 ( .Y(D16099_Y), .A(D10189_Y), .B(D16099_B),     .S0(D16016_Y));
KC_MXI2_X2 D16084 ( .Y(D16084_Y), .A(D13908_Q), .B(D16084_B),     .S0(D16016_Y));
KC_MXI2_X2 D16083 ( .Y(D16083_Y), .A(D13195_Q), .B(D16083_B),     .S0(D16016_Y));
KC_MXI2_X2 D16081 ( .Y(D16081_Y), .A(D10188_Y), .B(D16081_B),     .S0(D16016_Y));
KC_MXI2_X2 D16080 ( .Y(D16080_Y), .A(D16061_Y), .B(D16033_Y),     .S0(D15421_Y));
KC_MXI2_X2 D16076 ( .Y(D16076_Y), .A(D14512_Y), .B(D16076_B),     .S0(D16016_Y));
KC_MXI2_X2 D16075 ( .Y(D16075_Y), .A(D10190_Y), .B(D16075_B),     .S0(D16016_Y));
KC_MXI2_X2 D16074 ( .Y(D16074_Y), .A(D10172_Y), .B(D16074_B),     .S0(D2525_Y));
KC_MXI2_X2 D16073 ( .Y(D16073_Y), .A(D13907_Q), .B(D16073_B),     .S0(D16016_Y));
KC_MXI2_X2 D16072 ( .Y(D16072_Y), .A(D16053_Y), .B(D16088_Y),     .S0(D16090_Y));
KC_MXI2_X2 D16071 ( .Y(D16071_Y), .A(D16049_Y), .B(D16084_Y),     .S0(D16076_Y));
KC_MXI2_X2 D16046 ( .Y(D16046_Y), .A(D10169_Y), .B(D16046_B),     .S0(D16016_Y));
KC_MXI2_X2 D16039 ( .Y(D16039_Y), .A(D10126_Y), .B(D16039_B),     .S0(D2525_Y));
KC_MXI2_X2 D16038 ( .Y(D16038_Y), .A(D10113_Y), .B(D16038_B),     .S0(D2525_Y));
KC_MXI2_X2 D16037 ( .Y(D16037_Y), .A(D502_Y), .B(D16037_B),     .S0(D2525_Y));
KC_MXI2_X2 D16036 ( .Y(D16036_Y), .A(D14509_Y), .B(D16036_B),     .S0(D2525_Y));
KC_MXI2_X2 D16035 ( .Y(D16035_Y), .A(D10150_Y), .B(D16035_B),     .S0(D2525_Y));
KC_MXI2_X2 D16034 ( .Y(D16034_Y), .A(D12141_Y), .B(D16034_B),     .S0(D2525_Y));
KC_MXI2_X2 D16033 ( .Y(D16033_Y), .A(D10173_Y), .B(D16033_B),     .S0(D2525_Y));
KC_MXI2_X2 D16032 ( .Y(D16032_Y), .A(D2137_Y), .B(D16032_B),     .S0(D2525_Y));
KC_MXI2_X2 D16031 ( .Y(D16031_Y), .A(D10171_Y), .B(D16031_B),     .S0(D16016_Y));
KC_MXI2_X2 D16030 ( .Y(D16030_Y), .A(D14511_Y), .B(D16030_B),     .S0(D2525_Y));
KC_MXI2_X2 D16029 ( .Y(D16029_Y), .A(D10170_Y), .B(D16029_B),     .S0(D2525_Y));
KC_MXI2_X2 D16028 ( .Y(D16028_Y), .A(D10167_Y), .B(D16028_B),     .S0(D16016_Y));
KC_MXI2_X2 D16027 ( .Y(D16027_Y), .A(D10174_Y), .B(D16027_B),     .S0(D16016_Y));
KC_MXI2_X2 D16026 ( .Y(D16026_Y), .A(D10110_Y), .B(D16026_B),     .S0(D16016_Y));
KC_MXI2_X2 D16025 ( .Y(D16025_Y), .A(D10165_Y), .B(D16025_B),     .S0(D16016_Y));
KC_MXI2_X2 D16024 ( .Y(D16024_Y), .A(D15249_Y), .B(D16024_B),     .S0(D2525_Y));
KC_MXI2_X2 D16023 ( .Y(D16023_Y), .A(D14508_Y), .B(D16023_B),     .S0(D2525_Y));
KC_MXI2_X2 D16022 ( .Y(D16022_Y), .A(D10112_Y), .B(D16022_B),     .S0(D2525_Y));
KC_MXI2_X2 D16021 ( .Y(D16021_Y), .A(D14510_Y), .B(D16021_B),     .S0(D2525_Y));
KC_MXI2_X2 D16020 ( .Y(D16020_Y), .A(D10175_Y), .B(D16020_B),     .S0(D16016_Y));
KC_MXI2_X2 D16019 ( .Y(D16019_Y), .A(D10168_Y), .B(D16019_B),     .S0(D16016_Y));
KC_MXI2_X2 D16018 ( .Y(D16018_Y), .A(D10114_Y), .B(D16018_B),     .S0(D16016_Y));
KC_MXI2_X2 D15989 ( .Y(D15989_Y), .A(D16011_Q), .B(D15961_Y),     .S0(D15993_Q));
KC_MXI2_X2 D15946 ( .Y(D15946_Y), .A(D16393_Q), .B(D15910_Y),     .S0(D16390_Q));
KC_MXI2_X2 D15945 ( .Y(D15945_Y), .A(D15884_Y), .B(D16385_Q),     .S0(D15883_Y));
KC_MXI2_X2 D15866 ( .Y(D15866_Y), .A(D15820_Y), .B(D16356_Q),     .S0(D15831_Y));
KC_MXI2_X2 D15788 ( .Y(D15788_Y), .A(D15669_Q), .B(D15739_Y),     .S0(D1077_Q));
KC_MXI2_X2 D15705 ( .Y(D15705_Y), .A(D15472_Y), .B(D2616_Y),     .S0(D15621_Y));
KC_MXI2_X2 D15667 ( .Y(D15667_Y), .A(D15485_Y), .B(D15484_Y),     .S0(D15637_Y));
KC_MXI2_X2 D15666 ( .Y(D15666_Y), .A(D15485_Y), .B(D15484_Y),     .S0(D15620_Y));
KC_MXI2_X2 D15665 ( .Y(D15665_Y), .A(D2606_Y), .B(D15466_Y),     .S0(D14845_Y));
KC_MXI2_X2 D15566 ( .Y(D15566_Y), .A(D15378_Y), .B(D15367_Y),     .S0(D15517_Y));
KC_MXI2_X2 D15565 ( .Y(D15565_Y), .A(D15359_Y), .B(D15362_Y),     .S0(D15521_Y));
KC_MXI2_X2 D15564 ( .Y(D15564_Y), .A(D15487_Y), .B(D1273_Y),     .S0(D16242_Q));
KC_MXI2_X2 D15452 ( .Y(D15452_Y), .A(D15378_Y), .B(D15367_Y),     .S0(D15514_Y));
KC_MXI2_X2 D15449 ( .Y(D15449_Y), .A(D15390_Y), .B(D16037_Y),     .S0(D15389_Y));
KC_MXI2_X2 D15447 ( .Y(D15447_Y), .A(D10111_Y), .B(D1248_Y),     .S0(D16195_Y));
KC_MXI2_X2 D15446 ( .Y(D15446_Y), .A(D15348_Y), .B(D15376_Y),     .S0(D14777_Y));
KC_MXI2_X2 D15445 ( .Y(D15445_Y), .A(D15364_Y), .B(D15361_Y),     .S0(D15527_Y));
KC_MXI2_X2 D15444 ( .Y(D15444_Y), .A(D15365_Y), .B(D15354_Y),     .S0(D15519_Y));
KC_MXI2_X2 D15328 ( .Y(D15328_Y), .A(D2636_Y), .B(D15291_Y),     .S0(D14373_Y));
KC_MXI2_X2 D15252 ( .Y(D15252_Y), .A(D10166_Y), .B(D15252_B),     .S0(D2525_Y));
KC_MXI2_X2 D15251 ( .Y(D15251_Y), .A(D10634_Y), .B(D15251_B),     .S0(D2525_Y));
KC_MXI2_X2 D15211 ( .Y(D15211_Y), .A(D15172_Y), .B(D15236_Q),     .S0(D15165_Y));
KC_MXI2_X2 D14868 ( .Y(D14868_Y), .A(D14878_Q), .B(D14727_Y),     .S0(D14814_Q));
KC_MXI2_X2 D14516 ( .Y(D14516_Y), .A(D14687_Q), .B(D14532_Y),     .S0(D12173_Y));
KC_MXI2_X2 D14473 ( .Y(D14473_Y), .A(D16014_Q), .B(D14408_Y),     .S0(D14493_Q));
KC_MXI2_X2 D14472 ( .Y(D14472_Y), .A(D14413_Y), .B(D1375_Q),     .S0(D14430_Y));
KC_MXI2_X2 D14235 ( .Y(D14235_Y), .A(D14239_Q), .B(D14212_Y),     .S0(D14246_Q));
KC_MXI2_X2 D14234 ( .Y(D14234_Y), .A(D13655_Y), .B(D14237_Q),     .S0(D14222_Y));
KC_MXI2_X2 D14159 ( .Y(D14159_Y), .A(D14170_Q), .B(D14016_Y),     .S0(D14117_Q));
KC_MXI2_X2 D14090 ( .Y(D14090_Y), .A(D12688_Q), .B(D13906_Y),     .S0(D14711_Y));
KC_MXI2_X2 D14089 ( .Y(D14089_Y), .A(D12682_Q), .B(D12689_Q),     .S0(D14711_Y));
KC_MXI2_X2 D14088 ( .Y(D14088_Y), .A(D13991_Q), .B(D697_Q),     .S0(D2478_Y));
KC_MXI2_X2 D14087 ( .Y(D14087_Y), .A(D692_Q), .B(D691_Q),     .S0(D2478_Y));
KC_MXI2_X2 D14086 ( .Y(D14086_Y), .A(D691_Q), .B(D692_Q),     .S0(D14711_Y));
KC_MXI2_X2 D14085 ( .Y(D14085_Y), .A(D13279_Q), .B(D13976_Y),     .S0(D14711_Y));
KC_MXI2_X2 D14084 ( .Y(D14084_Y), .A(D13200_Q), .B(D2511_Y),     .S0(D14711_Y));
KC_MXI2_X2 D14083 ( .Y(D14083_Y), .A(D13279_Q), .B(D13976_Y),     .S0(D14711_Y));
KC_MXI2_X2 D14082 ( .Y(D14082_Y), .A(D12686_Q), .B(D13209_Q),     .S0(D14711_Y));
KC_MXI2_X2 D14081 ( .Y(D14081_Y), .A(D697_Q), .B(D13991_Q),     .S0(D14711_Y));
KC_MXI2_X2 D14004 ( .Y(D14004_Y), .A(D13271_Q), .B(D13272_Q),     .S0(D2478_Y));
KC_MXI2_X2 D14002 ( .Y(D14002_Y), .A(D13202_Q), .B(D13199_Q),     .S0(D14711_Y));
KC_MXI2_X2 D14001 ( .Y(D14001_Y), .A(D13199_Q), .B(D13202_Q),     .S0(D2478_Y));
KC_MXI2_X2 D13987 ( .Y(D13987_Y), .A(D12684_Q), .B(D13210_Q),     .S0(D14711_Y));
KC_MXI2_X2 D13986 ( .Y(D13986_Y), .A(D13992_Q), .B(D13989_Q),     .S0(D2478_Y));
KC_MXI2_X2 D13985 ( .Y(D13985_Y), .A(D13272_Q), .B(D13271_Q),     .S0(D14711_Y));
KC_MXI2_X2 D13984 ( .Y(D13984_Y), .A(D13990_Q), .B(D13998_Q),     .S0(D2478_Y));
KC_MXI2_X2 D13983 ( .Y(D13983_Y), .A(D13998_Q), .B(D13990_Q),     .S0(D14711_Y));
KC_MXI2_X2 D13982 ( .Y(D13982_Y), .A(D13989_Q), .B(D13992_Q),     .S0(D14711_Y));
KC_MXI2_X2 D13854 ( .Y(D13854_Y), .A(D2498_Y), .B(D13872_Q),     .S0(D2505_Y));
KC_MXI2_X2 D13797 ( .Y(D13797_Y), .A(D1185_Y), .B(D13805_Q),     .S0(D14455_Y));
KC_MXI2_X2 D13755 ( .Y(D13755_Y), .A(D13670_Y), .B(D14299_Q),     .S0(D13673_Y));
KC_MXI2_X2 D13391 ( .Y(D13391_Y), .A(D12687_Q), .B(D13259_Y),     .S0(D14711_Y));
KC_MXI2_X2 D13389 ( .Y(D13389_Y), .A(D13324_Y), .B(D13368_Y),     .S0(D13332_Y));
KC_MXI2_X2 D13282 ( .Y(D13282_Y), .A(D13270_Q), .B(D13274_Q),     .S0(D13938_Y));
KC_MXI2_X2 D13169 ( .Y(D13169_Y), .A(D7730_Y), .B(D723_Q),     .S0(D13190_Y));
KC_MXI2_X2 D13168 ( .Y(D13168_Y), .A(D7784_Y), .B(D13285_Y),     .S0(D2466_Y));
KC_MXI2_X2 D13167 ( .Y(D13167_Y), .A(D7784_Y), .B(D13285_Y),     .S0(D2463_Y));
KC_MXI2_X2 D13166 ( .Y(D13166_Y), .A(D7730_Y), .B(D723_Q),     .S0(D13158_Y));
KC_MXI2_X2 D13165 ( .Y(D13165_Y), .A(D10159_Y), .B(D13288_Y),     .S0(D13159_Y));
KC_MXI2_X2 D12911 ( .Y(D12911_Y), .A(D15774_Y), .B(D12936_Q),     .S0(D12776_Y));
KC_MXI2_X2 D12910 ( .Y(D12910_Y), .A(D15765_Y), .B(D12923_Q),     .S0(D12776_Y));
KC_MXI2_X2 D12909 ( .Y(D12909_Y), .A(D15774_Y), .B(D12925_Q),     .S0(D12774_Y));
KC_MXI2_X2 D12908 ( .Y(D12908_Y), .A(D15765_Y), .B(D12924_Q),     .S0(D12774_Y));
KC_MXI2_X2 D12845 ( .Y(D12845_Y), .A(D12789_Y), .B(D12826_Y),     .S0(D12351_Q));
KC_MXI2_X2 D12844 ( .Y(D12844_Y), .A(D15774_Y), .B(D12853_Q),     .S0(D12778_Y));
KC_MXI2_X2 D12842 ( .Y(D12842_Y), .A(D15774_Y), .B(D12850_Q),     .S0(D12775_Y));
KC_MXI2_X2 D12841 ( .Y(D12841_Y), .A(D15765_Y), .B(D12852_Q),     .S0(D12778_Y));
KC_MXI2_X2 D12744 ( .Y(D12744_Y), .A(D2353_Y), .B(D7669_Y),     .S0(D699_Q));
KC_MXI2_X2 D12652 ( .Y(D12652_Y), .A(D10142_Y), .B(D13171_Y),     .S0(D12676_Y));
KC_MXI2_X2 D12651 ( .Y(D12651_Y), .A(D10161_Y), .B(D12863_Y),     .S0(D12626_Y));
KC_MXI2_X2 D12650 ( .Y(D12650_Y), .A(D10160_Y), .B(D12763_Y),     .S0(D12628_Y));
KC_MXI2_X2 D12649 ( .Y(D12649_Y), .A(D481_Y), .B(D12764_Y),     .S0(D12629_Y));
KC_MXI2_X2 D12648 ( .Y(D12648_Y), .A(D10158_Y), .B(D12761_Y),     .S0(D12632_Y));
KC_MXI2_X2 D12647 ( .Y(D12647_Y), .A(D10161_Y), .B(D12863_Y),     .S0(D2465_Y));
KC_MXI2_X2 D12646 ( .Y(D12646_Y), .A(D9269_Y), .B(D13289_Y),     .S0(D13161_Y));
KC_MXI2_X2 D12645 ( .Y(D12645_Y), .A(D10142_Y), .B(D13171_Y),     .S0(D13160_Y));
KC_MXI2_X2 D12644 ( .Y(D12644_Y), .A(D10160_Y), .B(D12763_Y),     .S0(D12656_Y));
KC_MXI2_X2 D12643 ( .Y(D12643_Y), .A(D7713_Y), .B(D12762_Y),     .S0(D12224_Y));
KC_MXI2_X2 D12642 ( .Y(D12642_Y), .A(D7713_Y), .B(D12762_Y),     .S0(D12674_Y));
KC_MXI2_X2 D12641 ( .Y(D12641_Y), .A(D481_Y), .B(D12764_Y),     .S0(D694_Q));
KC_MXI2_X2 D12640 ( .Y(D12640_Y), .A(D9266_Y), .B(D13287_Y),     .S0(D13211_Q));
KC_MXI2_X2 D12639 ( .Y(D12639_Y), .A(D9268_Y), .B(D13280_Q),     .S0(D13162_Y));
KC_MXI2_X2 D12638 ( .Y(D12638_Y), .A(D9268_Y), .B(D13280_Q),     .S0(D13163_Y));
KC_MXI2_X2 D12636 ( .Y(D12636_Y), .A(D10162_Y), .B(D724_Y),     .S0(D12225_Y));
KC_MXI2_X2 D12635 ( .Y(D12635_Y), .A(D9269_Y), .B(D13289_Y),     .S0(D13191_Y));
KC_MXI2_X2 D12634 ( .Y(D12634_Y), .A(D10157_Y), .B(D12300_Y),     .S0(D12630_Y));
KC_MXI2_X2 D12633 ( .Y(D12633_Y), .A(D10157_Y), .B(D12300_Y),     .S0(D12683_Q));
KC_MXI2_X2 D12233 ( .Y(D12233_Y), .A(D9354_Y), .B(D12301_Y),     .S0(D12227_Y));
KC_MXI2_X2 D12232 ( .Y(D12232_Y), .A(D11660_Y), .B(D4747_Y),     .S0(D12235_Q));
KC_MXI2_X2 D12231 ( .Y(D12231_Y), .A(D10177_Y), .B(D6287_Y),     .S0(D12278_Q));
KC_MXI2_X2 D12230 ( .Y(D12230_Y), .A(D9354_Y), .B(D12301_Y),     .S0(D2390_Q));
KC_MXI2_X2 D12229 ( .Y(D12229_Y), .A(D11655_Y), .B(D6281_Y),     .S0(D12237_Q));
KC_MXI2_X2 D12228 ( .Y(D12228_Y), .A(D11657_Y), .B(D392_Y),     .S0(D12234_Q));
KC_MXI2_X2 D12172 ( .Y(D12172_Y), .A(D7785_Y), .B(D725_Y),     .S0(D9379_Y));
KC_MXI2_X2 D12171 ( .Y(D12171_Y), .A(D12131_Y), .B(D548_Q),     .S0(D12137_Y));
KC_MXI2_X2 D11652 ( .Y(D11652_Y), .A(D12201_Y), .B(D11646_Y),     .S0(D585_Y));
KC_MXI2_X2 D10346 ( .Y(D10346_Y), .A(D10319_Y), .B(D10360_Q),     .S0(D10359_Q));
KC_MXI2_X2 D10290 ( .Y(D10290_Y), .A(D10243_Y), .B(D10294_Q),     .S0(D10300_Q));
KC_MXI2_X2 D10289 ( .Y(D10289_Y), .A(D10247_Y), .B(D10302_Q),     .S0(D10290_Y));
KC_MXI2_X2 D10288 ( .Y(D10288_Y), .A(D10246_Y), .B(D10301_Q),     .S0(D10303_Q));
KC_MXI2_X2 D10287 ( .Y(D10287_Y), .A(D10244_Y), .B(D10299_Q),     .S0(D825_Q));
KC_MXI2_X2 D10286 ( .Y(D10286_Y), .A(D10244_Y), .B(D10299_Q),     .S0(D9580_Q));
KC_MXI2_X2 D10215 ( .Y(D10215_Y), .A(D9424_Y), .B(D10225_Q),     .S0(D827_Q));
KC_MXI2_X2 D10214 ( .Y(D10214_Y), .A(D2118_Y), .B(D10296_Q),     .S0(D10311_Q));
KC_MXI2_X2 D10213 ( .Y(D10213_Y), .A(D2118_Y), .B(D10296_Q),     .S0(D10226_Q));
KC_MXI2_X2 D10212 ( .Y(D10212_Y), .A(D10243_Y), .B(D10294_Q),     .S0(D9581_Q));
KC_MXI2_X2 D10211 ( .Y(D10211_Y), .A(D10246_Y), .B(D10301_Q),     .S0(D701_Q));
KC_MXI2_X2 D10094 ( .Y(D10094_Y), .A(D10080_Y), .B(D379_Y),     .S0(D9104_Y));
KC_MXI2_X2 D9573 ( .Y(D9573_Y), .A(D9578_Q), .B(D9522_Y), .S0(D484_Q));
KC_MXI2_X2 D9572 ( .Y(D9572_Y), .A(D9576_Q), .B(D9528_Y),     .S0(D2092_Q));
KC_MXI2_X2 D9571 ( .Y(D9571_Y), .A(D9579_Q), .B(D9514_Y),     .S0(D9278_Q));
KC_MXI2_X2 D9568 ( .Y(D9568_Y), .A(D9583_Y), .B(D761_Y), .S0(D9524_Y));
KC_MXI2_X2 D9567 ( .Y(D9567_Y), .A(D9568_Y), .B(D9497_Y),     .S0(D9565_Y));
KC_MXI2_X2 D9565 ( .Y(D9565_Y), .A(D9542_Y), .B(D9497_Y),     .S0(D9583_Y));
KC_MXI2_X2 D9467 ( .Y(D9467_Y), .A(D9581_Q), .B(D9423_Y), .S0(D482_Q));
KC_MXI2_X2 D9466 ( .Y(D9466_Y), .A(D700_Q), .B(D1994_Y), .S0(D7894_Q));
KC_MXI2_X2 D9465 ( .Y(D9465_Y), .A(D9580_Q), .B(D9415_Y), .S0(D451_Q));
KC_MXI2_X2 D9464 ( .Y(D9464_Y), .A(D701_Q), .B(D9414_Y), .S0(D449_Q));
KC_MXI2_X2 D9463 ( .Y(D9463_Y), .A(D9423_Y), .B(D9581_Q),     .S0(D9470_Q));
KC_MXI2_X2 D9462 ( .Y(D9462_Y), .A(D10226_Q), .B(D9422_Y),     .S0(D483_Q));
KC_MXI2_X2 D9461 ( .Y(D9461_Y), .A(D10225_Q), .B(D9424_Y),     .S0(D9325_Q));
KC_MXI2_X2 D9460 ( .Y(D9460_Y), .A(D9414_Y), .B(D701_Q), .S0(D702_Q));
KC_MXI2_X2 D9459 ( .Y(D9459_Y), .A(D1994_Y), .B(D700_Q), .S0(D9454_Y));
KC_MXI2_X2 D9456 ( .Y(D9456_Y), .A(D9006_Y), .B(D8149_Q),     .S0(D8079_Y));
KC_MXI2_X2 D9455 ( .Y(D9455_Y), .A(D9470_Q), .B(D9406_Y),     .S0(D2094_Q));
KC_MXI2_X2 D9454 ( .Y(D9454_Y), .A(D9415_Y), .B(D9580_Q),     .S0(D10226_Q));
KC_MXI2_X2 D9453 ( .Y(D9453_Y), .A(D1994_Y), .B(D700_Q), .S0(D825_Q));
KC_MXI2_X2 D9263 ( .Y(D9263_Y), .A(D9300_Y), .B(D9255_Y),     .S0(D9245_Y));
KC_MXI2_X2 D9213 ( .Y(D9213_Y), .A(D9179_Y), .B(D9216_Q),     .S0(D7497_Y));
KC_MXI2_X2 D9145 ( .Y(D9145_Y), .A(D9118_Y), .B(D273_Y),     .S0(D13171_Y));
KC_MXI2_X2 D9091 ( .Y(D9091_Y), .A(D8973_Y), .B(D8899_Q),     .S0(D13288_Y));
KC_MXI2_X2 D9090 ( .Y(D9090_Y), .A(D9033_Y), .B(D8951_Q),     .S0(D8064_Y));
KC_MXI2_X2 D9011 ( .Y(D9011_Y), .A(D9017_Y), .B(D8896_Q),     .S0(D12763_Y));
KC_MXI2_X2 D9010 ( .Y(D9010_Y), .A(D10043_Y), .B(D8895_Q),     .S0(D724_Y));
KC_MXI2_X2 D9009 ( .Y(D9009_Y), .A(D9016_Y), .B(D326_Q),     .S0(D12762_Y));
KC_MXI2_X2 D9008 ( .Y(D9008_Y), .A(D9012_Y), .B(D2090_Q),     .S0(D13285_Y));
KC_MXI2_X2 D9007 ( .Y(D9007_Y), .A(D9015_Y), .B(D8897_Q),     .S0(D12764_Y));
KC_MXI2_X2 D9005 ( .Y(D9005_Y), .A(D9014_Y), .B(D9023_Q),     .S0(D8063_Y));
KC_MXI2_X2 D9004 ( .Y(D9004_Y), .A(D2086_Y), .B(D272_Y),     .S0(D13289_Y));
KC_MXI2_X2 D8947 ( .Y(D8947_Y), .A(D272_Y), .B(D2086_Y), .S0(D7_Y));
KC_MXI2_X2 D8945 ( .Y(D8945_Y), .A(D8904_Y), .B(D8954_Q),     .S0(D8937_Y));
KC_MXI2_X2 D8944 ( .Y(D8944_Y), .A(D8948_Y), .B(D8955_Q),     .S0(D12761_Y));
KC_MXI2_X2 D8943 ( .Y(D8943_Y), .A(D9013_Y), .B(D305_Q),     .S0(D12300_Y));
KC_MXI2_X2 D8892 ( .Y(D8892_Y), .A(D9012_Y), .B(D2090_Q),     .S0(D8859_Y));
KC_MXI2_X2 D8891 ( .Y(D8891_Y), .A(D9015_Y), .B(D8897_Q),     .S0(D8874_Y));
KC_MXI2_X2 D8890 ( .Y(D8890_Y), .A(D8948_Y), .B(D8955_Q), .S0(D245_Y));
KC_MXI2_X2 D8814 ( .Y(D8814_Y), .A(D8698_Y), .B(D8700_Y), .S0(D231_Q));
KC_MXI2_X2 D8811 ( .Y(D8811_Y), .A(D8810_Y), .B(D8814_Y),     .S0(D9984_Q));
KC_MXI2_X2 D8810 ( .Y(D8810_Y), .A(D8809_Y), .B(D8808_Y), .S0(D231_Q));
KC_MXI2_X2 D8809 ( .Y(D8809_Y), .A(D8823_Q), .B(D9981_Q),     .S0(D8825_Q));
KC_MXI2_X2 D8808 ( .Y(D8808_Y), .A(D233_Q), .B(D9980_Q), .S0(D8825_Q));
KC_MXI2_X2 D8700 ( .Y(D8700_Y), .A(D9950_Q), .B(D8712_Q),     .S0(D8825_Q));
KC_MXI2_X2 D8698 ( .Y(D8698_Y), .A(D227_Q), .B(D9941_Q), .S0(D8825_Q));
KC_MXI2_X2 D8537 ( .Y(D8537_Y), .A(D8548_Q), .B(D8493_Y),     .S0(D16775_Y));
KC_MXI2_X2 D8536 ( .Y(D8536_Y), .A(D115_Q), .B(D8481_Y), .S0(D6917_Y));
KC_MXI2_X2 D8535 ( .Y(D8535_Y), .A(D8546_Q), .B(D8497_Y),     .S0(D8496_Y));
KC_MXI2_X2 D8457 ( .Y(D8457_Y), .A(D8394_Y), .B(D8392_Y),     .S0(D8440_Y));
KC_MXI2_X2 D8327 ( .Y(D8327_Y), .A(D6783_Y), .B(D8330_Q),     .S0(D6699_Y));
KC_MXI2_X2 D8325 ( .Y(D8325_Y), .A(D8381_Y), .B(D1838_Y),     .S0(D8327_Y));
KC_MXI2_X2 D8236 ( .Y(D8236_Y), .A(D8191_Y), .B(D8244_Q),     .S0(D8245_Q));
KC_MXI2_X2 D8233 ( .Y(D8233_Y), .A(D1931_Q), .B(D1824_Y),     .S0(D8173_Y));
KC_MXI2_X2 D8144 ( .Y(D8144_Y), .A(D8145_Q), .B(D8121_Y),     .S0(D8189_Y));
KC_MXI2_X2 D8143 ( .Y(D8143_Y), .A(D8117_Y), .B(D8107_Y),     .S0(D8091_Y));
KC_MXI2_X2 D7965 ( .Y(D7965_Y), .A(D7943_Y), .B(D7921_Y),     .S0(D7888_Q));
KC_MXI2_X2 D7881 ( .Y(D7881_Y), .A(D7888_Q), .B(D7839_Y),     .S0(D7845_Y));
KC_MXI2_X2 D7729 ( .Y(D7729_Y), .A(D13171_Y), .B(D10142_Y),     .S0(D364_Q));
KC_MXI2_X2 D7728 ( .Y(D7728_Y), .A(D12300_Y), .B(D10157_Y),     .S0(D384_Q));
KC_MXI2_X2 D7726 ( .Y(D7726_Y), .A(D12863_Y), .B(D10161_Y),     .S0(D4639_Q));
KC_MXI2_X2 D7725 ( .Y(D7725_Y), .A(D13280_Q), .B(D9268_Y),     .S0(D429_Q));
KC_MXI2_X2 D7724 ( .Y(D7724_Y), .A(D13285_Y), .B(D7784_Y),     .S0(D427_Q));
KC_MXI2_X2 D7722 ( .Y(D7722_Y), .A(D12301_Y), .B(D9354_Y),     .S0(D395_Q));
KC_MXI2_X2 D7721 ( .Y(D7721_Y), .A(D9266_Y), .B(D13287_Y),     .S0(D430_Q));
KC_MXI2_X2 D7720 ( .Y(D7720_Y), .A(D12761_Y), .B(D10158_Y),     .S0(D6357_Q));
KC_MXI2_X2 D7719 ( .Y(D7719_Y), .A(D7680_Y), .B(D9205_Y),     .S0(D7696_Y));
KC_MXI2_X2 D7718 ( .Y(D7718_Y), .A(D13288_Y), .B(D10159_Y),     .S0(D418_Q));
KC_MXI2_X2 D7717 ( .Y(D7717_Y), .A(D12764_Y), .B(D481_Y),     .S0(D6359_Q));
KC_MXI2_X2 D7716 ( .Y(D7716_Y), .A(D12763_Y), .B(D10160_Y),     .S0(D7741_Q));
KC_MXI2_X2 D7715 ( .Y(D7715_Y), .A(D724_Y), .B(D10162_Y), .S0(D167_Q));
KC_MXI2_X2 D7714 ( .Y(D7714_Y), .A(D725_Y), .B(D7785_Y), .S0(D6345_Q));
KC_MXI2_X2 D7650 ( .Y(D7650_Y), .A(D13289_Y), .B(D9269_Y),     .S0(D4641_Q));
KC_MXI2_X2 D7529 ( .Y(D7529_Y), .A(D282_Y), .B(D7479_Q), .S0(D8062_Y));
KC_MXI2_X2 D7528 ( .Y(D7528_Y), .A(D10045_Y), .B(D7_Y), .S0(D12863_Y));
KC_MXI2_X2 D7527 ( .Y(D7527_Y), .A(D7422_Y), .B(D4522_Y),     .S0(D6239_Y));
KC_MXI2_X2 D7525 ( .Y(D7525_Y), .A(D7730_Y), .B(D723_Q), .S0(D8824_Q));
KC_MXI2_X2 D7519 ( .Y(D7519_Y), .A(D7514_Y), .B(D6185_Y),     .S0(D7571_Y));
KC_MXI2_X2 D7467 ( .Y(D7467_Y), .A(D4116_Y), .B(D7442_Y),     .S0(D12863_Y));
KC_MXI2_X2 D7465 ( .Y(D7465_Y), .A(D303_Q), .B(D8949_Y),     .S0(D12301_Y));
KC_MXI2_X2 D7388 ( .Y(D7388_Y), .A(D7317_Y), .B(D7383_Y),     .S0(D7399_Y));
KC_MXI2_X2 D7294 ( .Y(D7294_Y), .A(D9476_Y), .B(D7183_Y),     .S0(D7166_Y));
KC_MXI2_X2 D7293 ( .Y(D7293_Y), .A(D9479_Y), .B(D8749_Y),     .S0(D1887_Y));
KC_MXI2_X2 D7292 ( .Y(D7292_Y), .A(D7172_Y), .B(D9475_Y),     .S0(D7167_Y));
KC_MXI2_X2 D7291 ( .Y(D7291_Y), .A(D9481_Y), .B(D2027_Y),     .S0(D7180_Y));
KC_MXI2_X2 D7139 ( .Y(D7139_Y), .A(D192_Q), .B(D7112_Y), .S0(D7115_Y));
KC_MXI2_X2 D6961 ( .Y(D6961_Y), .A(D6965_Q), .B(D6936_Y),     .S0(D6932_Y));
KC_MXI2_X2 D6960 ( .Y(D6960_Y), .A(D6963_Q), .B(D6925_Y),     .S0(D16777_Y));
KC_MXI2_X2 D6959 ( .Y(D6959_Y), .A(D6962_Q), .B(D6922_Y),     .S0(D6913_Y));
KC_MXI2_X2 D6812 ( .Y(D6812_Y), .A(D8328_Q), .B(D6766_Y), .S0(D863_Y));
KC_MXI2_X2 D6336 ( .Y(D6336_Y), .A(D6303_Y), .B(D6330_Y),     .S0(D6314_Y));
KC_MXI2_X2 D6335 ( .Y(D6335_Y), .A(D7704_Y), .B(D7674_Y),     .S0(D10204_Y));
KC_MXI2_X2 D6256 ( .Y(D6256_Y), .A(D6274_Y), .B(D6265_Y),     .S0(D13173_Y));
KC_MXI2_X2 D6116 ( .Y(D6116_Y), .A(D6165_Y), .B(D6104_Y),     .S0(D6103_Y));
KC_MXI2_X2 D6072 ( .Y(D6072_Y), .A(D7480_Q), .B(D726_Y), .S0(D5983_Y));
KC_MXI2_X2 D5680 ( .Y(D5680_Y), .A(D5649_Y), .B(D4119_Q),     .S0(D4092_Y));
KC_MXI2_X2 D5077 ( .Y(D5077_Y), .A(D3584_Y), .B(D5069_Y),     .S0(D3484_Q));
KC_MXI2_X2 D5075 ( .Y(D5075_Y), .A(D6507_Y), .B(D3502_Y),     .S0(D5082_Y));
KC_MXI2_X2 D4959 ( .Y(D4959_Y), .A(D4964_Y), .B(D3378_Y),     .S0(D3599_Y));
KC_MXI2_X2 D4810 ( .Y(D4810_Y), .A(D4788_Y), .B(D4775_Y),     .S0(D4820_Q));
KC_MXI2_X2 D4809 ( .Y(D4809_Y), .A(D4765_Y), .B(D4761_Y),     .S0(D4818_Q));
KC_MXI2_X2 D4805 ( .Y(D4805_Y), .A(D3372_Q), .B(D402_Y), .S0(D3311_Y));
KC_MXI2_X2 D4724 ( .Y(D4724_Y), .A(D1574_Y), .B(D2086_Y),     .S0(D3243_Y));
KC_MXI2_X2 D4723 ( .Y(D4723_Y), .A(D4684_Y), .B(D4666_Y), .S0(D391_Y));
KC_MXI2_X2 D4722 ( .Y(D4722_Y), .A(D4692_Y), .B(D3255_Y),     .S0(D4728_Q));
KC_MXI2_X2 D4631 ( .Y(D4631_Y), .A(D4602_Y), .B(D4552_Y),     .S0(D4497_Y));
KC_MXI2_X2 D4629 ( .Y(D4629_Y), .A(D4587_Y), .B(D4639_Q),     .S0(D4641_Q));
KC_MXI2_X2 D4477 ( .Y(D4477_Y), .A(D4434_Y), .B(D4484_Y),     .S0(D1717_Y));
KC_MXI2_X2 D4476 ( .Y(D4476_Y), .A(D4116_Y), .B(D4458_Y),     .S0(D5895_Y));
KC_MXI2_X2 D4475 ( .Y(D4475_Y), .A(D239_Q), .B(D4416_Y), .S0(D232_Q));
KC_MXI2_X2 D4474 ( .Y(D4474_Y), .A(D2878_Y), .B(D4434_Y),     .S0(D13289_Y));
KC_MXI2_X2 D4473 ( .Y(D4473_Y), .A(D165_Y), .B(D4417_Y), .S0(D4122_Q));
KC_MXI2_X2 D4472 ( .Y(D4472_Y), .A(D4470_Y), .B(D4449_Y),     .S0(D13171_Y));
KC_MXI2_X2 D4471 ( .Y(D4471_Y), .A(D8838_Y), .B(D1713_Y), .S0(D229_Q));
KC_MXI2_X2 D4469 ( .Y(D4469_Y), .A(D4150_Y), .B(D1787_Y),     .S0(D4136_Q));
KC_MXI2_X2 D4388 ( .Y(D4388_Y), .A(D4115_Y), .B(D255_Y), .S0(D4392_Y));
KC_MXI2_X2 D4387 ( .Y(D4387_Y), .A(D262_Y), .B(D4319_Y),     .S0(D13280_Q));
KC_MXI2_X2 D4386 ( .Y(D4386_Y), .A(D4270_Y), .B(D4286_Y),     .S0(D4302_Y));
KC_MXI2_X2 D4232 ( .Y(D4232_Y), .A(D4440_Y), .B(D5709_Y),     .S0(D5865_Y));
KC_MXI2_X2 D4230 ( .Y(D4230_Y), .A(D4187_Y), .B(D4246_Y),     .S0(D1582_Y));
KC_MXI2_X2 D4229 ( .Y(D4229_Y), .A(D4305_Y), .B(D4247_Y),     .S0(D1594_Y));
KC_MXI2_X2 D4228 ( .Y(D4228_Y), .A(D228_Q), .B(D4412_Y), .S0(D4119_Q));
KC_MXI2_X2 D4227 ( .Y(D4227_Y), .A(D4235_Q), .B(D4294_Y),     .S0(D4121_Q));
KC_MXI2_X2 D4114 ( .Y(D4114_Y), .A(D4096_Y), .B(D4118_Q),     .S0(D4095_Y));
KC_MXI2_X2 D4113 ( .Y(D4113_Y), .A(D4097_Y), .B(D4120_Q),     .S0(D4102_Y));
KC_MXI2_X2 D4112 ( .Y(D4112_Y), .A(D4122_Q), .B(D4094_Y), .S0(D176_Y));
KC_MXI2_X2 D3574 ( .Y(D3574_Y), .A(D3575_Q), .B(D3528_Y), .S0(D124_Q));
KC_MXI2_X2 D3478 ( .Y(D3478_Y), .A(D4893_Y), .B(D3516_Y), .S0(D69_Y));
KC_MXI2_X2 D3363 ( .Y(D3363_Y), .A(D3375_Q), .B(D3372_Q),     .S0(D3479_Y));
KC_MXI2_X2 D2994 ( .Y(D2994_Y), .A(D302_Q), .B(D4435_Y), .S0(D2708_Y));
KC_MXI2_X2 D2993 ( .Y(D2993_Y), .A(D3004_Q), .B(D2947_Y),     .S0(D2712_Y));
KC_MXI2_X2 D2992 ( .Y(D2992_Y), .A(D301_Q), .B(D2936_Y), .S0(D2711_Y));
KC_MXI2_X2 D2990 ( .Y(D2990_Y), .A(D2910_Y), .B(D2953_Y),     .S0(D2982_Y));
KC_MXI2_X2 D2988 ( .Y(D2988_Y), .A(D2816_Q), .B(D2848_Y),     .S0(D3082_Q));
KC_MXI2_X2 D2987 ( .Y(D2987_Y), .A(D2848_Y), .B(D2816_Q),     .S0(D1514_Q));
KC_MXI2_X2 D2986 ( .Y(D2986_Y), .A(D2848_Y), .B(D2816_Q),     .S0(D3093_Q));
KC_MXI2_X2 D2985 ( .Y(D2985_Y), .A(D2848_Y), .B(D2816_Q), .S0(D325_Q));
KC_MXI2_X2 D2879 ( .Y(D2879_Y), .A(D2844_Y), .B(D2737_Y),     .S0(D2846_Y));
KC_MXI2_X2 D2809 ( .Y(D2809_Y), .A(D2895_Y), .B(D2772_Y),     .S0(D2767_Y));
KC_MXI2_X2 D2673 ( .Y(D2673_Y), .A(D16083_Y), .B(D2653_Y),     .S0(D16028_Y));
KC_MXI2_X2 D2671 ( .Y(D2671_Y), .A(D618_Q), .B(D2671_B),     .S0(D16016_Y));
KC_MXI2_X2 D2670 ( .Y(D2670_Y), .A(D2171_Y), .B(D2670_B),     .S0(D16016_Y));
KC_MXI2_X2 D2668 ( .Y(D2668_Y), .A(D13921_Q), .B(D2668_B),     .S0(D16016_Y));
KC_MXI2_X2 D2667 ( .Y(D2667_Y), .A(D530_Q), .B(D2667_B),     .S0(D16016_Y));
KC_MXI2_X2 D2636 ( .Y(D2636_Y), .A(D13909_Q), .B(D2636_B),     .S0(D2525_Y));
KC_MXI2_X2 D2635 ( .Y(D2635_Y), .A(D15480_Y), .B(D15470_Y),     .S0(D15632_Y));
KC_MXI2_X2 D2634 ( .Y(D2634_Y), .A(D15479_Y), .B(D15468_Y),     .S0(D14863_Y));
KC_MXI2_X2 D2514 ( .Y(D2514_Y), .A(D13208_Q), .B(D13197_Q),     .S0(D2478_Y));
KC_MXI2_X2 D2400 ( .Y(D2400_Y), .A(D15765_Y), .B(D12917_Q),     .S0(D12775_Y));
KC_MXI2_X2 D2342 ( .Y(D2342_Y), .A(D7785_Y), .B(D725_Y),     .S0(D12675_Y));
KC_MXI2_X2 D2151 ( .Y(D2151_Y), .A(D10247_Y), .B(D10302_Q),     .S0(D10225_Q));
KC_MXI2_X2 D2077 ( .Y(D2077_Y), .A(D8904_Y), .B(D8954_Q),     .S0(D13280_Q));
KC_MXI2_X2 D2076 ( .Y(D2076_Y), .A(D8950_Y), .B(D151_Q),     .S0(D13287_Y));
KC_MXI2_X2 D2075 ( .Y(D2075_Y), .A(D8908_Y), .B(D334_Q), .S0(D8068_Y));
KC_MXI2_X2 D2074 ( .Y(D2074_Y), .A(D702_Q), .B(D10196_Y),     .S0(D2093_Q));
KC_MXI2_X2 D2073 ( .Y(D2073_Y), .A(D1994_Y), .B(D700_Q), .S0(D9531_Y));
KC_MXI2_X2 D1926 ( .Y(D1926_Y), .A(D1873_Y), .B(D7361_Y),     .S0(D7533_Q));
KC_MXI2_X2 D1924 ( .Y(D1924_Y), .A(D7449_Y), .B(D4499_Y),     .S0(D6239_Y));
KC_MXI2_X2 D1922 ( .Y(D1922_Y), .A(D538_Q), .B(D613_Q), .S0(D7973_Q));
KC_MXI2_X2 D1772 ( .Y(D1772_Y), .A(D6079_Y), .B(D4521_Y),     .S0(D6239_Y));
KC_MXI2_X2 D1632 ( .Y(D1632_Y), .A(D1629_Y), .B(D4306_Y), .S0(D723_Q));
KC_MXI2_X2 D1630 ( .Y(D1630_Y), .A(D4547_Y), .B(D4134_Y),     .S0(D4128_Y));
KC_MXI2_X2 D1491 ( .Y(D1491_Y), .A(D2848_Y), .B(D2816_Q), .S0(D150_Q));
KC_MXI2_X2 D1490 ( .Y(D1490_Y), .A(D2848_Y), .B(D2816_Q),     .S0(D3083_Q));
KC_MXI2_X2 D1489 ( .Y(D1489_Y), .A(D2816_Q), .B(D2848_Y),     .S0(D3081_Q));
KC_MXI2_X2 D1488 ( .Y(D1488_Y), .A(D2848_Y), .B(D2816_Q),     .S0(D3077_Q));
KC_MXI2_X2 D1117 ( .Y(D1117_Y), .A(D2679_Q), .B(D16347_Y),     .S0(D16353_Q));
KC_MXI2_X2 D1116 ( .Y(D1116_Y), .A(D6877_Y), .B(D8393_Y),     .S0(D8535_Y));
KC_MXI2_X2 D1115 ( .Y(D1115_Y), .A(D8541_Q), .B(D8488_Y),     .S0(D16776_Y));
KC_MXI2_X2 D895 ( .Y(D895_Y), .A(D8381_Y), .B(D1838_Y), .S0(D6812_Y));
KC_MXI2_X2 D783 ( .Y(D783_Y), .A(D12351_Q), .B(D12321_Y),     .S0(D12350_Q));
KC_MXI2_X2 D778 ( .Y(D778_Y), .A(D12681_Q), .B(D13203_Q),     .S0(D14711_Y));
KC_MXI2_X2 D777 ( .Y(D777_Y), .A(D12685_Q), .B(D13974_Y),     .S0(D14711_Y));
KC_MXI2_X2 D659 ( .Y(D659_Y), .A(D2137_Y), .B(D15710_Y),     .S0(D16195_Y));
KC_MXI2_X2 D658 ( .Y(D658_Y), .A(D13226_Y), .B(D12718_Y),     .S0(D13268_Q));
KC_MXI2_X2 D511 ( .Y(D511_Y), .A(D10162_Y), .B(D724_Y), .S0(D12680_Q));
KC_MXI2_X2 D510 ( .Y(D510_Y), .A(D10158_Y), .B(D12761_Y),     .S0(D12627_Y));
KC_MXI2_X2 D509 ( .Y(D509_Y), .A(D12178_Q), .B(D12132_Y),     .S0(D11183_Y));
KC_MXI2_X2 D505 ( .Y(D505_Y), .A(D10111_Y), .B(D505_B), .S0(D2525_Y));
KC_MXI2_X2 D379 ( .Y(D379_Y), .A(D10210_Y), .B(D727_Y), .S0(D10060_Q));
KC_MXI2_X2 D377 ( .Y(D377_Y), .A(D6211_Y), .B(D430_Q), .S0(D6357_Q));
KC_MXI2_X2 D351 ( .Y(D351_Y), .A(D13285_Y), .B(D7784_Y), .S0(D148_Q));
KC_MXI2_X2 D320 ( .Y(D320_Y), .A(D10044_Y), .B(D8898_Q), .S0(D725_Y));
KC_MXI2_X2 D295 ( .Y(D295_Y), .A(D8950_Y), .B(D151_Q), .S0(D283_Y));
KC_MXI2_X2 D225 ( .Y(D225_Y), .A(D4168_Y), .B(D4248_Y), .S0(D4278_Y));
KC_MXI2_X2 D110 ( .Y(D110_Y), .A(D569_Y), .B(D2668_Y), .S0(D584_Y));
KC_TLATHQN_X1 D16587 ( .D2(D16592_Y), .D1(D16582_Y), .QN(D16587_QN),     .GN(D1059_Y));
KC_TLATHQN_X1 D16515 ( .D2(D16525_Y), .D1(D16508_Y), .QN(D16515_QN),     .GN(D15867_Y));
KC_TLATHQN_X1 D15988 ( .D2(D16479_Y), .D1(D16446_Y), .QN(D15988_QN),     .GN(D2522_Y));
KC_TLATHQN_X1 D14162 ( .D2(D16766_Y), .D1(D2502_Y), .QN(D14162_QN),     .GN(D14177_Y));
KC_TLATHQN_X1 D14161 ( .D2(D2526_Y), .D1(D2491_Y), .QN(D14161_QN),     .GN(D833_Y));
KC_TLATHQN_X1 D14160 ( .D2(D14197_Y), .D1(D14126_Y), .QN(D14160_QN),     .GN(D833_Y));
KC_TLATHQN_X1 D14158 ( .D2(D16766_Y), .D1(D13405_Y), .QN(D14158_QN),     .GN(D14156_Y));
KC_TLATHQN_X1 D14157 ( .D2(D2526_Y), .D1(D2492_Y), .QN(D14157_QN),     .GN(D2458_Y));
KC_TLATHQN_X1 D14112 ( .D2(D14110_Y), .D1(D14116_Y), .QN(D14112_QN),     .GN(D14095_Y));
KC_TLATHQN_X1 D14080 ( .D2(D14110_Y), .D1(D14050_Y), .QN(D14080_QN),     .GN(D13404_Y));
KC_TLATHQN_X1 D13390 ( .D2(D14197_Y), .D1(D14129_Y), .QN(D13390_QN),     .GN(D2458_Y));
KC_TLATHQN_X1 D13388 ( .D2(D13408_Y), .D1(D13331_Y), .QN(D13388_QN),     .GN(D13404_Y));
KC_TLATHQN_X1 D13387 ( .D2(D16298_Y), .D1(D955_Y), .QN(D13387_QN),     .GN(D2458_Y));
KC_TLATHQN_X1 D13264 ( .D2(D13290_Y), .D1(D13247_Y), .QN(D13264_QN),     .GN(D13910_Y));
KC_TLATHQN_X1 D13263 ( .D2(D14006_Y), .D1(D13967_Y), .QN(D13263_QN),     .GN(D12859_Y));
KC_TLATHQN_X1 D13262 ( .D2(D13286_Y), .D1(D13241_Y), .QN(D13262_QN),     .GN(D15867_Y));
KC_TLATHQN_X1 D13261 ( .D2(D14110_Y), .D1(D14115_Y), .QN(D13261_QN),     .GN(D13276_Y));
KC_TLATHQN_X1 D13214 ( .D2(D13215_Y), .D1(D13187_Y), .QN(D13214_QN),     .GN(D13249_Y));
KC_TLATHQN_X1 D13193 ( .D2(D12691_Y), .D1(D2364_Y), .QN(D13193_QN),     .GN(D13205_Y));
KC_TLATHQN_X1 D12843 ( .D2(D12867_Y), .D1(D12824_Y), .QN(D12843_QN),     .GN(D12860_Y));
KC_TLATHQN_X1 D12746 ( .D2(D12758_Y), .D1(D12760_Y), .QN(D12746_QN),     .GN(D13249_Y));
KC_TLATHQN_X1 D12745 ( .D2(D12691_Y), .D1(D2377_Y), .QN(D12745_QN),     .GN(D12750_Y));
KC_TLATHQN_X1 D12742 ( .D2(D12867_Y), .D1(D12836_Y), .QN(D12742_QN),     .GN(D12860_Y));
KC_TLATHQN_X1 D12677 ( .D2(D12691_Y), .D1(D12667_Y), .QN(D12677_QN),     .GN(D12669_Y));
KC_TLATHQN_X1 D12571 ( .D2(D12128_Y), .D1(D11568_Y), .QN(D12571_QN),     .GN(D12084_Y));
KC_TLATHQN_X1 D12448 ( .D2(D11932_Y), .D1(D11893_Y), .QN(D12448_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D12447 ( .D2(D11932_Y), .D1(D11414_Y), .QN(D12447_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D12115 ( .D2(D12128_Y), .D1(D11588_Y), .QN(D12115_QN),     .GN(D12104_Y));
KC_TLATHQN_X1 D12114 ( .D2(D12129_Y), .D1(D11592_Y), .QN(D12114_QN),     .GN(D12104_Y));
KC_TLATHQN_X1 D12113 ( .D2(D12129_Y), .D1(D11587_Y), .QN(D12113_QN),     .GN(D11567_Y));
KC_TLATHQN_X1 D12085 ( .D2(D11590_Y), .D1(D11574_Y), .QN(D12085_QN),     .GN(D12084_Y));
KC_TLATHQN_X1 D12041 ( .D2(D11589_Y), .D1(D11569_Y), .QN(D12041_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D11916 ( .D2(D11933_Y), .D1(D11380_Y), .QN(D11916_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11915 ( .D2(D11931_Y), .D1(D11907_Y), .QN(D11915_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11914 ( .D2(D11932_Y), .D1(D11375_Y), .QN(D11914_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11913 ( .D2(D11931_Y), .D1(D11906_Y), .QN(D11913_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11912 ( .D2(D11931_Y), .D1(D1006_Y), .QN(D11912_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11911 ( .D2(D11932_Y), .D1(D11369_Y), .QN(D11911_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11910 ( .D2(D11931_Y), .D1(D11905_Y), .QN(D11910_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11909 ( .D2(D11932_Y), .D1(D11385_Y), .QN(D11909_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11714 ( .D2(D11676_Y), .D1(D11151_Y), .QN(D11714_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11713 ( .D2(D12240_Y), .D1(D12199_Y), .QN(D11713_QN),     .GN(D11711_Y));
KC_TLATHQN_X1 D11712 ( .D2(D11185_Y), .D1(D11700_Y), .QN(D11712_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11595 ( .D2(D11608_Y), .D1(D11556_Y), .QN(D11595_QN),     .GN(D12084_Y));
KC_TLATHQN_X1 D11583 ( .D2(D11589_Y), .D1(D11561_Y), .QN(D11583_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D11582 ( .D2(D11590_Y), .D1(D11573_Y), .QN(D11582_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D11581 ( .D2(D11589_Y), .D1(D11560_Y), .QN(D11581_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D11580 ( .D2(D11589_Y), .D1(D11570_Y), .QN(D11580_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D11579 ( .D2(D11589_Y), .D1(D11572_Y), .QN(D11579_QN),     .GN(D12104_Y));
KC_TLATHQN_X1 D11578 ( .D2(D11590_Y), .D1(D11571_Y), .QN(D11578_QN),     .GN(D12104_Y));
KC_TLATHQN_X1 D11577 ( .D2(D11590_Y), .D1(D11575_Y), .QN(D11577_QN),     .GN(D12084_Y));
KC_TLATHQN_X1 D11576 ( .D2(D11608_Y), .D1(D11545_Y), .QN(D11576_QN),     .GN(D12084_Y));
KC_TLATHQN_X1 D11387 ( .D2(D11933_Y), .D1(D11353_Y), .QN(D11387_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D11324 ( .D2(D10897_Y), .D1(D11348_Y), .QN(D11324_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D11323 ( .D2(D10897_Y), .D1(D11293_Y), .QN(D11323_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D11174 ( .D2(D11185_Y), .D1(D11161_Y), .QN(D11174_QN),     .GN(D11163_Y));
KC_TLATHQN_X1 D11173 ( .D2(D11184_Y), .D1(D2259_Y), .QN(D11173_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11171 ( .D2(D11185_Y), .D1(D11162_Y), .QN(D11171_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11170 ( .D2(D11186_Y), .D1(D11159_Y), .QN(D11170_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11169 ( .D2(D11186_Y), .D1(D11156_Y), .QN(D11169_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11168 ( .D2(D11186_Y), .D1(D11147_Y), .QN(D11168_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11167 ( .D2(D11279_Y), .D1(D11158_Y), .QN(D11167_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11166 ( .D2(D11186_Y), .D1(D11157_Y), .QN(D11166_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11165 ( .D2(D11279_Y), .D1(D11155_Y), .QN(D11165_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11164 ( .D2(D11186_Y), .D1(D11142_Y), .QN(D11164_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11134 ( .D2(D11117_Y), .D1(D11150_Y), .QN(D11134_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11115 ( .D2(D11117_Y), .D1(D2258_Y), .QN(D11115_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D11103 ( .D2(D11113_Y), .D1(D11099_Y), .QN(D11103_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D11102 ( .D2(D11113_Y), .D1(D11594_Y), .QN(D11102_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D11072 ( .D2(D11613_Y), .D1(D11559_Y), .QN(D11072_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D11071 ( .D2(D11089_Y), .D1(D11064_Y), .QN(D11071_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D11070 ( .D2(D11608_Y), .D1(D11558_Y), .QN(D11070_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D11069 ( .D2(D11089_Y), .D1(D1284_Y), .QN(D11069_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D11068 ( .D2(D11089_Y), .D1(D11562_Y), .QN(D11068_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D11067 ( .D2(D11613_Y), .D1(D11544_Y), .QN(D11067_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D11066 ( .D2(D11610_Y), .D1(D1338_Y), .QN(D11066_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D10939 ( .D2(D10897_Y), .D1(D11321_Y), .QN(D10939_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10879 ( .D2(D10895_Y), .D1(D10848_Y), .QN(D10879_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10878 ( .D2(D10898_Y), .D1(D10872_Y), .QN(D10878_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10877 ( .D2(D10896_Y), .D1(D10844_Y), .QN(D10877_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10876 ( .D2(D10896_Y), .D1(D10874_Y), .QN(D10876_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10875 ( .D2(D10898_Y), .D1(D10857_Y), .QN(D10875_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10593 ( .D2(D11610_Y), .D1(D1346_Y), .QN(D10593_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D10592 ( .D2(D11113_Y), .D1(D1267_Y), .QN(D10592_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D10543 ( .D2(D11088_Y), .D1(D2260_Y), .QN(D10543_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D10416 ( .D2(D10898_Y), .D1(D10866_Y), .QN(D10416_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10345 ( .D2(D10898_Y), .D1(D10894_Y), .QN(D10345_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D10107 ( .D2(D10129_Y), .D1(D431_Y), .QN(D10107_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D9783 ( .D2(D11088_Y), .D1(D11065_Y), .QN(D9783_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D9782 ( .D2(D11088_Y), .D1(D171_Y), .QN(D9782_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D9570 ( .D2(D9591_Y), .D1(D9585_Y), .QN(D9570_QN),     .GN(D534_Y));
KC_TLATHQN_X1 D9569 ( .D2(D9591_Y), .D1(D9560_Y), .QN(D9569_QN),     .GN(D10187_Y));
KC_TLATHQN_X1 D9468 ( .D2(D1973_Y), .D1(D7914_Y), .QN(D9468_QN),     .GN(D9474_Y));
KC_TLATHQN_X1 D9458 ( .D2(D8260_Y), .D1(D8174_Y), .QN(D9458_QN),     .GN(D2174_Q));
KC_TLATHQN_X1 D9212 ( .D2(D9229_Y), .D1(D411_Y), .QN(D9212_QN),     .GN(D9208_Y));
KC_TLATHQN_X1 D9211 ( .D2(D9229_Y), .D1(D9206_Y), .QN(D9211_QN),     .GN(D7520_Y));
KC_TLATHQN_X1 D9143 ( .D2(D9165_Y), .D1(D9103_Y), .QN(D9143_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D9142 ( .D2(D16757_Y), .D1(D71_Y), .QN(D9142_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D9141 ( .D2(D16757_Y), .D1(D9117_Y), .QN(D9141_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D9140 ( .D2(D9165_Y), .D1(D9112_Y), .QN(D9140_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D9139 ( .D2(D16757_Y), .D1(D9116_Y), .QN(D9139_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D8813 ( .D2(D8837_Y), .D1(D8736_Y), .QN(D8813_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D8235 ( .D2(D8263_Y), .D1(D8162_Y), .QN(D8235_QN),     .GN(D534_Y));
KC_TLATHQN_X1 D8142 ( .D2(D8167_Y), .D1(D8085_Y), .QN(D8142_QN),     .GN(D10187_Y));
KC_TLATHQN_X1 D7964 ( .D2(D7993_Y), .D1(D494_Y), .QN(D7964_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D7583 ( .D2(D7522_Y), .D1(D7550_Y), .QN(D7583_QN),     .GN(D7575_Y));
KC_TLATHQN_X1 D7530 ( .D2(D35_Y), .D1(D7498_Y), .QN(D7530_QN),     .GN(D7516_Y));
KC_TLATHQN_X1 D7524 ( .D2(D7561_Y), .D1(D7522_Y), .QN(D7524_QN),     .GN(VDD));
KC_TLATHQN_X1 D7518 ( .D2(D7561_Y), .D1(D1677_Y), .QN(D7518_QN),     .GN(VDD));
KC_TLATHQN_X1 D7468 ( .D2(D4_Y), .D1(D7457_Y), .QN(D7468_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D7466 ( .D2(D12_Y), .D1(D3_Y), .QN(D7466_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D7138 ( .D2(D7162_Y), .D1(D7378_Y), .QN(D7138_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D6817 ( .D2(D6832_Y), .D1(D6831_Y), .QN(D6817_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D6816 ( .D2(D6833_Y), .D1(D6776_Y), .QN(D6816_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D6815 ( .D2(D6832_Y), .D1(D6790_Y), .QN(D6815_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D6814 ( .D2(D6832_Y), .D1(D6779_Y), .QN(D6814_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D6811 ( .D2(D6832_Y), .D1(D6775_Y), .QN(D6811_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D6810 ( .D2(D6832_Y), .D1(D6778_Y), .QN(D6810_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D6538 ( .D2(D1819_Y), .D1(D1693_Y), .QN(D6538_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D6471 ( .D2(D6493_Y), .D1(D6495_Y), .QN(D6471_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D6468 ( .D2(D1673_Y), .D1(D5050_Y), .QN(D6468_QN),     .GN(D6461_Y));
KC_TLATHQN_X1 D6467 ( .D2(D1819_Y), .D1(D6420_Y), .QN(D6467_QN),     .GN(D536_Y));
KC_TLATHQN_X1 D6466 ( .D2(D6488_Y), .D1(D6456_Y), .QN(D6466_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D6374 ( .D2(D6488_Y), .D1(D6436_Y), .QN(D6374_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D6332 ( .D2(D6358_Y), .D1(D4789_Y), .QN(D6332_QN),     .GN(D6316_Y));
KC_TLATHQN_X1 D6258 ( .D2(D16147_Y), .D1(D6286_Y), .QN(D6258_QN),     .GN(D6242_Y));
KC_TLATHQN_X1 D5931 ( .D2(D5706_Y), .D1(D5875_Y), .QN(D5931_QN),     .GN(D7520_Y));
KC_TLATHQN_X1 D5800 ( .D2(D5701_Y), .D1(D5854_Y), .QN(D5800_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D5679 ( .D2(D5701_Y), .D1(D5919_Y), .QN(D5679_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D5559 ( .D2(D4031_Y), .D1(D3990_Y), .QN(D5559_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D5462 ( .D2(D6910_Y), .D1(D860_Y), .QN(D5462_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D5220 ( .D2(D5251_Y), .D1(D3710_Y), .QN(D5220_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D5219 ( .D2(D5252_Y), .D1(D3709_Y), .QN(D5219_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D5218 ( .D2(D5252_Y), .D1(D5249_Y), .QN(D5218_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D5217 ( .D2(D5250_Y), .D1(D1620_Y), .QN(D5217_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D5216 ( .D2(D5251_Y), .D1(D99_Y), .QN(D5216_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D5184 ( .D2(D3701_Y), .D1(D5181_Y), .QN(D5184_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D5183 ( .D2(D5251_Y), .D1(D5182_Y), .QN(D5183_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D4958 ( .D2(D4979_Y), .D1(D5052_Y), .QN(D4958_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D4957 ( .D2(D6488_Y), .D1(D6426_Y), .QN(D4957_QN),     .GN(D6461_Y));
KC_TLATHQN_X1 D4808 ( .D2(D6409_Y), .D1(D6408_Y), .QN(D4808_QN),     .GN(D536_Y));
KC_TLATHQN_X1 D4042 ( .D2(D4069_Y), .D1(D3998_Y), .QN(D4042_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4041 ( .D2(D4070_Y), .D1(D4026_Y), .QN(D4041_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4040 ( .D2(D4070_Y), .D1(D3994_Y), .QN(D4040_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4028 ( .D2(D4070_Y), .D1(D4003_Y), .QN(D4028_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4027 ( .D2(D4069_Y), .D1(D3995_Y), .QN(D4027_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4016 ( .D2(D4029_Y), .D1(D3996_Y), .QN(D4016_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4015 ( .D2(D4029_Y), .D1(D1523_Y), .QN(D4015_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4014 ( .D2(D4031_Y), .D1(D4006_Y), .QN(D4014_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4013 ( .D2(D4070_Y), .D1(D4005_Y), .QN(D4013_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4012 ( .D2(D4069_Y), .D1(D4004_Y), .QN(D4012_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4011 ( .D2(D4069_Y), .D1(D4001_Y), .QN(D4011_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4010 ( .D2(D4029_Y), .D1(D3997_Y), .QN(D4010_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4009 ( .D2(D4070_Y), .D1(D4002_Y), .QN(D4009_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D4008 ( .D2(D4029_Y), .D1(D3999_Y), .QN(D4008_QN),     .GN(D11063_Y));
KC_TLATHQN_X1 D4007 ( .D2(D4031_Y), .D1(D3989_Y), .QN(D4007_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D3873 ( .D2(D3889_Y), .D1(D3842_Y), .QN(D3873_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3872 ( .D2(D3890_Y), .D1(D3853_Y), .QN(D3872_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3871 ( .D2(D3889_Y), .D1(D3861_Y), .QN(D3871_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3870 ( .D2(D3891_Y), .D1(D3888_Y), .QN(D3870_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3868 ( .D2(D3892_Y), .D1(D3856_Y), .QN(D3868_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3867 ( .D2(D3892_Y), .D1(D3857_Y), .QN(D3867_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3866 ( .D2(D3891_Y), .D1(D3887_Y), .QN(D3866_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3865 ( .D2(D3892_Y), .D1(D3835_Y), .QN(D3865_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3864 ( .D2(D3892_Y), .D1(D3846_Y), .QN(D3864_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3798 ( .D2(D3891_Y), .D1(D3843_Y), .QN(D3798_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3797 ( .D2(D3891_Y), .D1(D3847_Y), .QN(D3797_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D3724 ( .D2(D3762_Y), .D1(D3657_Y), .QN(D3724_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D3723 ( .D2(D3762_Y), .D1(D3708_Y), .QN(D3723_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D3722 ( .D2(D3762_Y), .D1(D3761_Y), .QN(D3722_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D3671 ( .D2(D3701_Y), .D1(D3658_Y), .QN(D3671_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D3670 ( .D2(D3701_Y), .D1(D3656_Y), .QN(D3670_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D3669 ( .D2(D3701_Y), .D1(D3655_Y), .QN(D3669_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D3367 ( .D2(D3399_Y), .D1(D3335_Y), .QN(D3367_QN),     .GN(D10633_Y));
KC_TLATHQN_X1 D3271 ( .D2(D3297_Y), .D1(D3220_Y), .QN(D3271_QN),     .GN(D10633_Y));
KC_TLATHQN_X1 D3179 ( .D2(D3196_Y), .D1(D4635_Y), .QN(D3179_QN),     .GN(D10633_Y));
KC_TLATHQN_X1 D3178 ( .D2(D3201_Y), .D1(D367_Y), .QN(D3178_QN),     .GN(D10633_Y));
KC_TLATHQN_X1 D3177 ( .D2(D3201_Y), .D1(D3153_Y), .QN(D3177_QN),     .GN(D10633_Y));
KC_TLATHQN_X1 D3176 ( .D2(D3201_Y), .D1(D3239_Y), .QN(D3176_QN),     .GN(D10633_Y));
KC_TLATHQN_X1 D2791 ( .D2(D2811_Y), .D1(D2753_Y), .QN(D2791_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D2790 ( .D2(D2811_Y), .D1(D2776_Y), .QN(D2790_QN),     .GN(D1947_Y));
KC_TLATHQN_X1 D2513 ( .D2(D16336_Y), .D1(D16295_Y), .QN(D2513_QN),     .GN(D15867_Y));
KC_TLATHQN_X1 D2287 ( .D2(D11932_Y), .D1(D11364_Y), .QN(D2287_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D2286 ( .D2(D11996_Y), .D1(D11415_Y), .QN(D2286_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D2154 ( .D2(D10898_Y), .D1(D10850_Y), .QN(D2154_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D2153 ( .D2(D11088_Y), .D1(D11052_Y), .QN(D2153_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D2150 ( .D2(D10898_Y), .D1(D10868_Y), .QN(D2150_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D2071 ( .D2(D11113_Y), .D1(D1285_Y), .QN(D2071_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D1631 ( .D2(D1673_Y), .D1(D5046_Y), .QN(D1631_QN),     .GN(D536_Y));
KC_TLATHQN_X1 D1487 ( .D2(D4069_Y), .D1(D4000_Y), .QN(D1487_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D1486 ( .D2(D3889_Y), .D1(D3852_Y), .QN(D1486_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D1485 ( .D2(D3889_Y), .D1(D3854_Y), .QN(D1485_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D1484 ( .D2(D3891_Y), .D1(D3832_Y), .QN(D1484_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D1483 ( .D2(D3892_Y), .D1(D3858_Y), .QN(D1483_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D1402 ( .D2(D16592_Y), .D1(D16574_Y), .QN(D1402_QN),     .GN(D15867_Y));
KC_TLATHQN_X1 D1347 ( .D2(D12128_Y), .D1(D11555_Y), .QN(D1347_QN),     .GN(D12104_Y));
KC_TLATHQN_X1 D1287 ( .D2(D11590_Y), .D1(D11557_Y), .QN(D1287_QN),     .GN(D12104_Y));
KC_TLATHQN_X1 D1198 ( .D2(D11088_Y), .D1(D1330_Y), .QN(D1198_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D1197 ( .D2(D11089_Y), .D1(D11062_Y), .QN(D1197_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D1196 ( .D2(D4031_Y), .D1(D3988_Y), .QN(D1196_QN),     .GN(D5557_Y));
KC_TLATHQN_X1 D1120 ( .D2(D11996_Y), .D1(D11903_Y), .QN(D1120_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D1119 ( .D2(D11933_Y), .D1(D11381_Y), .QN(D1119_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D1118 ( .D2(D11996_Y), .D1(D11436_Y), .QN(D1118_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D1011 ( .D2(D11349_Y), .D1(D11303_Y), .QN(D1011_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D1010 ( .D2(D11933_Y), .D1(D11374_Y), .QN(D1010_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D1009 ( .D2(D6910_Y), .D1(D862_Y), .QN(D1009_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D901 ( .D2(D10897_Y), .D1(D10865_Y), .QN(D901_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D900 ( .D2(D10898_Y), .D1(D10867_Y), .QN(D900_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D899 ( .D2(D10896_Y), .D1(D2238_Y), .QN(D899_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D898 ( .D2(D10895_Y), .D1(D10853_Y), .QN(D898_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D897 ( .D2(D10897_Y), .D1(D10851_Y), .QN(D897_QN),     .GN(D10871_Y));
KC_TLATHQN_X1 D894 ( .D2(D3890_Y), .D1(D3844_Y), .QN(D894_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D893 ( .D2(D6833_Y), .D1(D6774_Y), .QN(D893_QN),     .GN(D6798_Y));
KC_TLATHQN_X1 D892 ( .D2(D1675_Y), .D1(D861_Y), .QN(D892_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D891 ( .D2(D1675_Y), .D1(D3855_Y), .QN(D891_QN),     .GN(D3860_Y));
KC_TLATHQN_X1 D782 ( .D2(D12867_Y), .D1(D12835_Y), .QN(D782_QN),     .GN(D12859_Y));
KC_TLATHQN_X1 D780 ( .D2(D12867_Y), .D1(D12833_Y), .QN(D780_QN),     .GN(D830_Y));
KC_TLATHQN_X1 D775 ( .D2(D8263_Y), .D1(D9430_Y), .QN(D775_QN),     .GN(D534_Y));
KC_TLATHQN_X1 D718 ( .D2(D11279_Y), .D1(D631_Y), .QN(D718_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D661 ( .D2(D11184_Y), .D1(D11710_Y), .QN(D661_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D660 ( .D2(D11279_Y), .D1(D11160_Y), .QN(D660_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D657 ( .D2(D5251_Y), .D1(D3721_Y), .QN(D657_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D656 ( .D2(D5251_Y), .D1(D3715_Y), .QN(D656_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D655 ( .D2(D5251_Y), .D1(D3720_Y), .QN(D655_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D588 ( .D2(D11135_Y), .D1(D11149_Y), .QN(D588_QN),     .GN(D11172_Y));
KC_TLATHQN_X1 D587 ( .D2(D3701_Y), .D1(D3667_Y), .QN(D587_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D586 ( .D2(D3701_Y), .D1(D575_Y), .QN(D586_QN),     .GN(D1663_Y));
KC_TLATHQN_X1 D507 ( .D2(D16768_Y), .D1(D14805_Y), .QN(D507_QN),     .GN(D13249_Y));
KC_TLATHQN_X1 D506 ( .D2(D13867_Y), .D1(D13889_Y), .QN(D506_QN),     .GN(D13910_Y));
KC_TLATHQN_X1 D503 ( .D2(D7993_Y), .D1(D7913_Y), .QN(D503_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D478 ( .D2(D6497_Y), .D1(D6496_Y), .QN(D478_QN),     .GN(D6484_Y));
KC_TLATHQN_X1 D443 ( .D2(D1972_Y), .D1(D7570_Y), .QN(D443_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D416 ( .D2(D7754_Y), .D1(D9207_Y), .QN(D416_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D415 ( .D2(D7754_Y), .D1(D375_Y), .QN(D415_QN),     .GN(D9224_Y));
KC_TLATHQN_X1 D380 ( .D2(D4742_Y), .D1(D3156_Y), .QN(D380_QN),     .GN(D10633_Y));
KC_TLATHQN_X1 D296 ( .D2(D270_Y), .D1(D7370_Y), .QN(D296_QN),     .GN(D7520_Y));
KC_TLATHQN_X1 D261 ( .D2(D2105_Y), .D1(D7400_Y), .QN(D261_QN),     .GN(D5812_Y));
KC_TLATHQN_X1 D226 ( .D2(D7161_Y), .D1(D7163_Y), .QN(D226_QN),     .GN(D7520_Y));
KC_TLATHQN_X1 D191 ( .D2(D7161_Y), .D1(D7126_Y), .QN(D191_QN),     .GN(D534_Y));
KC_TLATHQN_X1 D112 ( .D2(D11933_Y), .D1(D1005_Y), .QN(D112_QN),     .GN(D767_Y));
KC_TLATHQN_X1 D111 ( .D2(D11089_Y), .D1(D1286_Y), .QN(D111_QN),     .GN(D9699_Y));
KC_TLATHQN_X1 D108 ( .D2(D2811_Y), .D1(D2777_Y), .QN(D108_QN),     .GN(D7520_Y));
KC_XNOR2_X1 D16222 ( .Y(D16222_Y), .A(D16211_Y), .B(D16215_Y));
KC_XNOR2_X1 D16165 ( .Y(D16165_Y), .A(D16116_Y), .B(D16073_Y));
KC_XNOR2_X1 D16154 ( .Y(D16154_Y), .A(D16136_Y), .B(D16167_Y));
KC_XNOR2_X1 D14679 ( .Y(D14679_Y), .A(D16172_Y), .B(D14671_Y));
KC_XNOR2_X1 D14514 ( .Y(D14514_Y), .A(D14526_Y), .B(D7822_Y));
KC_XNOR2_X1 D14513 ( .Y(D14513_Y), .A(D14525_Y), .B(D7822_Y));
KC_XNOR2_X1 D349 ( .Y(D349_Y), .A(D13861_Y), .B(D2504_Y));
KC_XNOR2_X1 D13855 ( .Y(D13855_Y), .A(D13863_Y), .B(D2507_Y));
KC_XNOR2_X1 D13702 ( .Y(D13702_Y), .A(D13015_Y), .B(D16005_Y));
KC_XNOR2_X1 D12173 ( .Y(D12173_Y), .A(D2106_Y), .B(D490_Y));
KC_XNOR2_X1 D11654 ( .Y(D11654_Y), .A(D10181_Y), .B(D12197_Y));
KC_XNOR2_X1 D11653 ( .Y(D11653_Y), .A(D11654_Y), .B(D11645_Y));
KC_XNOR2_X1 D11101 ( .Y(D11101_Y), .A(D11073_Q), .B(D11098_Y));
KC_XNOR2_X1 D9566 ( .Y(D9566_Y), .A(D9593_Y), .B(D835_Q));
KC_XNOR2_X1 D9564 ( .Y(D9564_Y), .A(D9567_Y), .B(D857_Q));
KC_XNOR2_X1 D9264 ( .Y(D9264_Y), .A(D9263_Y), .B(D6301_Y));
KC_XNOR2_X1 D9210 ( .Y(D9210_Y), .A(D7686_Y), .B(D9230_Co));
KC_XNOR2_X1 D9146 ( .Y(D9146_Y), .A(D9121_Y), .B(D9136_Y));
KC_XNOR2_X1 D8812 ( .Y(D8812_Y), .A(D8799_Y), .B(D8804_Y));
KC_XNOR2_X1 D8704 ( .Y(D8704_Y), .A(D8706_Y), .B(D7125_Y));
KC_XNOR2_X1 D8702 ( .Y(D8702_Y), .A(D8726_Y), .B(D187_Y));
KC_XNOR2_X1 D8699 ( .Y(D8699_Y), .A(D8705_Y), .B(D8817_Y));
KC_XNOR2_X1 D8326 ( .Y(D8326_Y), .A(D8341_Q), .B(D8324_Y));
KC_XNOR2_X1 D8234 ( .Y(D8234_Y), .A(D8190_Y), .B(D8256_Y));
KC_XNOR2_X1 D7727 ( .Y(D7727_Y), .A(D420_Q), .B(D7690_Y));
KC_XNOR2_X1 D7723 ( .Y(D7723_Y), .A(D6335_Y), .B(D7682_Y));
KC_XNOR2_X1 D7656 ( .Y(D7656_Y), .A(D7626_Y), .B(D7659_Q));
KC_XNOR2_X1 D7654 ( .Y(D7654_Y), .A(D373_Y), .B(D7577_S));
KC_XNOR2_X1 D7652 ( .Y(D7652_Y), .A(D7630_Y), .B(D7651_Y));
KC_XNOR2_X1 D7651 ( .Y(D7651_Y), .A(D7658_Y), .B(D15451_Y));
KC_XNOR2_X1 D7584 ( .Y(D7584_Y), .A(D7554_Y), .B(D16156_Y));
KC_XNOR2_X1 D7582 ( .Y(D7582_Y), .A(D9264_Y), .B(D7574_Y));
KC_XNOR2_X1 D7581 ( .Y(D7581_Y), .A(D7548_Y), .B(D7543_Y));
KC_XNOR2_X1 D7521 ( .Y(D7521_Y), .A(D7556_Y), .B(D7513_Y));
KC_XNOR2_X1 D7141 ( .Y(D7141_Y), .A(D7145_Q), .B(D7131_Y));
KC_XNOR2_X1 D7140 ( .Y(D7140_Y), .A(D4105_Y), .B(D7147_Q));
KC_XNOR2_X1 D7137 ( .Y(D7137_Y), .A(D8687_Y), .B(D7150_Q));
KC_XNOR2_X1 D6469 ( .Y(D6469_Y), .A(D6450_Y), .B(D6452_Y));
KC_XNOR2_X1 D6338 ( .Y(D6338_Y), .A(D6322_Y), .B(D6331_Y));
KC_XNOR2_X1 D6337 ( .Y(D6337_Y), .A(D6297_Y), .B(D6300_Y));
KC_XNOR2_X1 D6261 ( .Y(D6261_Y), .A(D6304_Y), .B(D6243_Y));
KC_XNOR2_X1 D6257 ( .Y(D6257_Y), .A(D6277_Y), .B(D6225_Y));
KC_XNOR2_X1 D6174 ( .Y(D6174_Y), .A(D6352_Y), .B(D6141_Y));
KC_XNOR2_X1 D6171 ( .Y(D6171_Y), .A(D6135_Y), .B(D6133_Y));
KC_XNOR2_X1 D6170 ( .Y(D6170_Y), .A(D6136_Y), .B(D6284_Q));
KC_XNOR2_X1 D6169 ( .Y(D6169_Y), .A(D1704_Y), .B(D6163_Y));
KC_XNOR2_X1 D6115 ( .Y(D6115_Y), .A(D7531_Y), .B(D6100_Y));
KC_XNOR2_X1 D5393 ( .Y(D5393_Y), .A(D5404_Y), .B(D5343_Y));
KC_XNOR2_X1 D5076 ( .Y(D5076_Y), .A(D7954_Y), .B(D5051_Y));
KC_XNOR2_X1 D4806 ( .Y(D4806_Y), .A(D9352_Y), .B(D4681_Y));
KC_XNOR2_X1 D4630 ( .Y(D4630_Y), .A(D8152_Y), .B(D6137_Y));
KC_XNOR2_X1 D4628 ( .Y(D4628_Y), .A(D3175_Y), .B(D6210_Y));
KC_XNOR2_X1 D4551 ( .Y(D4551_Y), .A(D3051_Y), .B(D6144_Y));
KC_XNOR2_X1 D4470 ( .Y(D4470_Y), .A(D4460_Y), .B(D4491_Q));
KC_XNOR2_X1 D4466 ( .Y(D4466_Y), .A(D4481_Y), .B(D4411_Y));
KC_XNOR2_X1 D4231 ( .Y(D4231_Y), .A(D5693_Q), .B(D20_Y));
KC_XNOR2_X1 D4117 ( .Y(D4117_Y), .A(D4123_Y), .B(D4101_Y));
KC_XNOR2_X1 D3869 ( .Y(D3869_Y), .A(D3833_Y), .B(D3859_Y));
KC_XNOR2_X1 D3796 ( .Y(D3796_Y), .A(D3809_Q), .B(D3869_Y));
KC_XNOR2_X1 D3479 ( .Y(D3479_Y), .A(D3483_Q), .B(D3588_Y));
KC_XNOR2_X1 D3477 ( .Y(D3477_Y), .A(D16006_Y), .B(D3482_Q));
KC_XNOR2_X1 D3369 ( .Y(D3369_Y), .A(D3345_Y), .B(D3386_Q));
KC_XNOR2_X1 D3368 ( .Y(D3368_Y), .A(D4839_Y), .B(D3382_Q));
KC_XNOR2_X1 D3365 ( .Y(D3365_Y), .A(D1517_Q), .B(D3366_Y));
KC_XNOR2_X1 D3274 ( .Y(D3274_Y), .A(D4717_Y), .B(D3267_Y));
KC_XNOR2_X1 D3273 ( .Y(D3273_Y), .A(D3280_Q), .B(D4621_Y));
KC_XNOR2_X1 D3270 ( .Y(D3270_Y), .A(D7647_Q), .B(D3272_Y));
KC_XNOR2_X1 D3175 ( .Y(D3175_Y), .A(D3191_Y), .B(D3166_Y));
KC_XNOR2_X1 D3070 ( .Y(D3070_Y), .A(D2996_Y), .B(D2954_Y));
KC_XNOR2_X1 D3069 ( .Y(D3069_Y), .A(D3076_Y), .B(D1536_Q));
KC_XNOR2_X1 D3068 ( .Y(D3068_Y), .A(D3072_Y), .B(D3073_Y));
KC_XNOR2_X1 D2991 ( .Y(D2991_Y), .A(D2990_Y), .B(D2989_Y));
KC_XNOR2_X1 D2989 ( .Y(D2989_Y), .A(D2953_Y), .B(D2910_Y));
KC_XNOR2_X1 D2877 ( .Y(D2877_Y), .A(D2856_Y), .B(D2830_Y));
KC_XNOR2_X1 D2876 ( .Y(D2876_Y), .A(D2884_Q), .B(D2887_Q));
KC_XNOR2_X1 D2675 ( .Y(D2675_Y), .A(D16120_Y), .B(D2673_Y));
KC_XNOR2_X1 D2674 ( .Y(D2674_Y), .A(D84_Y), .B(D2671_Y));
KC_XNOR2_X1 D2637 ( .Y(D2637_Y), .A(D2618_Y), .B(D2667_Y));
KC_XNOR2_X1 D2155 ( .Y(D2155_Y), .A(D958_Y), .B(D10293_Q));
KC_XNOR2_X1 D2072 ( .Y(D2072_Y), .A(D9633_Y), .B(D2107_Y));
KC_XNOR2_X1 D1925 ( .Y(D1925_Y), .A(D6200_Y), .B(D7553_Y));
KC_XNOR2_X1 D1923 ( .Y(D1923_Y), .A(D7660_Y), .B(D7565_Y));
KC_XNOR2_X1 D1771 ( .Y(D1771_Y), .A(D6143_Y), .B(D6119_Y));
KC_XNOR2_X1 D1629 ( .Y(D1629_Y), .A(D194_Q), .B(D1630_Y));
KC_XNOR2_X1 D896 ( .Y(D896_Y), .A(D933_Q), .B(D8315_Y));
KC_XNOR2_X1 D776 ( .Y(D776_Y), .A(D15600_Y), .B(D851_Q));
KC_XNOR2_X1 D322 ( .Y(D322_Y), .A(D6143_Y), .B(D6102_Y));
KC_XNOR2_X1 D262 ( .Y(D262_Y), .A(D6066_Y), .B(D264_Q));
KC_XNOR2_X1 D189 ( .Y(D189_Y), .A(D193_Q), .B(D8795_Y));
KC_XNOR2_X1 D109 ( .Y(D109_Y), .A(D13174_Y), .B(D2459_Y));
KC_XNOR2_X1 D107 ( .Y(D107_Y), .A(D1419_Y), .B(D6306_Y));
KC_BUF_X3 D16381 ( .Y(D16381_Y), .A(D15608_Y));
KC_BUF_X3 D16351 ( .Y(D16351_Y), .A(D15649_Y));
KC_BUF_X3 D16309 ( .Y(D16309_Y), .A(D15548_Y));
KC_BUF_X3 D16284 ( .Y(D16284_Y), .A(D16297_Y));
KC_BUF_X3 D16283 ( .Y(D16283_Y), .A(D2660_Y));
KC_BUF_X3 D16282 ( .Y(D16282_Y), .A(D16280_Y));
KC_BUF_X3 D16280 ( .Y(D16280_Y), .A(D16258_Y));
KC_BUF_X3 D16278 ( .Y(D16278_Y), .A(D15595_Y));
KC_BUF_X3 D16140 ( .Y(D16140_Y), .A(D16119_Y));
KC_BUF_X3 D16017 ( .Y(D16017_Y), .A(D9951_Y));
KC_BUF_X3 D15987 ( .Y(D15987_Y), .A(D15163_Y));
KC_BUF_X3 D15944 ( .Y(D15944_Y), .A(D15674_Y));
KC_BUF_X3 D15864 ( .Y(D15864_Y), .A(D15830_Y));
KC_BUF_X3 D15863 ( .Y(D15863_Y), .A(D15828_Y));
KC_BUF_X3 D15787 ( .Y(D15787_Y), .A(D986_Y));
KC_BUF_X3 D15786 ( .Y(D15786_Y), .A(D15730_Y));
KC_BUF_X3 D15664 ( .Y(D15664_Y), .A(D15701_Y));
KC_BUF_X3 D15563 ( .Y(D15563_Y), .A(D16461_Y));
KC_BUF_X3 D15562 ( .Y(D15562_Y), .A(D16461_Y));
KC_BUF_X3 D15443 ( .Y(D15443_Y), .A(D14517_Y));
KC_BUF_X3 D15442 ( .Y(D15442_Y), .A(D14523_Y));
KC_BUF_X3 D15441 ( .Y(D15441_Y), .A(D15262_Y));
KC_BUF_X3 D15250 ( .Y(D15250_Y), .A(D15290_Y));
KC_BUF_X3 D15249 ( .Y(D15249_Y), .A(D10127_Y));
KC_BUF_X3 D15210 ( .Y(D15210_Y), .A(D15196_Y));
KC_BUF_X3 D15209 ( .Y(D15209_Y), .A(D15187_Y));
KC_BUF_X3 D15208 ( .Y(D15208_Y), .A(D15160_Y));
KC_BUF_X3 D15128 ( .Y(D15128_Y), .A(D15609_Y));
KC_BUF_X3 D15073 ( .Y(D15073_Y), .A(D15045_Y));
KC_BUF_X3 D14678 ( .Y(D14678_Y), .A(D15418_Y));
KC_BUF_X3 D14585 ( .Y(D14585_Y), .A(D608_Q));
KC_BUF_X3 D14584 ( .Y(D14584_Y), .A(D14520_Q));
KC_BUF_X3 D14512 ( .Y(D14512_Y), .A(D10122_Y));
KC_BUF_X3 D14511 ( .Y(D14511_Y), .A(D10141_Y));
KC_BUF_X3 D14510 ( .Y(D14510_Y), .A(D10151_Y));
KC_BUF_X3 D14509 ( .Y(D14509_Y), .A(D10117_Y));
KC_BUF_X3 D14508 ( .Y(D14508_Y), .A(D10124_Y));
KC_BUF_X3 D14294 ( .Y(D14294_Y), .A(D14937_Y));
KC_BUF_X3 D13981 ( .Y(D13981_Y), .A(D13942_Y));
KC_BUF_X3 D13980 ( .Y(D13980_Y), .A(D639_Y));
KC_BUF_X3 D13979 ( .Y(D13979_Y), .A(D13978_Y));
KC_BUF_X3 D13978 ( .Y(D13978_Y), .A(D13951_Y));
KC_BUF_X3 D13977 ( .Y(D13977_Y), .A(D13275_Q));
KC_BUF_X3 D13976 ( .Y(D13976_Y), .A(D694_Q));
KC_BUF_X3 D13975 ( .Y(D13975_Y), .A(D13994_Q));
KC_BUF_X3 D13974 ( .Y(D13974_Y), .A(D12683_Q));
KC_BUF_X3 D13906 ( .Y(D13906_Y), .A(D12680_Q));
KC_BUF_X3 D13796 ( .Y(D13796_Y), .A(D14457_Y));
KC_BUF_X3 D13795 ( .Y(D13795_Y), .A(D14449_Y));
KC_BUF_X3 D13752 ( .Y(D13752_Y), .A(D14477_Y));
KC_BUF_X3 D13751 ( .Y(D13751_Y), .A(D13720_Y));
KC_BUF_X3 D13750 ( .Y(D13750_Y), .A(D13721_Y));
KC_BUF_X3 D13701 ( .Y(D13701_Y), .A(D1090_Y));
KC_BUF_X3 D13260 ( .Y(D13260_Y), .A(D13943_Y));
KC_BUF_X3 D13259 ( .Y(D13259_Y), .A(D2390_Q));
KC_BUF_X3 D13258 ( .Y(D13258_Y), .A(D13895_Y));
KC_BUF_X3 D13257 ( .Y(D13257_Y), .A(D13236_Y));
KC_BUF_X3 D13192 ( .Y(D13192_Y), .A(D12280_Y));
KC_BUF_X3 D13191 ( .Y(D13191_Y), .A(D13202_Q));
KC_BUF_X3 D13190 ( .Y(D13190_Y), .A(D13990_Q));
KC_BUF_X3 D13164 ( .Y(D13164_Y), .A(D2464_Y));
KC_BUF_X3 D13163 ( .Y(D13163_Y), .A(D13272_Q));
KC_BUF_X3 D13162 ( .Y(D13162_Y), .A(D13271_Q));
KC_BUF_X3 D13161 ( .Y(D13161_Y), .A(D13199_Q));
KC_BUF_X3 D13160 ( .Y(D13160_Y), .A(D13991_Q));
KC_BUF_X3 D13159 ( .Y(D13159_Y), .A(D13197_Q));
KC_BUF_X3 D13158 ( .Y(D13158_Y), .A(D13998_Q));
KC_BUF_X3 D13157 ( .Y(D13157_Y), .A(D13208_Q));
KC_BUF_X3 D13030 ( .Y(D13030_Y), .A(D13712_Y));
KC_BUF_X3 D12840 ( .Y(D12840_Y), .A(D12796_Y));
KC_BUF_X3 D12676 ( .Y(D12676_Y), .A(D697_Q));
KC_BUF_X3 D12675 ( .Y(D12675_Y), .A(D12689_Q));
KC_BUF_X3 D12674 ( .Y(D12674_Y), .A(D13203_Q));
KC_BUF_X3 D12656 ( .Y(D12656_Y), .A(D13210_Q));
KC_BUF_X3 D12632 ( .Y(D12632_Y), .A(D13209_Q));
KC_BUF_X3 D12631 ( .Y(D12631_Y), .A(D13200_Q));
KC_BUF_X3 D12630 ( .Y(D12630_Y), .A(D12685_Q));
KC_BUF_X3 D12629 ( .Y(D12629_Y), .A(D13279_Q));
KC_BUF_X3 D12628 ( .Y(D12628_Y), .A(D12684_Q));
KC_BUF_X3 D12627 ( .Y(D12627_Y), .A(D12686_Q));
KC_BUF_X3 D12626 ( .Y(D12626_Y), .A(D692_Q));
KC_BUF_X3 D12227 ( .Y(D12227_Y), .A(D12687_Q));
KC_BUF_X3 D12226 ( .Y(D12226_Y), .A(D12682_Q));
KC_BUF_X3 D12225 ( .Y(D12225_Y), .A(D12688_Q));
KC_BUF_X3 D12224 ( .Y(D12224_Y), .A(D12681_Q));
KC_BUF_X3 D12223 ( .Y(D12223_Y), .A(D12156_Y));
KC_BUF_X3 D12222 ( .Y(D12222_Y), .A(D12223_Y));
KC_BUF_X3 D12170 ( .Y(D12170_Y), .A(D12158_Y));
KC_BUF_X3 D12169 ( .Y(D12169_Y), .A(D12152_Y));
KC_BUF_X3 D12168 ( .Y(D12168_Y), .A(D2338_Y));
KC_BUF_X3 D12167 ( .Y(D12167_Y), .A(D12222_Y));
KC_BUF_X3 D12166 ( .Y(D12166_Y), .A(D2339_Y));
KC_BUF_X3 D12165 ( .Y(D12165_Y), .A(D12169_Y));
KC_BUF_X3 D12164 ( .Y(D12164_Y), .A(D12163_Y));
KC_BUF_X3 D12163 ( .Y(D12163_Y), .A(D12151_Y));
KC_BUF_X3 D12162 ( .Y(D12162_Y), .A(D12160_Y));
KC_BUF_X3 D12161 ( .Y(D12161_Y), .A(D12155_Y));
KC_BUF_X3 D12160 ( .Y(D12160_Y), .A(D12159_Y));
KC_BUF_X3 D12159 ( .Y(D12159_Y), .A(D12171_Y));
KC_BUF_X3 D12158 ( .Y(D12158_Y), .A(D12153_Y));
KC_BUF_X3 D12157 ( .Y(D12157_Y), .A(D12167_Y));
KC_BUF_X3 D12156 ( .Y(D12156_Y), .A(D2340_Y));
KC_BUF_X3 D12155 ( .Y(D12155_Y), .A(D12170_Y));
KC_BUF_X3 D12154 ( .Y(D12154_Y), .A(D12165_Y));
KC_BUF_X3 D12153 ( .Y(D12153_Y), .A(D12154_Y));
KC_BUF_X3 D12152 ( .Y(D12152_Y), .A(D12164_Y));
KC_BUF_X3 D12151 ( .Y(D12151_Y), .A(D12162_Y));
KC_BUF_X3 D12150 ( .Y(D12150_Y), .A(D12161_Y));
KC_BUF_X3 D12149 ( .Y(D12149_Y), .A(D12147_Y));
KC_BUF_X3 D12148 ( .Y(D12148_Y), .A(D12182_Y));
KC_BUF_X3 D12147 ( .Y(D12147_Y), .A(D2863_Y));
KC_BUF_X3 D12146 ( .Y(D12146_Y), .A(D12145_Y));
KC_BUF_X3 D12145 ( .Y(D12145_Y), .A(D12142_Y));
KC_BUF_X3 D12144 ( .Y(D12144_Y), .A(D12149_Y));
KC_BUF_X3 D12142 ( .Y(D12142_Y), .A(D12148_Y));
KC_BUF_X3 D12141 ( .Y(D12141_Y), .A(D10121_Y));
KC_BUF_X3 D11970 ( .Y(D11970_Y), .A(D11958_Y));
KC_BUF_X3 D11969 ( .Y(D11969_Y), .A(D9555_Y));
KC_BUF_X3 D11626 ( .Y(D11626_Y), .A(D504_Y));
KC_BUF_X3 D11536 ( .Y(D11536_Y), .A(D621_Y));
KC_BUF_X3 D11535 ( .Y(D11535_Y), .A(D621_Y));
KC_BUF_X3 D11465 ( .Y(D11465_Y), .A(D621_Y));
KC_BUF_X3 D11386 ( .Y(D11386_Y), .A(D2244_Y));
KC_BUF_X3 D11322 ( .Y(D11322_Y), .A(D169_Y));
KC_BUF_X3 D11259 ( .Y(D11259_Y), .A(D8060_Y));
KC_BUF_X3 D11258 ( .Y(D11258_Y), .A(D621_Y));
KC_BUF_X3 D11257 ( .Y(D11257_Y), .A(D621_Y));
KC_BUF_X3 D11256 ( .Y(D11256_Y), .A(D621_Y));
KC_BUF_X3 D11255 ( .Y(D11255_Y), .A(D8177_Y));
KC_BUF_X3 D11024 ( .Y(D11024_Y), .A(D12070_Y));
KC_BUF_X3 D10990 ( .Y(D10990_Y), .A(D9555_Y));
KC_BUF_X3 D10788 ( .Y(D10788_Y), .A(D8013_Y));
KC_BUF_X3 D10787 ( .Y(D10787_Y), .A(D7990_Y));
KC_BUF_X3 D10344 ( .Y(D10344_Y), .A(D10335_Y));
KC_BUF_X3 D10343 ( .Y(D10343_Y), .A(D10320_Y));
KC_BUF_X3 D10342 ( .Y(D10342_Y), .A(D10320_Y));
KC_BUF_X3 D10341 ( .Y(D10341_Y), .A(D10334_Y));
KC_BUF_X3 D10340 ( .Y(D10340_Y), .A(D10337_Y));
KC_BUF_X3 D10339 ( .Y(D10339_Y), .A(D10332_Y));
KC_BUF_X3 D10338 ( .Y(D10338_Y), .A(D10342_Y));
KC_BUF_X3 D10337 ( .Y(D10337_Y), .A(D10343_Y));
KC_BUF_X3 D10336 ( .Y(D10336_Y), .A(D10333_Y));
KC_BUF_X3 D10335 ( .Y(D10335_Y), .A(D10340_Y));
KC_BUF_X3 D10334 ( .Y(D10334_Y), .A(D10336_Y));
KC_BUF_X3 D10333 ( .Y(D10333_Y), .A(D10338_Y));
KC_BUF_X3 D10332 ( .Y(D10332_Y), .A(D10320_Y));
KC_BUF_X3 D10331 ( .Y(D10331_Y), .A(D10320_Y));
KC_BUF_X3 D10330 ( .Y(D10330_Y), .A(D2148_Y));
KC_BUF_X3 D10329 ( .Y(D10329_Y), .A(D10339_Y));
KC_BUF_X3 D10328 ( .Y(D10328_Y), .A(D836_Q));
KC_BUF_X3 D10327 ( .Y(D10327_Y), .A(D10344_Y));
KC_BUF_X3 D10326 ( .Y(D10326_Y), .A(D10331_Y));
KC_BUF_X3 D10325 ( .Y(D10325_Y), .A(D10324_Y));
KC_BUF_X3 D10324 ( .Y(D10324_Y), .A(D10323_Y));
KC_BUF_X3 D10323 ( .Y(D10323_Y), .A(D10326_Y));
KC_BUF_X3 D10315 ( .Y(D10315_Y), .A(D2175_Q));
KC_BUF_X3 D10285 ( .Y(D10285_Y), .A(D10271_Y));
KC_BUF_X3 D10284 ( .Y(D10284_Y), .A(D10283_Y));
KC_BUF_X3 D10283 ( .Y(D10283_Y), .A(D10277_Y));
KC_BUF_X3 D10282 ( .Y(D10282_Y), .A(D10278_Y));
KC_BUF_X3 D10281 ( .Y(D10281_Y), .A(D10280_Y));
KC_BUF_X3 D10280 ( .Y(D10280_Y), .A(D10356_Y));
KC_BUF_X3 D10279 ( .Y(D10279_Y), .A(D10356_Y));
KC_BUF_X3 D10278 ( .Y(D10278_Y), .A(D10284_Y));
KC_BUF_X3 D10277 ( .Y(D10277_Y), .A(D10279_Y));
KC_BUF_X3 D10276 ( .Y(D10276_Y), .A(D10272_Y));
KC_BUF_X3 D10275 ( .Y(D10275_Y), .A(D10267_Y));
KC_BUF_X3 D10274 ( .Y(D10274_Y), .A(D10281_Y));
KC_BUF_X3 D10273 ( .Y(D10273_Y), .A(D10268_Y));
KC_BUF_X3 D10272 ( .Y(D10272_Y), .A(D10274_Y));
KC_BUF_X3 D10271 ( .Y(D10271_Y), .A(D10276_Y));
KC_BUF_X3 D10270 ( .Y(D10270_Y), .A(D10273_Y));
KC_BUF_X3 D10269 ( .Y(D10269_Y), .A(D10315_Y));
KC_BUF_X3 D10268 ( .Y(D10268_Y), .A(D10275_Y));
KC_BUF_X3 D10267 ( .Y(D10267_Y), .A(D10307_Q));
KC_BUF_X3 D10235 ( .Y(D10235_Y), .A(D10217_Q));
KC_BUF_X3 D10210 ( .Y(D10210_Y), .A(D9566_Y));
KC_BUF_X3 D9979 ( .Y(D9979_Y), .A(D9978_Y));
KC_BUF_X3 D9978 ( .Y(D9978_Y), .A(D8803_Y));
KC_BUF_X3 D9977 ( .Y(D9977_Y), .A(D10095_Y));
KC_BUF_X3 D9935 ( .Y(D9935_Y), .A(D9934_Y));
KC_BUF_X3 D9934 ( .Y(D9934_Y), .A(D9934_A));
KC_BUF_X3 D9933 ( .Y(D9933_Y), .A(D183_Y));
KC_BUF_X3 D9781 ( .Y(D9781_Y), .A(D621_Y));
KC_BUF_X3 D9636 ( .Y(D9636_Y), .A(D2067_Y));
KC_BUF_X3 D9605 ( .Y(D9605_Y), .A(D9604_Y));
KC_BUF_X3 D9604 ( .Y(D9604_Y), .A(D10362_Q));
KC_BUF_X3 D9603 ( .Y(D9603_Y), .A(D9602_Y));
KC_BUF_X3 D9602 ( .Y(D9602_Y), .A(D10362_Q));
KC_BUF_X3 D9601 ( .Y(D9601_Y), .A(D9600_Y));
KC_BUF_X3 D9600 ( .Y(D9600_Y), .A(D9603_Y));
KC_BUF_X3 D9563 ( .Y(D9563_Y), .A(D67_Y));
KC_BUF_X3 D9562 ( .Y(D9562_Y), .A(D8229_Y));
KC_BUF_X3 D9561 ( .Y(D9561_Y), .A(D9592_Y));
KC_BUF_X3 D9452 ( .Y(D9452_Y), .A(D10231_Q));
KC_BUF_X3 D9451 ( .Y(D9451_Y), .A(D9452_Y));
KC_BUF_X3 D9450 ( .Y(D9450_Y), .A(D9451_Y));
KC_BUF_X3 D9449 ( .Y(D9449_Y), .A(D10235_Y));
KC_BUF_X3 D9352 ( .Y(D9352_Y), .A(D16762_Y));
KC_BUF_X3 D9351 ( .Y(D9351_Y), .A(D9350_Y));
KC_BUF_X3 D9349 ( .Y(D9349_Y), .A(D9276_Q));
KC_BUF_X3 D9262 ( .Y(D9262_Y), .A(D9099_Y));
KC_BUF_X3 D9261 ( .Y(D9261_Y), .A(D7613_Y));
KC_BUF_X3 D9138 ( .Y(D9138_Y), .A(D2069_Y));
KC_BUF_X3 D9137 ( .Y(D9137_Y), .A(D9135_Y));
KC_BUF_X3 D9136 ( .Y(D9136_Y), .A(D7660_Y));
KC_BUF_X3 D9135 ( .Y(D9135_Y), .A(D41_Y));
KC_BUF_X3 D9134 ( .Y(D9134_Y), .A(D9133_Y));
KC_BUF_X3 D9133 ( .Y(D9133_Y), .A(D57_Y));
KC_BUF_X3 D9089 ( .Y(D9089_Y), .A(D40_Q));
KC_BUF_X3 D9088 ( .Y(D9088_Y), .A(D6248_Q));
KC_BUF_X3 D8806 ( .Y(D8806_Y), .A(D9298_Y));
KC_BUF_X3 D8805 ( .Y(D8805_Y), .A(D7257_Y));
KC_BUF_X3 D8803 ( .Y(D8803_Y), .A(D2147_Y));
KC_BUF_X3 D8697 ( .Y(D8697_Y), .A(D8770_Y));
KC_BUF_X3 D8534 ( .Y(D8534_Y), .A(D7974_Y));
KC_BUF_X3 D8533 ( .Y(D8533_Y), .A(D8013_Y));
KC_BUF_X3 D8532 ( .Y(D8532_Y), .A(D621_Y));
KC_BUF_X3 D8456 ( .Y(D8456_Y), .A(D3916_Y));
KC_BUF_X3 D8455 ( .Y(D8455_Y), .A(D8013_Y));
KC_BUF_X3 D8323 ( .Y(D8323_Y), .A(D7895_Y));
KC_BUF_X3 D8322 ( .Y(D8322_Y), .A(D8318_Y));
KC_BUF_X3 D8321 ( .Y(D8321_Y), .A(D9616_Y));
KC_BUF_X3 D8320 ( .Y(D8320_Y), .A(D8287_Y));
KC_BUF_X3 D8319 ( .Y(D8319_Y), .A(D8323_Y));
KC_BUF_X3 D8318 ( .Y(D8318_Y), .A(D7895_Y));
KC_BUF_X3 D8232 ( .Y(D8232_Y), .A(D8228_Y));
KC_BUF_X3 D8231 ( .Y(D8231_Y), .A(D8232_Y));
KC_BUF_X3 D8230 ( .Y(D8230_Y), .A(D8231_Y));
KC_BUF_X3 D8229 ( .Y(D8229_Y), .A(D8230_Y));
KC_BUF_X3 D8228 ( .Y(D8228_Y), .A(D8172_Y));
KC_BUF_X3 D8227 ( .Y(D8227_Y), .A(D8013_Y));
KC_BUF_X3 D8049 ( .Y(D8049_Y), .A(D621_Y));
KC_BUF_X3 D7880 ( .Y(D7880_Y), .A(D7795_Y));
KC_BUF_X3 D7649 ( .Y(D7649_Y), .A(D343_Y));
KC_BUF_X3 D7463 ( .Y(D7463_Y), .A(D7425_Y));
KC_BUF_X3 D7462 ( .Y(D7462_Y), .A(D13_Y));
KC_BUF_X3 D7133 ( .Y(D7133_Y), .A(D7245_Y));
KC_BUF_X3 D7132 ( .Y(D7132_Y), .A(D4198_Y));
KC_BUF_X3 D6958 ( .Y(D6958_Y), .A(D621_Y));
KC_BUF_X3 D6809 ( .Y(D6809_Y), .A(D6591_Y));
KC_BUF_X3 D6808 ( .Y(D6808_Y), .A(D6592_Y));
KC_BUF_X3 D6465 ( .Y(D6465_Y), .A(D1810_Y));
KC_BUF_X3 D6463 ( .Y(D6463_Y), .A(D7795_Y));
KC_BUF_X3 D6331 ( .Y(D6331_Y), .A(D6307_Y));
KC_BUF_X3 D6330 ( .Y(D6330_Y), .A(D7727_Y));
KC_BUF_X3 D6329 ( .Y(D6329_Y), .A(D4762_Y));
KC_BUF_X3 D6328 ( .Y(D6328_Y), .A(D6297_Y));
KC_BUF_X3 D6327 ( .Y(D6327_Y), .A(D6290_Y));
KC_BUF_X3 D6255 ( .Y(D6255_Y), .A(D16147_Y));
KC_BUF_X3 D6254 ( .Y(D6254_Y), .A(D6306_Y));
KC_BUF_X3 D5558 ( .Y(D5558_Y), .A(D621_Y));
KC_BUF_X3 D5461 ( .Y(D5461_Y), .A(D9555_Y));
KC_BUF_X3 D5392 ( .Y(D5392_Y), .A(D9555_Y));
KC_BUF_X3 D5391 ( .Y(D5391_Y), .A(D621_Y));
KC_BUF_X3 D5390 ( .Y(D5390_Y), .A(D621_Y));
KC_BUF_X3 D5389 ( .Y(D5389_Y), .A(D5102_Y));
KC_BUF_X3 D5388 ( .Y(D5388_Y), .A(D5104_Y));
KC_BUF_X3 D5387 ( .Y(D5387_Y), .A(D169_Y));
KC_BUF_X3 D5301 ( .Y(D5301_Y), .A(D8267_Y));
KC_BUF_X3 D5215 ( .Y(D5215_Y), .A(D621_Y));
KC_BUF_X3 D4627 ( .Y(D4627_Y), .A(D6213_Y));
KC_BUF_X3 D4548 ( .Y(D4548_Y), .A(D6031_Y));
KC_BUF_X3 D4547 ( .Y(D4547_Y), .A(D7816_Y));
KC_BUF_X3 D4546 ( .Y(D4546_Y), .A(D7820_Y));
KC_BUF_X3 D4385 ( .Y(D4385_Y), .A(D2873_Y));
KC_BUF_X3 D3862 ( .Y(D3862_Y), .A(D621_Y));
KC_BUF_X3 D3564 ( .Y(D3564_Y), .A(D1463_Y));
KC_BUF_X3 D3476 ( .Y(D3476_Y), .A(D3408_Y));
KC_BUF_X3 D3361 ( .Y(D3361_Y), .A(D6296_Y));
KC_BUF_X3 D3174 ( .Y(D3174_Y), .A(D6136_Y));
KC_BUF_X3 D3066 ( .Y(D3066_Y), .A(D1482_Y));
KC_BUF_X3 D3065 ( .Y(D3065_Y), .A(D3066_Y));
KC_BUF_X3 D3064 ( .Y(D3064_Y), .A(D3033_Y));
KC_BUF_X3 D3063 ( .Y(D3063_Y), .A(D3045_Y));
KC_BUF_X3 D3062 ( .Y(D3062_Y), .A(D4624_Y));
KC_BUF_X3 D2789 ( .Y(D2789_Y), .A(D2886_Q));
KC_BUF_X3 D2666 ( .Y(D2666_Y), .A(D15597_Y));
KC_BUF_X3 D2512 ( .Y(D2512_Y), .A(D14711_Y));
KC_BUF_X3 D2511 ( .Y(D2511_Y), .A(D13211_Q));
KC_BUF_X3 D2510 ( .Y(D2510_Y), .A(D14858_Y));
KC_BUF_X3 D2466 ( .Y(D2466_Y), .A(D13989_Q));
KC_BUF_X3 D2465 ( .Y(D2465_Y), .A(D691_Q));
KC_BUF_X3 D2464 ( .Y(D2464_Y), .A(D13239_Y));
KC_BUF_X3 D2463 ( .Y(D2463_Y), .A(D13992_Q));
KC_BUF_X3 D2341 ( .Y(D2341_Y), .A(D12168_Y));
KC_BUF_X3 D2340 ( .Y(D2340_Y), .A(D2341_Y));
KC_BUF_X3 D2339 ( .Y(D2339_Y), .A(D12157_Y));
KC_BUF_X3 D2338 ( .Y(D2338_Y), .A(D2337_Y));
KC_BUF_X3 D2337 ( .Y(D2337_Y), .A(D2336_Y));
KC_BUF_X3 D2336 ( .Y(D2336_Y), .A(D16128_Y));
KC_BUF_X3 D2244 ( .Y(D2244_Y), .A(D621_Y));
KC_BUF_X3 D2243 ( .Y(D2243_Y), .A(D169_Y));
KC_BUF_X3 D2242 ( .Y(D2242_Y), .A(D8267_Y));
KC_BUF_X3 D2149 ( .Y(D2149_Y), .A(D10282_Y));
KC_BUF_X3 D2148 ( .Y(D2148_Y), .A(D10329_Y));
KC_BUF_X3 D2147 ( .Y(D2147_Y), .A(D8958_Y));
KC_BUF_X3 D2070 ( .Y(D2070_Y), .A(D7313_Y));
KC_BUF_X3 D2069 ( .Y(D2069_Y), .A(D51_Y));
KC_BUF_X3 D2068 ( .Y(D2068_Y), .A(D106_Y));
KC_BUF_X3 D2067 ( .Y(D2067_Y), .A(D9605_Y));
KC_BUF_X3 D1919 ( .Y(D1919_Y), .A(D7974_Y));
KC_BUF_X3 D1769 ( .Y(D1769_Y), .A(D6143_Y));
KC_BUF_X3 D1628 ( .Y(D1628_Y), .A(D8267_Y));
KC_BUF_X3 D1482 ( .Y(D1482_Y), .A(D1481_Y));
KC_BUF_X3 D1481 ( .Y(D1481_Y), .A(D1626_Y));
KC_BUF_X3 D1480 ( .Y(D1480_Y), .A(D6137_Y));
KC_BUF_X3 D1479 ( .Y(D1479_Y), .A(D1465_Y));
KC_BUF_X3 D1478 ( .Y(D1478_Y), .A(D3939_Q));
KC_BUF_X3 D654 ( .Y(D654_Y), .A(D9449_Y));
KC_BUF_X3 D502 ( .Y(D502_Y), .A(D10119_Y));
KC_BUF_X3 D106 ( .Y(D106_Y), .A(D10370_Q));
KC_BUF_X3 D105 ( .Y(D105_Y), .A(D7554_Y));
KC_BUF_X2 D16720 ( .Y(D16720_Y), .A(D16715_Y));
KC_BUF_X2 D16704 ( .Y(D16704_Y), .A(D16772_Y));
KC_BUF_X2 D16697 ( .Y(D16697_Y), .A(D16772_Y));
KC_BUF_X2 D16649 ( .Y(D16649_Y), .A(D16639_Y));
KC_BUF_X2 D16575 ( .Y(D16575_Y), .A(D16588_Y));
KC_BUF_X2 D16455 ( .Y(D16455_Y), .A(D15867_Y));
KC_BUF_X2 D16349 ( .Y(D16349_Y), .A(D15867_Y));
KC_BUF_X2 D16348 ( .Y(D16348_Y), .A(D14157_QN));
KC_BUF_X2 D16308 ( .Y(D16308_Y), .A(D534_Y));
KC_BUF_X2 D16307 ( .Y(D16307_Y), .A(D16334_Y));
KC_BUF_X2 D16007 ( .Y(D16007_Y), .A(D15992_Q));
KC_BUF_X2 D15934 ( .Y(D15934_Y), .A(D14228_Y));
KC_BUF_X2 D15663 ( .Y(D15663_Y), .A(D13387_QN));
KC_BUF_X2 D15429 ( .Y(D15429_Y), .A(D15380_Y));
KC_BUF_X2 D15247 ( .Y(D15247_Y), .A(D9301_Y));
KC_BUF_X2 D15245 ( .Y(D15245_Y), .A(D9340_Y));
KC_BUF_X2 D15228 ( .Y(D15228_Y), .A(D13793_Y));
KC_BUF_X2 D15124 ( .Y(D15124_Y), .A(D15159_Y));
KC_BUF_X2 D15123 ( .Y(D15123_Y), .A(D15159_Y));
KC_BUF_X2 D14992 ( .Y(D14992_Y), .A(D14228_Y));
KC_BUF_X2 D14987 ( .Y(D14987_Y), .A(D14161_QN));
KC_BUF_X2 D14983 ( .Y(D14983_Y), .A(D14160_QN));
KC_BUF_X2 D14675 ( .Y(D14675_Y), .A(D14712_Y));
KC_BUF_X2 D14674 ( .Y(D14674_Y), .A(D14712_Y));
KC_BUF_X2 D14579 ( .Y(D14579_Y), .A(D507_QN));
KC_BUF_X2 D14469 ( .Y(D14469_Y), .A(D14160_QN));
KC_BUF_X2 D14466 ( .Y(D14466_Y), .A(D14161_QN));
KC_BUF_X2 D14231 ( .Y(D14231_Y), .A(D13390_QN));
KC_BUF_X2 D14229 ( .Y(D14229_Y), .A(D14157_QN));
KC_BUF_X2 D14228 ( .Y(D14228_Y), .A(D14158_QN));
KC_BUF_X2 D14156 ( .Y(D14156_Y), .A(D14155_Y));
KC_BUF_X2 D14155 ( .Y(D14155_Y), .A(D14154_Y));
KC_BUF_X2 D14154 ( .Y(D14154_Y), .A(D885_Y));
KC_BUF_X2 D13818 ( .Y(D13818_Y), .A(D13843_Y));
KC_BUF_X2 D13817 ( .Y(D13817_Y), .A(D13843_Y));
KC_BUF_X2 D13794 ( .Y(D13794_Y), .A(D14228_Y));
KC_BUF_X2 D13747 ( .Y(D13747_Y), .A(D14148_Y));
KC_BUF_X2 D13745 ( .Y(D13745_Y), .A(D13390_QN));
KC_BUF_X2 D13698 ( .Y(D13698_Y), .A(D14228_Y));
KC_BUF_X2 D13605 ( .Y(D13605_Y), .A(D1076_Y));
KC_BUF_X2 D13604 ( .Y(D13604_Y), .A(D1076_Y));
KC_BUF_X2 D13511 ( .Y(D13511_Y), .A(D14228_Y));
KC_BUF_X2 D13509 ( .Y(D13509_Y), .A(D12743_Y));
KC_BUF_X2 D13376 ( .Y(D13376_Y), .A(D12333_Y));
KC_BUF_X2 D13251 ( .Y(D13251_Y), .A(D12860_Y));
KC_BUF_X2 D13249 ( .Y(D13249_Y), .A(D13248_Y));
KC_BUF_X2 D13248 ( .Y(D13248_Y), .A(D1059_Y));
KC_BUF_X2 D13155 ( .Y(D13155_Y), .A(D10097_Y));
KC_BUF_X2 D13079 ( .Y(D13079_Y), .A(D13094_Y));
KC_BUF_X2 D12975 ( .Y(D12975_Y), .A(D14228_Y));
KC_BUF_X2 D12903 ( .Y(D12903_Y), .A(D13387_QN));
KC_BUF_X2 D12838 ( .Y(D12838_Y), .A(D12280_Y));
KC_BUF_X2 D12831 ( .Y(D12831_Y), .A(D13387_QN));
KC_BUF_X2 D12827 ( .Y(D12827_Y), .A(D13387_QN));
KC_BUF_X2 D12740 ( .Y(D12740_Y), .A(D13249_Y));
KC_BUF_X2 D12670 ( .Y(D12670_Y), .A(D10131_Y));
KC_BUF_X2 D12669 ( .Y(D12669_Y), .A(D12668_Y));
KC_BUF_X2 D12668 ( .Y(D12668_Y), .A(D833_Y));
KC_BUF_X2 D12267 ( .Y(D12267_Y), .A(D6248_Q));
KC_BUF_X2 D12263 ( .Y(D12263_Y), .A(D12304_Y));
KC_BUF_X2 D12262 ( .Y(D12262_Y), .A(D12304_Y));
KC_BUF_X2 D12112 ( .Y(D12112_Y), .A(D11612_Y));
KC_BUF_X2 D12084 ( .Y(D12084_Y), .A(D11567_Y));
KC_BUF_X2 D11711 ( .Y(D11711_Y), .A(D15004_Y));
KC_BUF_X2 D11651 ( .Y(D11651_Y), .A(D10179_Y));
KC_BUF_X2 D11625 ( .Y(D11625_Y), .A(D11617_Y));
KC_BUF_X2 D11624 ( .Y(D11624_Y), .A(D11636_Q));
KC_BUF_X2 D11622 ( .Y(D11622_Y), .A(D2284_Y));
KC_BUF_X2 D11621 ( .Y(D11621_Y), .A(D11618_Y));
KC_BUF_X2 D11620 ( .Y(D11620_Y), .A(D2285_Y));
KC_BUF_X2 D11618 ( .Y(D11618_Y), .A(D11620_Y));
KC_BUF_X2 D11617 ( .Y(D11617_Y), .A(D501_Y));
KC_BUF_X2 D11593 ( .Y(D11593_Y), .A(D11612_Y));
KC_BUF_X2 D11567 ( .Y(D11567_Y), .A(D9440_Y));
KC_BUF_X2 D11316 ( .Y(D11316_Y), .A(D11417_Y));
KC_BUF_X2 D11315 ( .Y(D11315_Y), .A(D11417_Y));
KC_BUF_X2 D11163 ( .Y(D11163_Y), .A(D6615_Y));
KC_BUF_X2 D11124 ( .Y(D11124_Y), .A(D11122_Y));
KC_BUF_X2 D11123 ( .Y(D11123_Y), .A(D10644_Y));
KC_BUF_X2 D11122 ( .Y(D11122_Y), .A(D11123_Y));
KC_BUF_X2 D11063 ( .Y(D11063_Y), .A(D9440_Y));
KC_BUF_X2 D11023 ( .Y(D11023_Y), .A(D11055_Y));
KC_BUF_X2 D11022 ( .Y(D11022_Y), .A(D11055_Y));
KC_BUF_X2 D10938 ( .Y(D10938_Y), .A(D9701_Y));
KC_BUF_X2 D10871 ( .Y(D10871_Y), .A(D9440_Y));
KC_BUF_X2 D10786 ( .Y(D10786_Y), .A(D9563_Y));
KC_BUF_X2 D10784 ( .Y(D10784_Y), .A(D10236_Y));
KC_BUF_X2 D10707 ( .Y(D10707_Y), .A(D10705_Y));
KC_BUF_X2 D10706 ( .Y(D10706_Y), .A(D11133_Y));
KC_BUF_X2 D10705 ( .Y(D10705_Y), .A(D10704_Y));
KC_BUF_X2 D10704 ( .Y(D10704_Y), .A(D652_Y));
KC_BUF_X2 D10648 ( .Y(D10648_Y), .A(D540_Q));
KC_BUF_X2 D10647 ( .Y(D10647_Y), .A(D10648_Y));
KC_BUF_X2 D10646 ( .Y(D10646_Y), .A(D10641_Y));
KC_BUF_X2 D10645 ( .Y(D10645_Y), .A(D10646_Y));
KC_BUF_X2 D10644 ( .Y(D10644_Y), .A(D10645_Y));
KC_BUF_X2 D10643 ( .Y(D10643_Y), .A(D10182_Y));
KC_BUF_X2 D10642 ( .Y(D10642_Y), .A(D10643_Y));
KC_BUF_X2 D10641 ( .Y(D10641_Y), .A(D10642_Y));
KC_BUF_X2 D10494 ( .Y(D10494_Y), .A(D9701_Y));
KC_BUF_X2 D10412 ( .Y(D10412_Y), .A(D9701_Y));
KC_BUF_X2 D10411 ( .Y(D10411_Y), .A(D9701_Y));
KC_BUF_X2 D10208 ( .Y(D10208_Y), .A(D709_Y));
KC_BUF_X2 D10182 ( .Y(D10182_Y), .A(D10647_Y));
KC_BUF_X2 D10156 ( .Y(D10156_Y), .A(D414_Q));
KC_BUF_X2 D10140 ( .Y(D10140_Y), .A(D442_Q));
KC_BUF_X2 D10005 ( .Y(D10005_Y), .A(D265_Q));
KC_BUF_X2 D9900 ( .Y(D9900_Y), .A(D8663_Y));
KC_BUF_X2 D9899 ( .Y(D9899_Y), .A(D8663_Y));
KC_BUF_X2 D9701 ( .Y(D9701_Y), .A(D9468_QN));
KC_BUF_X2 D9700 ( .Y(D9700_Y), .A(D8478_Y));
KC_BUF_X2 D9699 ( .Y(D9699_Y), .A(D9440_Y));
KC_BUF_X2 D9559 ( .Y(D9559_Y), .A(D9446_Y));
KC_BUF_X2 D9555 ( .Y(D9555_Y), .A(D1761_Y));
KC_BUF_X2 D9554 ( .Y(D9554_Y), .A(D8264_Y));
KC_BUF_X2 D9448 ( .Y(D9448_Y), .A(D9701_Y));
KC_BUF_X2 D9447 ( .Y(D9447_Y), .A(D1663_Y));
KC_BUF_X2 D9443 ( .Y(D9443_Y), .A(D9423_Y));
KC_BUF_X2 D9440 ( .Y(D9440_Y), .A(D11627_Y));
KC_BUF_X2 D9348 ( .Y(D9348_Y), .A(D9260_Q));
KC_BUF_X2 D9347 ( .Y(D9347_Y), .A(D11627_Y));
KC_BUF_X2 D9346 ( .Y(D9346_Y), .A(D11711_Y));
KC_BUF_X2 D9315 ( .Y(D9315_Y), .A(D2104_Q));
KC_BUF_X2 D9257 ( .Y(D9257_Y), .A(D9315_Y));
KC_BUF_X2 D9254 ( .Y(D9254_Y), .A(D7654_Y));
KC_BUF_X2 D9208 ( .Y(D9208_Y), .A(D9257_Y));
KC_BUF_X2 D8797 ( .Y(D8797_Y), .A(D7272_Y));
KC_BUF_X2 D8793 ( .Y(D8793_Y), .A(D9017_Y));
KC_BUF_X2 D8791 ( .Y(D8791_Y), .A(D431_Y));
KC_BUF_X2 D8790 ( .Y(D8790_Y), .A(D9099_Y));
KC_BUF_X2 D8696 ( .Y(D8696_Y), .A(D8696_A));
KC_BUF_X2 D8695 ( .Y(D8695_Y), .A(D8695_A));
KC_BUF_X2 D8692 ( .Y(D8692_Y), .A(D36_Y));
KC_BUF_X2 D8579 ( .Y(D8579_Y), .A(D8607_Y));
KC_BUF_X2 D8569 ( .Y(D8569_Y), .A(D8607_Y));
KC_BUF_X2 D8453 ( .Y(D8453_Y), .A(D10237_Y));
KC_BUF_X2 D8441 ( .Y(D8441_Y), .A(D9701_Y));
KC_BUF_X2 D8310 ( .Y(D8310_Y), .A(D947_Q));
KC_BUF_X2 D8222 ( .Y(D8222_Y), .A(D8045_Y));
KC_BUF_X2 D7962 ( .Y(D7962_Y), .A(D2174_Q));
KC_BUF_X2 D7712 ( .Y(D7712_Y), .A(D9224_Y));
KC_BUF_X2 D7706 ( .Y(D7706_Y), .A(D7686_Y));
KC_BUF_X2 D7704 ( .Y(D7704_Y), .A(D7690_Y));
KC_BUF_X2 D7575 ( .Y(D7575_Y), .A(D7712_Y));
KC_BUF_X2 D7574 ( .Y(D7574_Y), .A(D7577_S));
KC_BUF_X2 D7572 ( .Y(D7572_Y), .A(D4807_Y));
KC_BUF_X2 D7516 ( .Y(D7516_Y), .A(D5812_Y));
KC_BUF_X2 D7514 ( .Y(D7514_Y), .A(D102_Y));
KC_BUF_X2 D7381 ( .Y(D7381_Y), .A(D7588_Y));
KC_BUF_X2 D6954 ( .Y(D6954_Y), .A(D9701_Y));
KC_BUF_X2 D6889 ( .Y(D6889_Y), .A(D6856_Y));
KC_BUF_X2 D6798 ( .Y(D6798_Y), .A(D536_Y));
KC_BUF_X2 D6735 ( .Y(D6735_Y), .A(D9701_Y));
KC_BUF_X2 D6647 ( .Y(D6647_Y), .A(D8138_Y));
KC_BUF_X2 D6646 ( .Y(D6646_Y), .A(D16753_Y));
KC_BUF_X2 D6534 ( .Y(D6534_Y), .A(D6467_QN));
KC_BUF_X2 D6525 ( .Y(D6525_Y), .A(D6467_QN));
KC_BUF_X2 D6522 ( .Y(D6522_Y), .A(D16696_Y));
KC_BUF_X2 D6520 ( .Y(D6520_Y), .A(D16696_Y));
KC_BUF_X2 D6462 ( .Y(D6462_Y), .A(D6484_Y));
KC_BUF_X2 D6461 ( .Y(D6461_Y), .A(D6460_Y));
KC_BUF_X2 D6460 ( .Y(D6460_Y), .A(D6615_Y));
KC_BUF_X2 D6373 ( .Y(D6373_Y), .A(D14591_Y));
KC_BUF_X2 D6372 ( .Y(D6372_Y), .A(D14591_Y));
KC_BUF_X2 D6326 ( .Y(D6326_Y), .A(D6304_Y));
KC_BUF_X2 D6322 ( .Y(D6322_Y), .A(D6268_Y));
KC_BUF_X2 D6321 ( .Y(D6321_Y), .A(D4808_QN));
KC_BUF_X2 D6319 ( .Y(D6319_Y), .A(D9266_Y));
KC_BUF_X2 D6316 ( .Y(D6316_Y), .A(D11640_Q));
KC_BUF_X2 D6253 ( .Y(D6253_Y), .A(D6232_Y));
KC_BUF_X2 D6252 ( .Y(D6252_Y), .A(D7660_Y));
KC_BUF_X2 D6250 ( .Y(D6250_Y), .A(D6173_Y));
KC_BUF_X2 D6249 ( .Y(D6249_Y), .A(D6305_Y));
KC_BUF_X2 D6205 ( .Y(D6205_Y), .A(D6139_Y));
KC_BUF_X2 D6166 ( .Y(D6166_Y), .A(D1008_Y));
KC_BUF_X2 D6165 ( .Y(D6165_Y), .A(D6223_Y));
KC_BUF_X2 D6064 ( .Y(D6064_Y), .A(D6078_Y));
KC_BUF_X2 D5799 ( .Y(D5799_Y), .A(D226_QN));
KC_BUF_X2 D5557 ( .Y(D5557_Y), .A(D9440_Y));
KC_BUF_X2 D5460 ( .Y(D5460_Y), .A(D5489_Y));
KC_BUF_X2 D5459 ( .Y(D5459_Y), .A(D5489_Y));
KC_BUF_X2 D5383 ( .Y(D5383_Y), .A(D5343_Y));
KC_BUF_X2 D4799 ( .Y(D4799_Y), .A(D10633_Y));
KC_BUF_X2 D4717 ( .Y(D4717_Y), .A(D7134_Y));
KC_BUF_X2 D4716 ( .Y(D4716_Y), .A(D6197_Y));
KC_BUF_X2 D4714 ( .Y(D4714_Y), .A(D4668_Y));
KC_BUF_X2 D4618 ( .Y(D4618_Y), .A(D6197_Y));
KC_BUF_X2 D4545 ( .Y(D4545_Y), .A(D297_Q));
KC_BUF_X2 D4544 ( .Y(D4544_Y), .A(D302_Q));
KC_BUF_X2 D4543 ( .Y(D4543_Y), .A(D108_QN));
KC_BUF_X2 D4539 ( .Y(D4539_Y), .A(D3003_Q));
KC_BUF_X2 D4538 ( .Y(D4538_Y), .A(D2999_Q));
KC_BUF_X2 D4537 ( .Y(D4537_Y), .A(D4485_Q));
KC_BUF_X2 D4535 ( .Y(D4535_Y), .A(D40_Q));
KC_BUF_X2 D4534 ( .Y(D4534_Y), .A(D300_Q));
KC_BUF_X2 D4533 ( .Y(D4533_Y), .A(D2883_Q));
KC_BUF_X2 D4532 ( .Y(D4532_Y), .A(D301_Q));
KC_BUF_X2 D4531 ( .Y(D4531_Y), .A(D298_Q));
KC_BUF_X2 D4530 ( .Y(D4530_Y), .A(D4486_Q));
KC_BUF_X2 D4527 ( .Y(D4527_Y), .A(D4808_QN));
KC_BUF_X2 D4462 ( .Y(D4462_Y), .A(D226_QN));
KC_BUF_X2 D4461 ( .Y(D4461_Y), .A(D9358_Y));
KC_BUF_X2 D4459 ( .Y(D4459_Y), .A(D6128_Y));
KC_BUF_X2 D4106 ( .Y(D4106_Y), .A(D4431_Y));
KC_BUF_X2 D4039 ( .Y(D4039_Y), .A(D4072_Y));
KC_BUF_X2 D4038 ( .Y(D4038_Y), .A(D62_Y));
KC_BUF_X2 D4034 ( .Y(D4034_Y), .A(D4072_Y));
KC_BUF_X2 D3958 ( .Y(D3958_Y), .A(D4571_Y));
KC_BUF_X2 D3860 ( .Y(D3860_Y), .A(D6615_Y));
KC_BUF_X2 D3719 ( .Y(D3719_Y), .A(D4406_Y));
KC_BUF_X2 D3718 ( .Y(D3718_Y), .A(D4406_Y));
KC_BUF_X2 D3668 ( .Y(D3668_Y), .A(D1663_Y));
KC_BUF_X2 D3353 ( .Y(D3353_Y), .A(D4782_Y));
KC_BUF_X2 D3352 ( .Y(D3352_Y), .A(D3528_Y));
KC_BUF_X2 D3267 ( .Y(D3267_Y), .A(D6268_Y));
KC_BUF_X2 D3265 ( .Y(D3265_Y), .A(D1825_Y));
KC_BUF_X2 D3259 ( .Y(D3259_Y), .A(D3211_Y));
KC_BUF_X2 D3170 ( .Y(D3170_Y), .A(D6171_Y));
KC_BUF_X2 D3057 ( .Y(D3057_Y), .A(D3000_Q));
KC_BUF_X2 D3056 ( .Y(D3056_Y), .A(D3004_Q));
KC_BUF_X2 D3055 ( .Y(D3055_Y), .A(D3001_Q));
KC_BUF_X2 D3054 ( .Y(D3054_Y), .A(D3002_Q));
KC_BUF_X2 D3052 ( .Y(D3052_Y), .A(D3013_Y));
KC_BUF_X2 D3049 ( .Y(D3049_Y), .A(D7784_Y));
KC_BUF_X2 D2982 ( .Y(D2982_Y), .A(D6136_Y));
KC_BUF_X2 D2956 ( .Y(D2956_Y), .A(D6185_Y));
KC_BUF_X2 D2955 ( .Y(D2955_Y), .A(D2962_Y));
KC_BUF_X2 D2864 ( .Y(D2864_Y), .A(D108_QN));
KC_BUF_X2 D2788 ( .Y(D2788_Y), .A(D2770_Y));
KC_BUF_X2 D2783 ( .Y(D2783_Y), .A(D2744_Y));
KC_BUF_X2 D2717 ( .Y(D2717_Y), .A(D4086_Y));
KC_BUF_X2 D2694 ( .Y(D2694_Y), .A(D16715_Y));
KC_BUF_X2 D2631 ( .Y(D2631_Y), .A(D13390_QN));
KC_BUF_X2 D2586 ( .Y(D2586_Y), .A(D15867_Y));
KC_BUF_X2 D2571 ( .Y(D2571_Y), .A(D14501_Y));
KC_BUF_X2 D2568 ( .Y(D2568_Y), .A(D15867_Y));
KC_BUF_X2 D2460 ( .Y(D2460_Y), .A(D13214_QN));
KC_BUF_X2 D2458 ( .Y(D2458_Y), .A(D14156_Y));
KC_BUF_X2 D2285 ( .Y(D2285_Y), .A(D11622_Y));
KC_BUF_X2 D2284 ( .Y(D2284_Y), .A(D11637_Q));
KC_BUF_X2 D2211 ( .Y(D2211_Y), .A(D9701_Y));
KC_BUF_X2 D2144 ( .Y(D2144_Y), .A(D9209_Q));
KC_BUF_X2 D2059 ( .Y(D2059_Y), .A(D9701_Y));
KC_BUF_X2 D2056 ( .Y(D2056_Y), .A(D233_Q));
KC_BUF_X2 D1764 ( .Y(D1764_Y), .A(D1825_Y));
KC_BUF_X2 D1625 ( .Y(D1625_Y), .A(D6128_Y));
KC_BUF_X2 D1469 ( .Y(D1469_Y), .A(D3167_Y));
KC_BUF_X2 D1460 ( .Y(D1460_Y), .A(D4571_Y));
KC_BUF_X2 D1345 ( .Y(D1345_Y), .A(D14157_QN));
KC_BUF_X2 D885 ( .Y(D885_Y), .A(D13509_Y));
KC_BUF_X2 D884 ( .Y(D884_Y), .A(D9701_Y));
KC_BUF_X2 D767 ( .Y(D767_Y), .A(D9440_Y));
KC_BUF_X2 D652 ( .Y(D652_Y), .A(D10208_Y));
KC_BUF_X2 D501 ( .Y(D501_Y), .A(D11621_Y));
KC_BUF_X2 D499 ( .Y(D499_Y), .A(D13097_Q));
KC_BUF_X2 D316 ( .Y(D316_Y), .A(D4536_Y));
KC_BUF_X2 D315 ( .Y(D315_Y), .A(D299_Q));
KC_BUF_X2 D224 ( .Y(D224_Y), .A(D6275_Y));
KC_BUF_X2 D185 ( .Y(D185_Y), .A(D6275_Y));
KC_BUF_X2 D104 ( .Y(D104_Y), .A(D13094_Y));
KC_NOR2B_X1 D16680 ( .B(D16570_Y), .Y(D16680_Y), .AN(D16686_Y));
KC_NOR2B_X1 D16679 ( .B(D16570_Y), .Y(D16679_Y), .AN(D16685_Y));
KC_NOR2B_X1 D16678 ( .B(D16570_Y), .Y(D16678_Y), .AN(D16687_Y));
KC_NOR2B_X1 D16675 ( .B(D16570_Y), .Y(D16675_Y), .AN(D15435_Y));
KC_NOR2B_X1 D16674 ( .B(D16570_Y), .Y(D16674_Y), .AN(D16662_Y));
KC_NOR2B_X1 D16673 ( .B(D16570_Y), .Y(D16673_Y), .AN(D1399_Y));
KC_NOR2B_X1 D16651 ( .B(D16570_Y), .Y(D16651_Y), .AN(D16663_Y));
KC_NOR2B_X1 D16648 ( .B(D16570_Y), .Y(D16648_Y), .AN(D16664_Y));
KC_NOR2B_X1 D16627 ( .B(D16570_Y), .Y(D16627_Y), .AN(D2690_Y));
KC_NOR2B_X1 D16626 ( .B(D16570_Y), .Y(D16626_Y), .AN(D16638_Y));
KC_NOR2B_X1 D16625 ( .B(D16570_Y), .Y(D16625_Y), .AN(D1398_Y));
KC_NOR2B_X1 D16609 ( .B(D16599_Q), .Y(D16609_Y), .AN(D1396_Q));
KC_NOR2B_X1 D16548 ( .B(D16531_Y), .Y(D16548_Y), .AN(D16560_Y));
KC_NOR2B_X1 D16513 ( .B(D16469_Y), .Y(D16513_Y), .AN(D16510_Y));
KC_NOR2B_X1 D16512 ( .B(D1344_Y), .Y(D16512_Y), .AN(D16546_Y));
KC_NOR2B_X1 D16196 ( .B(D7609_Y), .Y(D16196_Y), .AN(D16225_Q));
KC_NOR2B_X1 D16138 ( .B(D7609_Y), .Y(D16138_Y), .AN(D16138_AN));
KC_NOR2B_X1 D16133 ( .B(D7609_Y), .Y(D16133_Y), .AN(D539_Q));
KC_NOR2B_X1 D16005 ( .B(D16078_Y), .Y(D16005_Y), .AN(D16004_Y));
KC_NOR2B_X1 D15784 ( .B(D2639_Q), .Y(D15784_Y), .AN(D925_Q));
KC_NOR2B_X1 D15006 ( .B(D1065_Q), .Y(D15006_Y), .AN(D1054_Q));
KC_NOR2B_X1 D14991 ( .B(D14903_Q), .Y(D14991_Y), .AN(D14874_Q));
KC_NOR2B_X1 D14077 ( .B(D14065_Y), .Y(D14077_Y), .AN(D2478_Y));
KC_NOR2B_X1 D13973 ( .B(D14017_Y), .Y(D13973_Y), .AN(D13993_Q));
KC_NOR2B_X1 D13853 ( .B(D14000_Y), .Y(D13853_Y), .AN(D13861_Y));
KC_NOR2B_X1 D13852 ( .B(D14000_Y), .Y(D13852_Y), .AN(D13862_Y));
KC_NOR2B_X1 D13851 ( .B(D14000_Y), .Y(D13851_Y), .AN(D2498_Y));
KC_NOR2B_X1 D13850 ( .B(D14000_Y), .Y(D13850_Y), .AN(D13863_Y));
KC_NOR2B_X1 D13849 ( .B(D14000_Y), .Y(D13849_Y), .AN(D10206_Y));
KC_NOR2B_X1 D13513 ( .B(D12861_Y), .Y(D13513_Y), .AN(D930_Q));
KC_NOR2B_X1 D13377 ( .B(D699_Q), .Y(D13377_Y), .AN(D12732_Y));
KC_NOR2B_X1 D13256 ( .B(D7609_Y), .Y(D13256_Y), .AN(D6107_Y));
KC_NOR2B_X1 D13252 ( .B(D13245_Y), .Y(D13252_Y), .AN(D13977_Y));
KC_NOR2B_X1 D12839 ( .B(D12837_Y), .Y(D12839_Y), .AN(D12697_Y));
KC_NOR2B_X1 D12828 ( .B(D12829_Y), .Y(D12828_Y), .AN(D12697_Y));
KC_NOR2B_X1 D12739 ( .B(D7305_Y), .Y(D12739_Y), .AN(D12260_Y));
KC_NOR2B_X1 D12220 ( .B(D12196_Y), .Y(D12220_Y), .AN(D10179_Y));
KC_NOR2B_X1 D12219 ( .B(D12196_Y), .Y(D12219_Y), .AN(D11657_Y));
KC_NOR2B_X1 D12217 ( .B(D12196_Y), .Y(D12217_Y), .AN(D11655_Y));
KC_NOR2B_X1 D12216 ( .B(D12196_Y), .Y(D12216_Y), .AN(D11660_Y));
KC_NOR2B_X1 D12215 ( .B(D12196_Y), .Y(D12215_Y), .AN(D9371_Y));
KC_NOR2B_X1 D12138 ( .B(D12183_Y), .Y(D12138_Y), .AN(D11672_Q));
KC_NOR2B_X1 D12040 ( .B(D8465_Y), .Y(D12040_Y), .AN(D1246_Q));
KC_NOR2B_X1 D12037 ( .B(D8465_Y), .Y(D12037_Y), .AN(D1224_Q));
KC_NOR2B_X1 D12034 ( .B(D8465_Y), .Y(D12034_Y), .AN(D12043_Q));
KC_NOR2B_X1 D12033 ( .B(D8465_Y), .Y(D12033_Y), .AN(D12042_Q));
KC_NOR2B_X1 D11845 ( .B(D2222_Y), .Y(D11845_Y), .AN(D11859_Q));
KC_NOR2B_X1 D11780 ( .B(D2222_Y), .Y(D11780_Y), .AN(D136_Q));
KC_NOR2B_X1 D11619 ( .B(D2304_Q), .Y(D11619_Y), .AN(D8903_Y));
KC_NOR2B_X1 D11533 ( .B(D8465_Y), .Y(D11533_Y), .AN(D11543_Q));
KC_NOR2B_X1 D11530 ( .B(D8465_Y), .Y(D11530_Y), .AN(D1219_Q));
KC_NOR2B_X1 D11529 ( .B(D8465_Y), .Y(D11529_Y), .AN(D11542_Q));
KC_NOR2B_X1 D11528 ( .B(D8465_Y), .Y(D11528_Y), .AN(D11541_Q));
KC_NOR2B_X1 D11527 ( .B(D8465_Y), .Y(D11527_Y), .AN(D11537_Q));
KC_NOR2B_X1 D11464 ( .B(D8465_Y), .Y(D11464_Y), .AN(D1218_Q));
KC_NOR2B_X1 D11463 ( .B(D8465_Y), .Y(D11463_Y), .AN(D2251_Q));
KC_NOR2B_X1 D11462 ( .B(D8465_Y), .Y(D11462_Y), .AN(D131_Q));
KC_NOR2B_X1 D11461 ( .B(D8465_Y), .Y(D11461_Y), .AN(D2249_Q));
KC_NOR2B_X1 D11460 ( .B(D8465_Y), .Y(D11460_Y), .AN(D11539_Q));
KC_NOR2B_X1 D11459 ( .B(D8465_Y), .Y(D11459_Y), .AN(D2250_Q));
KC_NOR2B_X1 D11457 ( .B(D8465_Y), .Y(D11457_Y), .AN(D11469_Q));
KC_NOR2B_X1 D11452 ( .B(D8465_Y), .Y(D11452_Y), .AN(D2253_Q));
KC_NOR2B_X1 D11450 ( .B(D8465_Y), .Y(D11450_Y), .AN(D11466_Q));
KC_NOR2B_X1 D11448 ( .B(D8465_Y), .Y(D11448_Y), .AN(D11468_Q));
KC_NOR2B_X1 D11320 ( .B(D2222_Y), .Y(D11320_Y), .AN(D11341_Q));
KC_NOR2B_X1 D11319 ( .B(D2222_Y), .Y(D11319_Y), .AN(D11326_Q));
KC_NOR2B_X1 D11318 ( .B(D2222_Y), .Y(D11318_Y), .AN(D11392_Q));
KC_NOR2B_X1 D11314 ( .B(D2222_Y), .Y(D11314_Y), .AN(D11342_Q));
KC_NOR2B_X1 D11313 ( .B(D2222_Y), .Y(D11313_Y), .AN(D11340_Q));
KC_NOR2B_X1 D11251 ( .B(D2222_Y), .Y(D11251_Y), .AN(D11262_Q));
KC_NOR2B_X1 D11250 ( .B(D2222_Y), .Y(D11250_Y), .AN(D11264_Q));
KC_NOR2B_X1 D11249 ( .B(D2222_Y), .Y(D11249_Y), .AN(D11265_Q));
KC_NOR2B_X1 D11245 ( .B(D2222_Y), .Y(D11245_Y), .AN(D11263_Q));
KC_NOR2B_X1 D11242 ( .B(D2222_Y), .Y(D11242_Y), .AN(D11261_Q));
KC_NOR2B_X1 D11240 ( .B(D2222_Y), .Y(D11240_Y), .AN(D2256_Q));
KC_NOR2B_X1 D10780 ( .B(D2222_Y), .Y(D10780_Y), .AN(D797_Q));
KC_NOR2B_X1 D10779 ( .B(D2202_Y), .Y(D10779_Y), .AN(D10793_Q));
KC_NOR2B_X1 D10778 ( .B(D2202_Y), .Y(D10778_Y), .AN(D10791_Q));
KC_NOR2B_X1 D10777 ( .B(D2202_Y), .Y(D10777_Y), .AN(D10789_Q));
KC_NOR2B_X1 D10505 ( .B(D8363_Y), .Y(D10505_Y), .AN(D10978_Y));
KC_NOR2B_X1 D10209 ( .B(D10218_Q), .Y(D10209_Y), .AN(D10217_Q));
KC_NOR2B_X1 D10141 ( .B(D2162_Y), .Y(D10141_Y), .AN(D10033_Q));
KC_NOR2B_X1 D9558 ( .B(D9513_Y), .Y(D9558_Y), .AN(D9505_Y));
KC_NOR2B_X1 D9556 ( .B(D8175_Y), .Y(D9556_Y), .AN(D837_Q));
KC_NOR2B_X1 D9255 ( .B(D9234_Y), .Y(D9255_Y), .AN(D9282_Y));
KC_NOR2B_X1 D9205 ( .B(D70_Y), .Y(D9205_Y), .AN(D2002_Y));
KC_NOR2B_X1 D9000 ( .B(D9159_Q), .Y(D9000_Y), .AN(D9216_Q));
KC_NOR2B_X1 D8794 ( .B(D8798_S), .Y(D8794_Y), .AN(D8774_Y));
KC_NOR2B_X1 D8788 ( .B(D8772_Y), .Y(D8788_Y), .AN(D8754_Y));
KC_NOR2B_X1 D8693 ( .B(D188_Y), .Y(D8693_Y), .AN(D9928_Y));
KC_NOR2B_X1 D8690 ( .B(D190_Y), .Y(D8690_Y), .AN(D8675_Y));
KC_NOR2B_X1 D8582 ( .B(D8422_Y), .Y(D8582_Y), .AN(D8589_Q));
KC_NOR2B_X1 D8578 ( .B(D8422_Y), .Y(D8578_Y), .AN(D7005_Q));
KC_NOR2B_X1 D8577 ( .B(D8422_Y), .Y(D8577_Y), .AN(D1927_Q));
KC_NOR2B_X1 D8576 ( .B(D8422_Y), .Y(D8576_Y), .AN(D8594_Q));
KC_NOR2B_X1 D8528 ( .B(D8422_Y), .Y(D8528_Y), .AN(D8538_Q));
KC_NOR2B_X1 D8448 ( .B(D8395_Y), .Y(D8448_Y), .AN(D1779_Q));
KC_NOR2B_X1 D8439 ( .B(D8395_Y), .Y(D8439_Y), .AN(D1928_Q));
KC_NOR2B_X1 D8306 ( .B(D1932_Y), .Y(D8306_Y), .AN(D6829_Q));
KC_NOR2B_X1 D8305 ( .B(D1932_Y), .Y(D8305_Y), .AN(D6825_Q));
KC_NOR2B_X1 D8304 ( .B(D1932_Y), .Y(D8304_Y), .AN(D1930_Q));
KC_NOR2B_X1 D8226 ( .B(D9559_Y), .Y(D8226_Y), .AN(D8261_Y));
KC_NOR2B_X1 D8225 ( .B(D8219_Y), .Y(D8225_Y), .AN(D8190_Y));
KC_NOR2B_X1 D8224 ( .B(D9559_Y), .Y(D8224_Y), .AN(D8261_Y));
KC_NOR2B_X1 D8141 ( .B(D8007_Y), .Y(D8141_Y), .AN(D676_Q));
KC_NOR2B_X1 D8138 ( .B(D8109_Y), .Y(D8138_Y), .AN(D4137_Q));
KC_NOR2B_X1 D8043 ( .B(D8007_Y), .Y(D8043_Y), .AN(D669_Q));
KC_NOR2B_X1 D8041 ( .B(D8007_Y), .Y(D8041_Y), .AN(D8052_Q));
KC_NOR2B_X1 D8040 ( .B(D8007_Y), .Y(D8040_Y), .AN(D8054_Q));
KC_NOR2B_X1 D8037 ( .B(D8007_Y), .Y(D8037_Y), .AN(D8053_Q));
KC_NOR2B_X1 D8036 ( .B(D8007_Y), .Y(D8036_Y), .AN(D8055_Q));
KC_NOR2B_X1 D8033 ( .B(D8007_Y), .Y(D8033_Y), .AN(D672_Q));
KC_NOR2B_X1 D7960 ( .B(D6431_Y), .Y(D7960_Y), .AN(D7915_Y));
KC_NOR2B_X1 D7959 ( .B(D8044_Y), .Y(D7959_Y), .AN(D8272_Y));
KC_NOR2B_X1 D7958 ( .B(D8044_Y), .Y(D7958_Y), .AN(D8277_Y));
KC_NOR2B_X1 D7957 ( .B(D8044_Y), .Y(D7957_Y), .AN(D8270_Y));
KC_NOR2B_X1 D7877 ( .B(D7830_Y), .Y(D7877_Y), .AN(D7953_Y));
KC_NOR2B_X1 D7875 ( .B(D1852_Y), .Y(D7875_Y), .AN(D7838_Y));
KC_NOR2B_X1 D7780 ( .B(D9281_Y), .Y(D7780_Y), .AN(D9241_Y));
KC_NOR2B_X1 D7779 ( .B(D382_Y), .Y(D7779_Y), .AN(D18_Y));
KC_NOR2B_X1 D7710 ( .B(D7751_Q), .Y(D7710_Y), .AN(D7732_Q));
KC_NOR2B_X1 D7709 ( .B(D7742_Q), .Y(D7709_Y), .AN(D7733_Q));
KC_NOR2B_X1 D7648 ( .B(D7686_Y), .Y(D7648_Y), .AN(D7642_Y));
KC_NOR2B_X1 D7460 ( .B(D7402_Y), .Y(D7460_Y), .AN(D9473_Y));
KC_NOR2B_X1 D7459 ( .B(D23_Y), .Y(D7459_Y), .AN(D7505_Y));
KC_NOR2B_X1 D7382 ( .B(D7381_Y), .Y(D7382_Y), .AN(D5908_Y));
KC_NOR2B_X1 D7380 ( .B(D5827_Y), .Y(D7380_Y), .AN(D8050_Y));
KC_NOR2B_X1 D7290 ( .B(D7240_Y), .Y(D7290_Y), .AN(D7215_Y));
KC_NOR2B_X1 D7288 ( .B(D7183_Y), .Y(D7288_Y), .AN(D7166_Y));
KC_NOR2B_X1 D7130 ( .B(D7116_Y), .Y(D7130_Y), .AN(D7115_Y));
KC_NOR2B_X1 D6953 ( .B(D8395_Y), .Y(D6953_Y), .AN(D1126_Q));
KC_NOR2B_X1 D6951 ( .B(D8395_Y), .Y(D6951_Y), .AN(D6970_Q));
KC_NOR2B_X1 D6948 ( .B(D8395_Y), .Y(D6948_Y), .AN(D1774_Q));
KC_NOR2B_X1 D6804 ( .B(D1932_Y), .Y(D6804_Y), .AN(D8238_Q));
KC_NOR2B_X1 D6801 ( .B(D1932_Y), .Y(D6801_Y), .AN(D6826_Q));
KC_NOR2B_X1 D6800 ( .B(D6260_Y), .Y(D6800_Y), .AN(D8031_Y));
KC_NOR2B_X1 D6741 ( .B(D1932_Y), .Y(D6741_Y), .AN(D796_Q));
KC_NOR2B_X1 D6740 ( .B(D1932_Y), .Y(D6740_Y), .AN(D6750_Q));
KC_NOR2B_X1 D6737 ( .B(D1932_Y), .Y(D6737_Y), .AN(D6754_Q));
KC_NOR2B_X1 D6734 ( .B(D1932_Y), .Y(D6734_Y), .AN(D6744_Q));
KC_NOR2B_X1 D6733 ( .B(D1932_Y), .Y(D6733_Y), .AN(D789_Q));
KC_NOR2B_X1 D6730 ( .B(D1932_Y), .Y(D6730_Y), .AN(D785_Q));
KC_NOR2B_X1 D6651 ( .B(D1932_Y), .Y(D6651_Y), .AN(D8051_Q));
KC_NOR2B_X1 D6644 ( .B(D1932_Y), .Y(D6644_Y), .AN(D6758_Q));
KC_NOR2B_X1 D6643 ( .B(D1932_Y), .Y(D6643_Y), .AN(D664_Q));
KC_NOR2B_X1 D6371 ( .B(D153_Q), .Y(D6371_Y), .AN(D1847_Y));
KC_NOR2B_X1 D6325 ( .B(D6330_Y), .Y(D6325_Y), .AN(D6315_Y));
KC_NOR2B_X1 D6324 ( .B(D1945_Y), .Y(D6324_Y), .AN(D427_Q));
KC_NOR2B_X1 D6323 ( .B(D1945_Y), .Y(D6323_Y), .AN(D429_Q));
KC_NOR2B_X1 D6317 ( .B(D1945_Y), .Y(D6317_Y), .AN(D6359_Q));
KC_NOR2B_X1 D6168 ( .B(D6196_Y), .Y(D6168_Y), .AN(D6167_Y));
KC_NOR2B_X1 D6114 ( .B(D8838_Y), .Y(D6114_Y), .AN(D266_Y));
KC_NOR2B_X1 D6113 ( .B(D4489_Q), .Y(D6113_Y), .AN(D12678_Y));
KC_NOR2B_X1 D6071 ( .B(D1724_Y), .Y(D6071_Y), .AN(D288_Y));
KC_NOR2B_X1 D6068 ( .B(D5970_Y), .Y(D6068_Y), .AN(D5982_Y));
KC_NOR2B_X1 D6065 ( .B(D4409_Y), .Y(D6065_Y), .AN(D5962_Y));
KC_NOR2B_X1 D5925 ( .B(D5841_Y), .Y(D5925_Y), .AN(D5980_Y));
KC_NOR2B_X1 D5678 ( .B(D5675_Y), .Y(D5678_Y), .AN(D5689_Q));
KC_NOR2B_X1 D5677 ( .B(D5676_Y), .Y(D5677_Y), .AN(D5652_Y));
KC_NOR2B_X1 D5073 ( .B(D5067_Y), .Y(D5073_Y), .AN(D5030_Y));
KC_NOR2B_X1 D4952 ( .B(D6381_Q), .Y(D4952_Y), .AN(D6371_Y));
KC_NOR2B_X1 D4803 ( .B(D4772_Y), .Y(D4803_Y), .AN(D4828_Y));
KC_NOR2B_X1 D4802 ( .B(D4835_Y), .Y(D4802_Y), .AN(D4779_Y));
KC_NOR2B_X1 D4800 ( .B(D413_Y), .Y(D4800_Y), .AN(D4833_Y));
KC_NOR2B_X1 D4797 ( .B(D4780_Y), .Y(D4797_Y), .AN(D4812_Y));
KC_NOR2B_X1 D4795 ( .B(D413_Y), .Y(D4795_Y), .AN(D425_Y));
KC_NOR2B_X1 D4794 ( .B(D413_Y), .Y(D4794_Y), .AN(D4831_Y));
KC_NOR2B_X1 D4793 ( .B(D413_Y), .Y(D4793_Y), .AN(D4832_Y));
KC_NOR2B_X1 D4792 ( .B(D413_Y), .Y(D4792_Y), .AN(D4829_Y));
KC_NOR2B_X1 D4791 ( .B(D413_Y), .Y(D4791_Y), .AN(D4550_Y));
KC_NOR2B_X1 D4790 ( .B(D413_Y), .Y(D4790_Y), .AN(D4830_Y));
KC_NOR2B_X1 D4711 ( .B(D4712_Y), .Y(D4711_Y), .AN(D4702_Y));
KC_NOR2B_X1 D4626 ( .B(D1945_Y), .Y(D4626_Y), .AN(D4649_Q));
KC_NOR2B_X1 D4624 ( .B(D1945_Y), .Y(D4624_Y), .AN(D4641_Q));
KC_NOR2B_X1 D4623 ( .B(D4610_Y), .Y(D4623_Y), .AN(D4651_Y));
KC_NOR2B_X1 D4621 ( .B(D4633_Y), .Y(D4621_Y), .AN(D4623_Y));
KC_NOR2B_X1 D4536 ( .B(D1945_Y), .Y(D4536_Y), .AN(D4467_Y));
KC_NOR2B_X1 D4529 ( .B(D1945_Y), .Y(D4529_Y), .AN(D4560_Q));
KC_NOR2B_X1 D4528 ( .B(D3026_Y), .Y(D4528_Y), .AN(D3024_Y));
KC_NOR2B_X1 D4460 ( .B(D4482_Y), .Y(D4460_Y), .AN(D4492_Y));
KC_NOR2B_X1 D4384 ( .B(D4348_Y), .Y(D4384_Y), .AN(D4345_Y));
KC_NOR2B_X1 D4381 ( .B(D4314_Y), .Y(D4381_Y), .AN(D4283_Y));
KC_NOR2B_X1 D4380 ( .B(D165_Y), .Y(D4380_Y), .AN(D4456_Y));
KC_NOR2B_X1 D4110 ( .B(D4104_Y), .Y(D4110_Y), .AN(D4103_Y));
KC_NOR2B_X1 D4109 ( .B(D16135_Y), .Y(D4109_Y), .AN(D4123_Y));
KC_NOR2B_X1 D3623 ( .B(D1953_Y), .Y(D3623_Y), .AN(D3638_Q));
KC_NOR2B_X1 D3621 ( .B(D1953_Y), .Y(D3621_Y), .AN(D3635_Q));
KC_NOR2B_X1 D3620 ( .B(D1953_Y), .Y(D3620_Y), .AN(D1518_Q));
KC_NOR2B_X1 D3619 ( .B(D1953_Y), .Y(D3619_Y), .AN(D3637_Q));
KC_NOR2B_X1 D3617 ( .B(D1953_Y), .Y(D3617_Y), .AN(D3645_Q));
KC_NOR2B_X1 D3616 ( .B(D1953_Y), .Y(D3616_Y), .AN(D3648_Q));
KC_NOR2B_X1 D3615 ( .B(D1953_Y), .Y(D3615_Y), .AN(D3636_Q));
KC_NOR2B_X1 D3614 ( .B(D1953_Y), .Y(D3614_Y), .AN(D3646_Q));
KC_NOR2B_X1 D3613 ( .B(D1953_Y), .Y(D3613_Y), .AN(D3642_Q));
KC_NOR2B_X1 D3612 ( .B(D1953_Y), .Y(D3612_Y), .AN(D3640_Q));
KC_NOR2B_X1 D3608 ( .B(D1953_Y), .Y(D3608_Y), .AN(D3641_Q));
KC_NOR2B_X1 D3606 ( .B(D1953_Y), .Y(D3606_Y), .AN(D3643_Q));
KC_NOR2B_X1 D3605 ( .B(D1953_Y), .Y(D3605_Y), .AN(D3644_Q));
KC_NOR2B_X1 D3559 ( .B(D3517_Y), .Y(D3559_Y), .AN(D3571_Y));
KC_NOR2B_X1 D3472 ( .B(D3476_Y), .Y(D3472_Y), .AN(D3411_Y));
KC_NOR2B_X1 D3360 ( .B(D3369_Y), .Y(D3360_Y), .AN(D3323_Y));
KC_NOR2B_X1 D3359 ( .B(D3357_Y), .Y(D3359_Y), .AN(D3314_Y));
KC_NOR2B_X1 D3358 ( .B(D413_Y), .Y(D3358_Y), .AN(D426_Y));
KC_NOR2B_X1 D3357 ( .B(D3342_Y), .Y(D3357_Y), .AN(D1454_Y));
KC_NOR2B_X1 D3268 ( .B(D2995_Y), .Y(D3268_Y), .AN(D4718_S));
KC_NOR2B_X1 D3266 ( .B(D1480_Y), .Y(D3266_Y), .AN(D3265_Y));
KC_NOR2B_X1 D3261 ( .B(D3245_Y), .Y(D3261_Y), .AN(D3360_Y));
KC_NOR2B_X1 D3258 ( .B(D3350_Y), .Y(D3258_Y), .AN(D3329_Y));
KC_NOR2B_X1 D3172 ( .B(D3132_Y), .Y(D3172_Y), .AN(D3140_Y));
KC_NOR2B_X1 D3168 ( .B(D7641_Y), .Y(D3168_Y), .AN(D3105_Y));
KC_NOR2B_X1 D3053 ( .B(D3087_Y), .Y(D3053_Y), .AN(D3064_Y));
KC_NOR2B_X1 D3047 ( .B(D7641_Y), .Y(D3047_Y), .AN(D1608_Y));
KC_NOR2B_X1 D2873 ( .B(D4392_Y), .Y(D2873_Y), .AN(D4310_Y));
KC_NOR2B_X1 D2867 ( .B(D2868_Y), .Y(D2867_Y), .AN(D2853_Y));
KC_NOR2B_X1 D2784 ( .B(D2772_Y), .Y(D2784_Y), .AN(D2901_Y));
KC_NOR2B_X1 D2632 ( .B(D14871_Q), .Y(D2632_Y), .AN(D15670_Q));
KC_NOR2B_X1 D2282 ( .B(D2222_Y), .Y(D2282_Y), .AN(D11260_Q));
KC_NOR2B_X1 D2241 ( .B(D2222_Y), .Y(D2241_Y), .AN(D11328_Q));
KC_NOR2B_X1 D2240 ( .B(D2222_Y), .Y(D2240_Y), .AN(D11327_Q));
KC_NOR2B_X1 D2237 ( .B(D2202_Y), .Y(D2237_Y), .AN(D11389_Q));
KC_NOR2B_X1 D2212 ( .B(D2222_Y), .Y(D2212_Y), .AN(D135_Q));
KC_NOR2B_X1 D2210 ( .B(D2202_Y), .Y(D2210_Y), .AN(D10790_Q));
KC_NOR2B_X1 D2209 ( .B(D2202_Y), .Y(D2209_Y), .AN(D2221_Q));
KC_NOR2B_X1 D2146 ( .B(D2135_Y), .Y(D2146_Y), .AN(D98_Y));
KC_NOR2B_X1 D2063 ( .B(D263_Y), .Y(D2063_Y), .AN(D16_Y));
KC_NOR2B_X1 D2061 ( .B(D1895_Y), .Y(D2061_Y), .AN(D10361_Q));
KC_NOR2B_X1 D2058 ( .B(D8717_Y), .Y(D2058_Y), .AN(D8672_Y));
KC_NOR2B_X1 D1917 ( .B(D7865_Y), .Y(D1917_Y), .AN(D7985_Y));
KC_NOR2B_X1 D1915 ( .B(D8246_Q), .Y(D1915_Y), .AN(D8201_Y));
KC_NOR2B_X1 D1765 ( .B(D4804_Y), .Y(D1765_Y), .AN(D1764_Y));
KC_NOR2B_X1 D1758 ( .B(D1932_Y), .Y(D1758_Y), .AN(D784_Q));
KC_NOR2B_X1 D1755 ( .B(D8395_Y), .Y(D1755_Y), .AN(D7008_Q));
KC_NOR2B_X1 D1627 ( .B(D6010_Y), .Y(D1627_Y), .AN(D5726_Y));
KC_NOR2B_X1 D1534 ( .B(D1953_Y), .Y(D1534_Y), .AN(D3579_Q));
KC_NOR2B_X1 D1467 ( .B(D4948_Y), .Y(D1467_Y), .AN(D5005_Y));
KC_NOR2B_X1 D1465 ( .B(D3634_Y), .Y(D1465_Y), .AN(D3500_Y));
KC_NOR2B_X1 D1464 ( .B(D1953_Y), .Y(D1464_Y), .AN(D3580_Q));
KC_NOR2B_X1 D1462 ( .B(D1953_Y), .Y(D1462_Y), .AN(D3700_Q));
KC_NOR2B_X1 D1461 ( .B(D1953_Y), .Y(D1461_Y), .AN(D3639_Q));
KC_NOR2B_X1 D1195 ( .B(D8465_Y), .Y(D1195_Y), .AN(D11538_Q));
KC_NOR2B_X1 D1111 ( .B(D15835_Y), .Y(D1111_Y), .AN(D2678_Q));
KC_NOR2B_X1 D890 ( .B(D2222_Y), .Y(D890_Y), .AN(D11329_Q));
KC_NOR2B_X1 D886 ( .B(D2395_Y), .Y(D886_Y), .AN(D954_Q));
KC_NOR2B_X1 D881 ( .B(D1932_Y), .Y(D881_Y), .AN(D8459_Q));
KC_NOR2B_X1 D880 ( .B(D1932_Y), .Y(D880_Y), .AN(D903_Q));
KC_NOR2B_X1 D772 ( .B(D2222_Y), .Y(D772_Y), .AN(D10792_Q));
KC_NOR2B_X1 D768 ( .B(D13302_Y), .Y(D768_Y), .AN(D12279_Q));
KC_NOR2B_X1 D581 ( .B(D7782_Y), .Y(D581_Y), .AN(D9341_Y));
KC_NOR2B_X1 D500 ( .B(D14000_Y), .Y(D500_Y), .AN(D13174_Y));
KC_NOR2B_X1 D413 ( .B(D369_Y), .Y(D413_Y), .AN(D3321_Y));
KC_NOR2B_X1 D412 ( .B(D413_Y), .Y(D412_Y), .AN(D4834_Y));
KC_NOR2B_X1 D187 ( .B(D8693_Y), .Y(D187_Y), .AN(D8686_Y));
KC_NOR2B_X1 D102 ( .B(D235_Y), .Y(D102_Y), .AN(D6114_Y));
KC_MXI2_X1 D15561 ( .Y(D15561_Y), .A(D15350_Y), .BN(D15402_Y),     .S0(D15554_Y));
KC_MXI2_X1 D15560 ( .Y(D15560_Y), .A(D15483_Y), .BN(D2614_Y),     .S0(D14862_Y));
KC_MXI2_X1 D14985 ( .Y(D14985_Y), .A(D14872_Q), .BN(D16315_Q),     .S0(D16362_Q));
KC_MXI2_X1 D14812 ( .Y(D14812_Y), .A(D16234_Y), .BN(D14889_Y),     .S0(D13971_Y));
KC_MXI2_X1 D14783 ( .Y(D14783_Y), .A(D720_Y), .BN(D14191_Y),     .S0(D13971_Y));
KC_MXI2_X1 D14782 ( .Y(D14782_Y), .A(D846_Y), .BN(D14192_Y),     .S0(D13971_Y));
KC_MXI2_X1 D14781 ( .Y(D14781_Y), .A(D16235_Y), .BN(D14892_Y),     .S0(D13971_Y));
KC_MXI2_X1 D14780 ( .Y(D14780_Y), .A(D16228_Y), .BN(D14898_Y),     .S0(D13971_Y));
KC_MXI2_X1 D14779 ( .Y(D14779_Y), .A(D16230_Y), .BN(D14902_Y),     .S0(D13971_Y));
KC_MXI2_X1 D14778 ( .Y(D14778_Y), .A(D16241_Y), .BN(D14899_Y),     .S0(D13971_Y));
KC_MXI2_X1 D14232 ( .Y(D14232_Y), .A(D1066_Q), .BN(D14236_Q),     .S0(D14243_Q));
KC_MXI2_X1 D12837 ( .Y(D12837_Y), .A(D12858_Q), .BN(D12259_Y),     .S0(D13348_Y));
KC_MXI2_X1 D12829 ( .Y(D12829_Y), .A(D12855_Q), .BN(D12257_Y),     .S0(D13221_Y));
KC_MXI2_X1 D10322 ( .Y(D10322_Y), .A(D10361_Q), .BN(D10361_Q),     .S0(D10318_Y));
KC_MXI2_X1 D9259 ( .Y(D9259_Y), .A(D9222_Y), .BN(D9243_Y),     .S0(D163_Y));
KC_MXI2_X1 D8796 ( .Y(D8796_Y), .A(D8805_Y), .BN(D8774_Y),     .S0(D8755_Y));
KC_MXI2_X1 D8133 ( .Y(D8133_Y), .A(D8092_Y), .BN(D8148_Q),     .S0(D8090_Y));
KC_MXI2_X1 D8048 ( .Y(D8048_Y), .A(D7670_Y), .BN(D7971_Q),     .S0(D8073_Q));
KC_MXI2_X1 D8047 ( .Y(D8047_Y), .A(D7668_Y), .BN(D7970_Q),     .S0(D8073_Q));
KC_MXI2_X1 D8045 ( .Y(D8045_Y), .A(D392_Y), .BN(D6472_Q),     .S0(D8073_Q));
KC_MXI2_X1 D8034 ( .Y(D8034_Y), .A(D6288_Y), .BN(D7969_Q),     .S0(D8073_Q));
KC_MXI2_X1 D7387 ( .Y(D7387_Y), .A(D5938_Y), .BN(D8903_Y),     .S0(D5915_Y));
KC_MXI2_X1 D6592 ( .Y(D6592_Y), .A(D6287_Y), .BN(D6474_Q),     .S0(D8073_Q));
KC_MXI2_X1 D6591 ( .Y(D6591_Y), .A(D6281_Y), .BN(D6476_Q),     .S0(D8073_Q));
KC_MXI2_X1 D6521 ( .Y(D6521_Y), .A(D392_Y), .BN(D523_Q), .S0(D8073_Q));
KC_MXI2_X1 D6110 ( .Y(D6110_Y), .A(D332_Y), .BN(D6085_Y),     .S0(D6813_Y));
KC_MXI2_X1 D5122 ( .Y(D5122_Y), .A(D6505_Y), .BN(D1644_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5121 ( .Y(D5121_Y), .A(D6509_Y), .BN(D5140_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5120 ( .Y(D5120_Y), .A(D6509_Y), .BN(D5078_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5119 ( .Y(D5119_Y), .A(D6506_Y), .BN(D522_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5118 ( .Y(D5118_Y), .A(D6508_Y), .BN(D5137_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5117 ( .Y(D5117_Y), .A(D6508_Y), .BN(D5139_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5116 ( .Y(D5116_Y), .A(D5098_Y), .BN(D520_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5115 ( .Y(D5115_Y), .A(D6504_Y), .BN(D5135_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5114 ( .Y(D5114_Y), .A(D7908_Y), .BN(D518_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5113 ( .Y(D5113_Y), .A(D6501_Y), .BN(D5133_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5112 ( .Y(D5112_Y), .A(D6498_Y), .BN(D5134_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5111 ( .Y(D5111_Y), .A(D6504_Y), .BN(D5136_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5110 ( .Y(D5110_Y), .A(D6503_Y), .BN(D5130_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5109 ( .Y(D5109_Y), .A(D6502_Y), .BN(D516_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5108 ( .Y(D5108_Y), .A(D6503_Y), .BN(D5124_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5107 ( .Y(D5107_Y), .A(D6499_Y), .BN(D5129_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5106 ( .Y(D5106_Y), .A(D6501_Y), .BN(D5125_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5105 ( .Y(D5105_Y), .A(D6498_Y), .BN(D5132_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5104 ( .Y(D5104_Y), .A(D6281_Y), .BN(D125_Q),     .S0(D8073_Q));
KC_MXI2_X1 D5103 ( .Y(D5103_Y), .A(D1692_Y), .BN(D512_Q),     .S0(D5079_Y));
KC_MXI2_X1 D5102 ( .Y(D5102_Y), .A(D6287_Y), .BN(D5138_Q),     .S0(D8073_Q));
KC_MXI2_X1 D5101 ( .Y(D5101_Y), .A(D6502_Y), .BN(D5123_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5100 ( .Y(D5100_Y), .A(D1692_Y), .BN(D1641_Q),     .S0(D5082_Y));
KC_MXI2_X1 D5099 ( .Y(D5099_Y), .A(D6499_Y), .BN(D5128_Q),     .S0(D5082_Y));
KC_MXI2_X1 D4955 ( .Y(D4955_Y), .A(D4924_Y), .BN(D4940_Y),     .S0(D454_Y));
KC_MXI2_X1 D4719 ( .Y(D4719_Y), .A(D3257_Y), .BN(D4726_Y),     .S0(D390_Y));
KC_MXI2_X1 D4463 ( .Y(D4463_Y), .A(D4297_Y), .BN(D4490_Q),     .S0(D4403_Y));
KC_MXI2_X1 D3622 ( .Y(D3622_Y), .A(D6506_Y), .BN(D3631_Q),     .S0(D5082_Y));
KC_MXI2_X1 D3618 ( .Y(D3618_Y), .A(D5098_Y), .BN(D3630_Q),     .S0(D5082_Y));
KC_MXI2_X1 D3611 ( .Y(D3611_Y), .A(D7910_Y), .BN(D514_Q),     .S0(D5079_Y));
KC_MXI2_X1 D3610 ( .Y(D3610_Y), .A(D7908_Y), .BN(D3628_Q),     .S0(D5082_Y));
KC_MXI2_X1 D3609 ( .Y(D3609_Y), .A(D7909_Y), .BN(D3629_Q),     .S0(D5079_Y));
KC_MXI2_X1 D3607 ( .Y(D3607_Y), .A(D7910_Y), .BN(D123_Q),     .S0(D5082_Y));
KC_MXI2_X1 D3604 ( .Y(D3604_Y), .A(D7909_Y), .BN(D3624_Q),     .S0(D5082_Y));
KC_MXI2_X1 D3355 ( .Y(D3355_Y), .A(D3334_Y), .BN(D4797_Y),     .S0(D4796_Y));
KC_MXI2_X1 D3264 ( .Y(D3264_Y), .A(D1574_Y), .BN(D3224_Y),     .S0(D3222_Y));
KC_MXI2_X1 D2055 ( .Y(D2055_Y), .A(D8699_Y), .BN(D8807_Y),     .S0(D2057_S));
KC_MXI2_X1 D1761 ( .Y(D1761_Y), .A(D4747_Y), .BN(D6475_Q),     .S0(D8073_Q));
KC_MXI2_X1 D1621 ( .Y(D1621_Y), .A(D6507_Y), .BN(D124_Q),     .S0(D5079_Y));
KC_MXI2_X1 D1463 ( .Y(D1463_Y), .A(D6505_Y), .BN(D3632_Q),     .S0(D5082_Y));
KC_MXI2_X1 D101 ( .Y(D101_Y), .A(D4747_Y), .BN(D6552_Q), .S0(D8073_Q));
KC_AND2_X1 D16514 ( .B(D16540_Y), .A(D16539_Y), .Y(D16514_Y));
KC_AND2_X1 D16468 ( .B(D16382_Y), .A(D16428_Y), .Y(D16468_Y));
KC_AND2_X1 D16131 ( .B(D15315_Y), .A(D16188_Y), .Y(D16131_Y));
KC_AND2_X1 D15327 ( .B(D15283_Y), .A(D15282_Y), .Y(D15327_Y));
KC_AND2_X1 D15326 ( .B(D15280_Y), .A(D15262_Y), .Y(D15326_Y));
KC_AND2_X1 D15320 ( .B(D16089_Y), .A(D15262_Y), .Y(D15320_Y));
KC_AND2_X1 D14676 ( .B(D14653_Y), .A(D13973_Y), .Y(D14676_Y));
KC_AND2_X1 D14673 ( .B(D14531_Y), .A(D15504_Y), .Y(D14673_Y));
KC_AND2_X1 D14576 ( .B(D14518_Q), .A(D14544_Y), .Y(D14576_Y));
KC_AND2_X1 D14488 ( .B(D14481_Y), .A(D13804_Q), .Y(D14488_Y));
KC_AND2_X1 D14468 ( .B(D14455_Y), .A(D13807_Q), .Y(D14468_Y));
KC_AND2_X1 D14467 ( .B(D13774_Y), .A(D13811_Q), .Y(D14467_Y));
KC_AND2_X1 D14465 ( .B(D13779_Y), .A(D13809_Q), .Y(D14465_Y));
KC_AND2_X1 D14372 ( .B(D13717_Y), .A(D13760_Q), .Y(D14372_Y));
KC_AND2_X1 D14371 ( .B(D13729_Y), .A(D13764_Q), .Y(D14371_Y));
KC_AND2_X1 D14079 ( .B(D13236_Y), .A(D11228_Y), .Y(D14079_Y));
KC_AND2_X1 D14078 ( .B(D13236_Y), .A(D10751_Y), .Y(D14078_Y));
KC_AND2_X1 D14075 ( .B(D13236_Y), .A(D12319_Y), .Y(D14075_Y));
KC_AND2_X1 D14069 ( .B(D13236_Y), .A(D12320_Y), .Y(D14069_Y));
KC_AND2_X1 D13905 ( .B(D13275_Q), .A(D13198_Q), .Y(D13905_Y));
KC_AND2_X1 D13904 ( .B(D13257_Y), .A(D13188_Y), .Y(D13904_Y));
KC_AND2_X1 D13746 ( .B(D13716_Y), .A(D13762_Q), .Y(D13746_Y));
KC_AND2_X1 D13699 ( .B(D13694_S), .A(D12422_Y), .Y(D13699_Y));
KC_AND2_X1 D13697 ( .B(D13693_S), .A(D949_Y), .Y(D13697_Y));
KC_AND2_X1 D13696 ( .B(D13695_S), .A(D950_Y), .Y(D13696_Y));
KC_AND2_X1 D13512 ( .B(D13748_S), .A(D162_Y), .Y(D13512_Y));
KC_AND2_X1 D13386 ( .B(D13236_Y), .A(D10291_Y), .Y(D13386_Y));
KC_AND2_X1 D13384 ( .B(D13236_Y), .A(D10794_Y), .Y(D13384_Y));
KC_AND2_X1 D13383 ( .B(D13346_Y), .A(D13395_Q), .Y(D13383_Y));
KC_AND2_X1 D13379 ( .B(D13328_Y), .A(D13361_Y), .Y(D13379_Y));
KC_AND2_X1 D13378 ( .B(D699_Q), .A(D12732_Y), .Y(D13378_Y));
KC_AND2_X1 D13375 ( .B(D13302_Y), .A(D12279_Q), .Y(D13375_Y));
KC_AND2_X1 D13254 ( .B(D13257_Y), .A(D2454_Y), .Y(D13254_Y));
KC_AND2_X1 D13253 ( .B(D12678_Y), .A(D693_Q), .Y(D13253_Y));
KC_AND2_X1 D13250 ( .B(D13257_Y), .A(D10681_Y), .Y(D13250_Y));
KC_AND2_X1 D13189 ( .B(D13275_Q), .A(D13201_Q), .Y(D13189_Y));
KC_AND2_X1 D13188 ( .B(D2363_Y), .A(D12659_Y), .Y(D13188_Y));
KC_AND2_X1 D13028 ( .B(D2456_S), .A(D12421_Y), .Y(D13028_Y));
KC_AND2_X1 D13027 ( .B(D2457_S), .A(D12420_Y), .Y(D13027_Y));
KC_AND2_X1 D12974 ( .B(D12951_Y), .A(D13566_Y), .Y(D12974_Y));
KC_AND2_X1 D12970 ( .B(D13749_S), .A(D12834_Y), .Y(D12970_Y));
KC_AND2_X1 D12906 ( .B(D14057_Y), .A(D15765_Y), .Y(D12906_Y));
KC_AND2_X1 D12905 ( .B(D12879_Y), .A(D12790_Y), .Y(D12905_Y));
KC_AND2_X1 D12832 ( .B(D14057_Y), .A(D15774_Y), .Y(D12832_Y));
KC_AND2_X1 D12826 ( .B(D12858_Q), .A(D12856_Q), .Y(D12826_Y));
KC_AND2_X1 D12741 ( .B(D13236_Y), .A(D10701_Y), .Y(D12741_Y));
KC_AND2_X1 D12673 ( .B(D13236_Y), .A(D2119_Y), .Y(D12673_Y));
KC_AND2_X1 D12672 ( .B(D13236_Y), .A(D10201_Y), .Y(D12672_Y));
KC_AND2_X1 D12671 ( .B(D13236_Y), .A(D10178_Y), .Y(D12671_Y));
KC_AND2_X1 D12666 ( .B(D13257_Y), .A(D11146_Y), .Y(D12666_Y));
KC_AND2_X1 D12665 ( .B(D13236_Y), .A(D11212_Y), .Y(D12665_Y));
KC_AND2_X1 D12268 ( .B(D12207_Y), .A(D2310_Y), .Y(D12268_Y));
KC_AND2_X1 D12213 ( .B(D10179_Y), .A(D11660_Y), .Y(D12213_Y));
KC_AND2_X1 D11968 ( .B(D11458_Y), .A(D11465_Y), .Y(D11968_Y));
KC_AND2_X1 D11967 ( .B(D11444_Y), .A(D11465_Y), .Y(D11967_Y));
KC_AND2_X1 D11966 ( .B(D1112_Y), .A(D11465_Y), .Y(D11966_Y));
KC_AND2_X1 D11908 ( .B(D10413_Y), .A(D2244_Y), .Y(D11908_Y));
KC_AND2_X1 D11854 ( .B(D11853_Y), .A(D2244_Y), .Y(D11854_Y));
KC_AND2_X1 D11852 ( .B(D11850_Y), .A(D2244_Y), .Y(D11852_Y));
KC_AND2_X1 D11851 ( .B(D889_Y), .A(D2244_Y), .Y(D11851_Y));
KC_AND2_X1 D11849 ( .B(D11843_Y), .A(D2244_Y), .Y(D11849_Y));
KC_AND2_X1 D11848 ( .B(D887_Y), .A(D2244_Y), .Y(D11848_Y));
KC_AND2_X1 D11847 ( .B(D11317_Y), .A(D2244_Y), .Y(D11847_Y));
KC_AND2_X1 D11846 ( .B(D11844_Y), .A(D2244_Y), .Y(D11846_Y));
KC_AND2_X1 D11787 ( .B(D11248_Y), .A(D11257_Y), .Y(D11787_Y));
KC_AND2_X1 D11786 ( .B(D11247_Y), .A(D11257_Y), .Y(D11786_Y));
KC_AND2_X1 D11785 ( .B(D773_Y), .A(D11257_Y), .Y(D11785_Y));
KC_AND2_X1 D11784 ( .B(D11782_Y), .A(D11257_Y), .Y(D11784_Y));
KC_AND2_X1 D11783 ( .B(D11781_Y), .A(D11257_Y), .Y(D11783_Y));
KC_AND2_X1 D11779 ( .B(D2280_Y), .A(D11257_Y), .Y(D11779_Y));
KC_AND2_X1 D11778 ( .B(D11777_Y), .A(D11257_Y), .Y(D11778_Y));
KC_AND2_X1 D11623 ( .B(D12253_Y), .A(D9345_Y), .Y(D11623_Y));
KC_AND2_X1 D11534 ( .B(D11532_Y), .A(D11535_Y), .Y(D11534_Y));
KC_AND2_X1 D11454 ( .B(D11478_Y), .A(D2244_Y), .Y(D11454_Y));
KC_AND2_X1 D11453 ( .B(D11451_Y), .A(D2244_Y), .Y(D11453_Y));
KC_AND2_X1 D11384 ( .B(D8444_Y), .A(D11386_Y), .Y(D11384_Y));
KC_AND2_X1 D11383 ( .B(D8447_Y), .A(D11386_Y), .Y(D11383_Y));
KC_AND2_X1 D11382 ( .B(D8443_Y), .A(D11386_Y), .Y(D11382_Y));
KC_AND2_X1 D11254 ( .B(D11243_Y), .A(D11257_Y), .Y(D11254_Y));
KC_AND2_X1 D11253 ( .B(D11241_Y), .A(D11257_Y), .Y(D11253_Y));
KC_AND2_X1 D11252 ( .B(D2239_Y), .A(D11257_Y), .Y(D11252_Y));
KC_AND2_X1 D11246 ( .B(D11244_Y), .A(D11257_Y), .Y(D11246_Y));
KC_AND2_X1 D11114 ( .B(D12252_Y), .A(D9345_Y), .Y(D11114_Y));
KC_AND2_X1 D10873 ( .B(D8454_Y), .A(D11256_Y), .Y(D10873_Y));
KC_AND2_X1 D10870 ( .B(D10864_Y), .A(D2223_Y), .Y(D10870_Y));
KC_AND2_X1 D10783 ( .B(D10782_Y), .A(D11257_Y), .Y(D10783_Y));
KC_AND2_X1 D10629 ( .B(D12256_Y), .A(D9345_Y), .Y(D10629_Y));
KC_AND2_X1 D10542 ( .B(D9778_Y), .A(D8532_Y), .Y(D10542_Y));
KC_AND2_X1 D10507 ( .B(D10499_Y), .A(D9781_Y), .Y(D10507_Y));
KC_AND2_X1 D10503 ( .B(D10501_Y), .A(D9781_Y), .Y(D10503_Y));
KC_AND2_X1 D10502 ( .B(D10506_Y), .A(D9781_Y), .Y(D10502_Y));
KC_AND2_X1 D10498 ( .B(D10500_Y), .A(D9781_Y), .Y(D10498_Y));
KC_AND2_X1 D10496 ( .B(D10497_Y), .A(D9781_Y), .Y(D10496_Y));
KC_AND2_X1 D10492 ( .B(D10493_Y), .A(D9781_Y), .Y(D10492_Y));
KC_AND2_X1 D10415 ( .B(D10495_Y), .A(D9781_Y), .Y(D10415_Y));
KC_AND2_X1 D10414 ( .B(D10504_Y), .A(D9781_Y), .Y(D10414_Y));
KC_AND2_X1 D9976 ( .B(D10197_Y), .A(D10095_Y), .Y(D9976_Y));
KC_AND2_X1 D9833 ( .B(D9772_Y), .A(D8532_Y), .Y(D9833_Y));
KC_AND2_X1 D9832 ( .B(D9798_Y), .A(D8532_Y), .Y(D9832_Y));
KC_AND2_X1 D9780 ( .B(D9771_Y), .A(D8532_Y), .Y(D9780_Y));
KC_AND2_X1 D9777 ( .B(D9776_Y), .A(D9781_Y), .Y(D9777_Y));
KC_AND2_X1 D9702 ( .B(D9694_Y), .A(D9781_Y), .Y(D9702_Y));
KC_AND2_X1 D9698 ( .B(D9692_Y), .A(D9781_Y), .Y(D9698_Y));
KC_AND2_X1 D9697 ( .B(D9779_Y), .A(D9781_Y), .Y(D9697_Y));
KC_AND2_X1 D9696 ( .B(D8446_Y), .A(D9781_Y), .Y(D9696_Y));
KC_AND2_X1 D9695 ( .B(D9693_Y), .A(D9781_Y), .Y(D9695_Y));
KC_AND2_X1 D9446 ( .B(D9444_Y), .A(D9381_Y), .Y(D9446_Y));
KC_AND2_X1 D9442 ( .B(D9492_Y), .A(D8105_Y), .Y(D9442_Y));
KC_AND2_X1 D9441 ( .B(D9399_Y), .A(D9550_Y), .Y(D9441_Y));
KC_AND2_X1 D9378 ( .B(D9341_Y), .A(D7782_Y), .Y(D9378_Y));
KC_AND2_X1 D9376 ( .B(D9380_Y), .A(D8056_Y), .Y(D9376_Y));
KC_AND2_X1 D8799 ( .B(D8828_Y), .A(D8842_Y), .Y(D8799_Y));
KC_AND2_X1 D8795 ( .B(D8843_Y), .A(D8830_Y), .Y(D8795_Y));
KC_AND2_X1 D8789 ( .B(D7166_Y), .A(D8773_Y), .Y(D8789_Y));
KC_AND2_X1 D8694 ( .B(D2056_Y), .A(D8728_Y), .Y(D8694_Y));
KC_AND2_X1 D8691 ( .B(D7133_Y), .A(D7132_Y), .Y(D8691_Y));
KC_AND2_X1 D8688 ( .B(D8691_Y), .A(D8691_Y), .Y(D8688_Y));
KC_AND2_X1 D8629 ( .B(D8524_Y), .A(D8532_Y), .Y(D8629_Y));
KC_AND2_X1 D8628 ( .B(D8523_Y), .A(D8532_Y), .Y(D8628_Y));
KC_AND2_X1 D8627 ( .B(D8522_Y), .A(D8532_Y), .Y(D8627_Y));
KC_AND2_X1 D8626 ( .B(D1109_Y), .A(D8532_Y), .Y(D8626_Y));
KC_AND2_X1 D8585 ( .B(D8525_Y), .A(D8532_Y), .Y(D8585_Y));
KC_AND2_X1 D8584 ( .B(D8527_Y), .A(D8532_Y), .Y(D8584_Y));
KC_AND2_X1 D8583 ( .B(D8526_Y), .A(D8532_Y), .Y(D8583_Y));
KC_AND2_X1 D8581 ( .B(D1912_Y), .A(D8532_Y), .Y(D8581_Y));
KC_AND2_X1 D8580 ( .B(D1913_Y), .A(D8532_Y), .Y(D8580_Y));
KC_AND2_X1 D8573 ( .B(D8531_Y), .A(D8532_Y), .Y(D8573_Y));
KC_AND2_X1 D8572 ( .B(D8574_Y), .A(D8532_Y), .Y(D8572_Y));
KC_AND2_X1 D8571 ( .B(D8529_Y), .A(D8532_Y), .Y(D8571_Y));
KC_AND2_X1 D8570 ( .B(D8530_Y), .A(D8532_Y), .Y(D8570_Y));
KC_AND2_X1 D8440 ( .B(D545_Y), .A(D10994_Q), .Y(D8440_Y));
KC_AND2_X1 D8312 ( .B(D8283_Y), .A(D8310_Y), .Y(D8312_Y));
KC_AND2_X1 D8038 ( .B(D8042_Y), .A(D8049_Y), .Y(D8038_Y));
KC_AND2_X1 D7963 ( .B(D7941_Y), .A(D7948_Y), .Y(D7963_Y));
KC_AND2_X1 D7702 ( .B(D7735_Q), .A(D7734_Q), .Y(D7702_Y));
KC_AND2_X1 D7578 ( .B(D37_Y), .A(D37_Y), .Y(D7578_Y));
KC_AND2_X1 D7573 ( .B(D7610_Y), .A(D7616_Y), .Y(D7573_Y));
KC_AND2_X1 D7515 ( .B(D6100_Y), .A(D6086_Y), .Y(D7515_Y));
KC_AND2_X1 D7513 ( .B(D7524_QN), .A(D7518_QN), .Y(D7513_Y));
KC_AND2_X1 D7461 ( .B(D5671_Y), .A(D10753_Q), .Y(D7461_Y));
KC_AND2_X1 D7131 ( .B(D7158_Y), .A(D7156_Y), .Y(D7131_Y));
KC_AND2_X1 D7003 ( .B(D6949_Y), .A(D6958_Y), .Y(D7003_Y));
KC_AND2_X1 D7002 ( .B(D8575_Y), .A(D6958_Y), .Y(D7002_Y));
KC_AND2_X1 D6957 ( .B(D1757_Y), .A(D6958_Y), .Y(D6957_Y));
KC_AND2_X1 D6956 ( .B(D6886_Y), .A(D6958_Y), .Y(D6956_Y));
KC_AND2_X1 D6952 ( .B(D1756_Y), .A(D6958_Y), .Y(D6952_Y));
KC_AND2_X1 D6891 ( .B(D8445_Y), .A(D5391_Y), .Y(D6891_Y));
KC_AND2_X1 D6890 ( .B(D6856_Y), .A(D5391_Y), .Y(D6890_Y));
KC_AND2_X1 D6888 ( .B(D781_Y), .A(D781_Y), .Y(D6888_Y));
KC_AND2_X1 D6805 ( .B(D6803_Y), .A(D8049_Y), .Y(D6805_Y));
KC_AND2_X1 D6797 ( .B(D6796_Y), .A(D5391_Y), .Y(D6797_Y));
KC_AND2_X1 D6742 ( .B(D6732_Y), .A(D8049_Y), .Y(D6742_Y));
KC_AND2_X1 D6731 ( .B(D6727_Y), .A(D8049_Y), .Y(D6731_Y));
KC_AND2_X1 D6649 ( .B(D6648_Y), .A(D8049_Y), .Y(D6649_Y));
KC_AND2_X1 D6645 ( .B(D6642_Y), .A(D8049_Y), .Y(D6645_Y));
KC_AND2_X1 D6320 ( .B(D6301_Y), .A(D6319_Y), .Y(D6320_Y));
KC_AND2_X1 D6247 ( .B(D6254_Y), .A(D6238_Y), .Y(D6247_Y));
KC_AND2_X1 D6167 ( .B(D6160_Y), .A(D6205_Y), .Y(D6167_Y));
KC_AND2_X1 D6109 ( .B(D6102_Y), .A(D6084_Y), .Y(D6109_Y));
KC_AND2_X1 D6066 ( .B(D6042_Y), .A(D6064_Y), .Y(D6066_Y));
KC_AND2_X1 D5556 ( .B(D6950_Y), .A(D6958_Y), .Y(D5556_Y));
KC_AND2_X1 D5555 ( .B(D6955_Y), .A(D6958_Y), .Y(D5555_Y));
KC_AND2_X1 D5458 ( .B(D8303_Y), .A(D5390_Y), .Y(D5458_Y));
KC_AND2_X1 D5457 ( .B(D8452_Y), .A(D5390_Y), .Y(D5457_Y));
KC_AND2_X1 D5456 ( .B(D8451_Y), .A(D5390_Y), .Y(D5456_Y));
KC_AND2_X1 D5455 ( .B(D8450_Y), .A(D5390_Y), .Y(D5455_Y));
KC_AND2_X1 D5386 ( .B(D6799_Y), .A(D5390_Y), .Y(D5386_Y));
KC_AND2_X1 D5385 ( .B(D5404_Y), .A(D5481_Y), .Y(D5385_Y));
KC_AND2_X1 D5382 ( .B(D6806_Y), .A(D5390_Y), .Y(D5382_Y));
KC_AND2_X1 D5381 ( .B(D6807_Y), .A(D5390_Y), .Y(D5381_Y));
KC_AND2_X1 D5380 ( .B(D8307_Y), .A(D5390_Y), .Y(D5380_Y));
KC_AND2_X1 D5379 ( .B(D8311_Y), .A(D5390_Y), .Y(D5379_Y));
KC_AND2_X1 D5300 ( .B(D6738_Y), .A(D5390_Y), .Y(D5300_Y));
KC_AND2_X1 D5299 ( .B(D6739_Y), .A(D5390_Y), .Y(D5299_Y));
KC_AND2_X1 D5298 ( .B(D6736_Y), .A(D5390_Y), .Y(D5298_Y));
KC_AND2_X1 D5297 ( .B(D6729_Y), .A(D5390_Y), .Y(D5297_Y));
KC_AND2_X1 D5296 ( .B(D6728_Y), .A(D5390_Y), .Y(D5296_Y));
KC_AND2_X1 D4950 ( .B(D4887_Y), .A(D4871_Y), .Y(D4950_Y));
KC_AND2_X1 D4712 ( .B(D4714_Y), .A(D4664_Y), .Y(D4712_Y));
KC_AND2_X1 D4622 ( .B(D3169_Y), .A(D4608_Y), .Y(D4622_Y));
KC_AND2_X1 D4541 ( .B(D2746_Y), .A(D150_Q), .Y(D4541_Y));
KC_AND2_X1 D4540 ( .B(D2896_Q), .A(D4563_Q), .Y(D4540_Y));
KC_AND2_X1 D4036 ( .B(D4038_Y), .A(D4032_Y), .Y(D4036_Y));
KC_AND2_X1 D4035 ( .B(D4038_Y), .A(D4032_Y), .Y(D4035_Y));
KC_AND2_X1 D3269 ( .B(D3267_Y), .A(D3268_Y), .Y(D3269_Y));
KC_AND2_X1 D3263 ( .B(D3264_Y), .A(D3224_Y), .Y(D3263_Y));
KC_AND2_X1 D3173 ( .B(D3143_Y), .A(D4625_Y), .Y(D3173_Y));
KC_AND2_X1 D3060 ( .B(D2746_Y), .A(D3081_Q), .Y(D3060_Y));
KC_AND2_X1 D3059 ( .B(D2746_Y), .A(D3083_Q), .Y(D3059_Y));
KC_AND2_X1 D3058 ( .B(D2746_Y), .A(D3093_Q), .Y(D3058_Y));
KC_AND2_X1 D3051 ( .B(D3090_Y), .A(D4557_Y), .Y(D3051_Y));
KC_AND2_X1 D3050 ( .B(D3036_Y), .A(D3049_Y), .Y(D3050_Y));
KC_AND2_X1 D3048 ( .B(D3039_Y), .A(D44_Y), .Y(D3048_Y));
KC_AND2_X1 D2983 ( .B(D2998_Y), .A(D2953_Y), .Y(D2983_Y));
KC_AND2_X1 D2981 ( .B(D2941_Y), .A(D2894_Y), .Y(D2981_Y));
KC_AND2_X1 D2980 ( .B(D2945_Y), .A(D2894_Y), .Y(D2980_Y));
KC_AND2_X1 D2977 ( .B(D2940_Y), .A(D2894_Y), .Y(D2977_Y));
KC_AND2_X1 D2868 ( .B(D2853_Y), .A(D2880_Y), .Y(D2868_Y));
KC_AND2_X1 D2509 ( .B(D13257_Y), .A(D13902_Y), .Y(D2509_Y));
KC_AND2_X1 D2508 ( .B(D13257_Y), .A(D2330_Y), .Y(D2508_Y));
KC_AND2_X1 D2507 ( .B(D13275_Q), .A(D13918_Q), .Y(D2507_Y));
KC_AND2_X1 D2506 ( .B(D13275_Q), .A(D13920_Q), .Y(D2506_Y));
KC_AND2_X1 D2505 ( .B(D13275_Q), .A(D13860_Q), .Y(D2505_Y));
KC_AND2_X1 D2504 ( .B(D13275_Q), .A(D619_Q), .Y(D2504_Y));
KC_AND2_X1 D2462 ( .B(D13257_Y), .A(D13218_Y), .Y(D2462_Y));
KC_AND2_X1 D2461 ( .B(D13257_Y), .A(D13229_Y), .Y(D2461_Y));
KC_AND2_X1 D2459 ( .B(D13275_Q), .A(D607_Q), .Y(D2459_Y));
KC_AND2_X1 D2283 ( .B(D2281_Y), .A(D11257_Y), .Y(D2283_Y));
KC_AND2_X1 D1918 ( .B(D7736_Q), .A(D7745_Q), .Y(D1918_Y));
KC_AND2_X1 D1766 ( .B(D1764_Y), .A(D6245_Y), .Y(D1766_Y));
KC_AND2_X1 D1760 ( .B(D1916_Y), .A(D8049_Y), .Y(D1760_Y));
KC_AND2_X1 D1759 ( .B(D6802_Y), .A(D8049_Y), .Y(D1759_Y));
KC_AND2_X1 D1626 ( .B(D2746_Y), .A(D727_Y), .Y(D1626_Y));
KC_AND2_X1 D1619 ( .B(D8308_Y), .A(D5390_Y), .Y(D1619_Y));
KC_AND2_X1 D1618 ( .B(D882_Y), .A(D5390_Y), .Y(D1618_Y));
KC_AND2_X1 D19 ( .B(D2746_Y), .A(D3077_Q), .Y(D19_Y));
KC_AND2_X1 D1470 ( .B(D2746_Y), .A(D3082_Q), .Y(D1470_Y));
KC_AND2_X1 D1113 ( .B(D9775_Y), .A(D9781_Y), .Y(D1113_Y));
KC_AND2_X1 D1007 ( .B(D9773_Y), .A(D9781_Y), .Y(D1007_Y));
KC_AND2_X1 D1004 ( .B(D11456_Y), .A(D11386_Y), .Y(D1004_Y));
KC_AND2_X1 D1003 ( .B(D8442_Y), .A(D9781_Y), .Y(D1003_Y));
KC_AND2_X1 D1002 ( .B(D1001_Y), .A(D5391_Y), .Y(D1002_Y));
KC_AND2_X1 D585 ( .B(D11648_Y), .A(D11653_Y), .Y(D585_Y));
KC_AND2_X1 D580 ( .B(D8035_Y), .A(D8049_Y), .Y(D580_Y));
KC_AND2_X1 D579 ( .B(D8039_Y), .A(D8049_Y), .Y(D579_Y));
KC_AND2_X1 D577 ( .B(D578_Y), .A(D8049_Y), .Y(D577_Y));
KC_AND2_X1 D576 ( .B(D6593_Y), .A(D8049_Y), .Y(D576_Y));
KC_AND2_X1 D317 ( .B(D2746_Y), .A(D325_Q), .Y(D317_Y));
KC_AND2_X1 D188 ( .B(D9928_Y), .A(D9986_Y), .Y(D188_Y));
KC_AND2_X1 D186 ( .B(D6334_Y), .A(D7256_Y), .Y(D186_Y));
KC_AND2_X1 D100 ( .B(D8134_Y), .A(D8049_Y), .Y(D100_Y));
KC_OAI21_X2 D16596 ( .B0(D16590_Q), .B1(D16563_Y), .A(D16600_Y),     .Y(D16596_Y));
KC_OAI21_X2 D16137 ( .B0(D15267_Y), .B1(D2654_Y), .A(D16087_Y),     .Y(D16137_Y));
KC_OAI21_X2 D16136 ( .B0(D16110_Y), .B1(D16122_Y), .A(D16037_Y),     .Y(D16136_Y));
KC_OAI21_X2 D16134 ( .B0(D16105_Y), .B1(D16188_Y), .A(D16131_Y),     .Y(D16134_Y));
KC_OAI21_X2 D15941 ( .B0(D15994_Q), .B1(D15961_Y), .A(D15917_Y),     .Y(D15941_Y));
KC_OAI21_X2 D15940 ( .B0(D16010_Q), .B1(D15882_Y), .A(D15912_Y),     .Y(D15940_Y));
KC_OAI21_X2 D15938 ( .B0(D15948_Q), .B1(D15897_Y), .A(D2595_Y),     .Y(D15938_Y));
KC_OAI21_X2 D15933 ( .B0(D16388_Q), .B1(D15883_Y), .A(D15901_Y),     .Y(D15933_Y));
KC_OAI21_X2 D15932 ( .B0(D15947_Q), .B1(D15888_Y), .A(D15893_Y),     .Y(D15932_Y));
KC_OAI21_X2 D15777 ( .B0(D145_Q), .B1(D15728_Y), .A(D15788_Y),     .Y(D15777_Y));
KC_OAI21_X2 D15436 ( .B0(D15408_Y), .B1(D15407_Y), .A(D2629_Y),     .Y(D15436_Y));
KC_OAI21_X2 D15321 ( .B0(D16060_Y), .B1(D15288_Y), .A(D16052_Y),     .Y(D15321_Y));
KC_OAI21_X2 D15125 ( .B0(D15133_Q), .B1(D15094_Y), .A(D15096_Y),     .Y(D15125_Y));
KC_OAI21_X2 D15069 ( .B0(D1158_Q), .B1(D15099_Y), .A(D15014_Y),     .Y(D15069_Y));
KC_OAI21_X2 D14866 ( .B0(D14808_Q), .B1(D815_Q), .A(D14081_Y),     .Y(D14866_Y));
KC_OAI21_X2 D14865 ( .B0(D14790_Q), .B1(D14876_Q), .A(D16765_Y),     .Y(D14865_Y));
KC_OAI21_X2 D14677 ( .B0(D14687_Q), .B1(D14557_Y), .A(D14637_Y),     .Y(D14677_Y));
KC_OAI21_X2 D14672 ( .B0(D636_Y), .B1(D14615_Y), .A(D634_Y),     .Y(D14672_Y));
KC_OAI21_X2 D14582 ( .B0(D14557_Y), .B1(D14556_Y), .A(D14805_Y),     .Y(D14582_Y));
KC_OAI21_X2 D14581 ( .B0(D14520_Q), .B1(D14557_Y), .A(D14560_Y),     .Y(D14581_Y));
KC_OAI21_X2 D14577 ( .B0(D14542_Y), .B1(D14557_Y), .A(D14805_Y),     .Y(D14577_Y));
KC_OAI21_X2 D14507 ( .B0(D14502_Y), .B1(D14500_Y), .A(D14497_Y),     .Y(D14507_Y));
KC_OAI21_X2 D14230 ( .B0(D14305_Q), .B1(D2419_Y), .A(D14084_Y),     .Y(D14230_Y));
KC_OAI21_X2 D14076 ( .B0(D14089_Y), .B1(D14097_Y), .A(D14036_Y),     .Y(D14076_Y));
KC_OAI21_X2 D14074 ( .B0(D13391_Y), .B1(D14097_Y), .A(D758_Y),     .Y(D14074_Y));
KC_OAI21_X2 D14073 ( .B0(D778_Y), .B1(D14097_Y), .A(D14040_Y),     .Y(D14073_Y));
KC_OAI21_X2 D14072 ( .B0(D14084_Y), .B1(D14097_Y), .A(D14032_Y),     .Y(D14072_Y));
KC_OAI21_X2 D14071 ( .B0(D14090_Y), .B1(D14097_Y), .A(D14042_Y),     .Y(D14071_Y));
KC_OAI21_X2 D14070 ( .B0(D14083_Y), .B1(D14097_Y), .A(D14037_Y),     .Y(D14070_Y));
KC_OAI21_X2 D14068 ( .B0(D13987_Y), .B1(D14097_Y), .A(D14035_Y),     .Y(D14068_Y));
KC_OAI21_X2 D14067 ( .B0(D14082_Y), .B1(D14097_Y), .A(D14096_Y),     .Y(D14067_Y));
KC_OAI21_X2 D13514 ( .B0(D13471_Y), .B1(D13477_Y), .A(D13476_Y),     .Y(D13514_Y));
KC_OAI21_X2 D13510 ( .B0(D13434_Y), .B1(D13446_Y), .A(D13445_Y),     .Y(D13510_Y));
KC_OAI21_X2 D13385 ( .B0(D7305_Y), .B1(D13380_Y), .A(D13323_Y),     .Y(D13385_Y));
KC_OAI21_X2 D13380 ( .B0(D13338_Y), .B1(D12892_Y), .A(D13393_Y),     .Y(D13380_Y));
KC_OAI21_X2 D13255 ( .B0(D15508_Y), .B1(D13372_Y), .A(D12731_Y),     .Y(D13255_Y));
KC_OAI21_X2 D13187 ( .B0(D2409_Y), .B1(D12195_Y), .A(D13257_Y),     .Y(D13187_Y));
KC_OAI21_X2 D13029 ( .B0(D2397_Y), .B1(D13010_Y), .A(D12947_Y),     .Y(D13029_Y));
KC_OAI21_X2 D12973 ( .B0(D814_Q), .B1(D13709_Y), .A(D12949_Y),     .Y(D12973_Y));
KC_OAI21_X2 D12972 ( .B0(D13452_Y), .B1(D13010_Y), .A(D12947_Y),     .Y(D12972_Y));
KC_OAI21_X2 D12971 ( .B0(D12988_Y), .B1(D12943_Y), .A(D12951_Y),     .Y(D12971_Y));
KC_OAI21_X2 D12969 ( .B0(D12942_Y), .B1(D13010_Y), .A(D12947_Y),     .Y(D12969_Y));
KC_OAI21_X2 D12968 ( .B0(D12941_Y), .B1(D13010_Y), .A(D12947_Y),     .Y(D12968_Y));
KC_OAI21_X2 D12967 ( .B0(D2398_Y), .B1(D13010_Y), .A(D12947_Y),     .Y(D12967_Y));
KC_OAI21_X2 D12907 ( .B0(D12857_Q), .B1(D12785_Y), .A(D12777_Y),     .Y(D12907_Y));
KC_OAI21_X2 D12902 ( .B0(D12749_Q), .B1(D12785_Y), .A(D12777_Y),     .Y(D12902_Y));
KC_OAI21_X2 D12836 ( .B0(D13330_Y), .B1(D12795_Y), .A(D14057_Y),     .Y(D12836_Y));
KC_OAI21_X2 D12835 ( .B0(D13330_Y), .B1(D12810_Y), .A(D14057_Y),     .Y(D12835_Y));
KC_OAI21_X2 D12833 ( .B0(D13330_Y), .B1(D14730_Y), .A(D14057_Y),     .Y(D12833_Y));
KC_OAI21_X2 D12830 ( .B0(D843_Q), .B1(D12785_Y), .A(D12777_Y),     .Y(D12830_Y));
KC_OAI21_X2 D12824 ( .B0(D13330_Y), .B1(D15498_Y), .A(D14057_Y),     .Y(D12824_Y));
KC_OAI21_X2 D12738 ( .B0(D12739_Y), .B1(D12717_Y), .A(D12255_Y),     .Y(D12738_Y));
KC_OAI21_X2 D12737 ( .B0(D12755_Q), .B1(D12357_Q), .A(D12707_Y),     .Y(D12737_Y));
KC_OAI21_X2 D12736 ( .B0(D12813_Y), .B1(D12704_Y), .A(D12296_Y),     .Y(D12736_Y));
KC_OAI21_X2 D12735 ( .B0(D819_Q), .B1(D13363_Y), .A(D13228_Y),     .Y(D12735_Y));
KC_OAI21_X2 D12667 ( .B0(D2362_Y), .B1(D12195_Y), .A(D13257_Y),     .Y(D12667_Y));
KC_OAI21_X2 D12625 ( .B0(D12631_Y), .B1(D13287_Y), .A(D12623_Y),     .Y(D12625_Y));
KC_OAI21_X2 D12335 ( .B0(D12854_Q), .B1(D821_Q), .A(D12245_Y),     .Y(D12335_Y));
KC_OAI21_X2 D12334 ( .B0(D12857_Q), .B1(D823_Q), .A(D12247_Y),     .Y(D12334_Y));
KC_OAI21_X2 D12266 ( .B0(D716_Q), .B1(D12275_Q), .A(D12245_Y),     .Y(D12266_Y));
KC_OAI21_X2 D12265 ( .B0(D12657_Y), .B1(D12276_Y), .A(D12725_Y),     .Y(D12265_Y));
KC_OAI21_X2 D12264 ( .B0(D12752_Q), .B1(D12360_Q), .A(D12247_Y),     .Y(D12264_Y));
KC_OAI21_X2 D12212 ( .B0(D10177_Y), .B1(D12192_Y), .A(D12213_Y),     .Y(D12212_Y));
KC_OAI21_X2 D11907 ( .B0(D980_Y), .B1(D11377_Y), .A(D11386_Y),     .Y(D11907_Y));
KC_OAI21_X2 D11906 ( .B0(D981_Y), .B1(D11377_Y), .A(D2244_Y),     .Y(D11906_Y));
KC_OAI21_X2 D11905 ( .B0(D11365_Y), .B1(D980_Y), .A(D11386_Y),     .Y(D11905_Y));
KC_OAI21_X2 D11594 ( .B0(D11552_Y), .B1(D11591_Y), .A(D11536_Y),     .Y(D11594_Y));
KC_OAI21_X2 D11575 ( .B0(D11553_Y), .B1(D11563_Y), .A(D11535_Y),     .Y(D11575_Y));
KC_OAI21_X2 D11574 ( .B0(D11550_Y), .B1(D11563_Y), .A(D11535_Y),     .Y(D11574_Y));
KC_OAI21_X2 D11573 ( .B0(D11554_Y), .B1(D11553_Y), .A(D11535_Y),     .Y(D11573_Y));
KC_OAI21_X2 D11572 ( .B0(D11553_Y), .B1(D11564_Y), .A(D11535_Y),     .Y(D11572_Y));
KC_OAI21_X2 D11571 ( .B0(D11549_Y), .B1(D11553_Y), .A(D11535_Y),     .Y(D11571_Y));
KC_OAI21_X2 D11570 ( .B0(D11549_Y), .B1(D11550_Y), .A(D11535_Y),     .Y(D11570_Y));
KC_OAI21_X2 D11569 ( .B0(D11550_Y), .B1(D11564_Y), .A(D11535_Y),     .Y(D11569_Y));
KC_OAI21_X2 D11568 ( .B0(D11554_Y), .B1(D11550_Y), .A(D11535_Y),     .Y(D11568_Y));
KC_OAI21_X2 D11385 ( .B0(D11358_Y), .B1(D981_Y), .A(D11386_Y),     .Y(D11385_Y));
KC_OAI21_X2 D11381 ( .B0(D981_Y), .B1(D11379_Y), .A(D11386_Y),     .Y(D11381_Y));
KC_OAI21_X2 D11380 ( .B0(D980_Y), .B1(D11379_Y), .A(D11386_Y),     .Y(D11380_Y));
KC_OAI21_X2 D11321 ( .B0(D10852_Y), .B1(D11305_Y), .A(D11256_Y),     .Y(D11321_Y));
KC_OAI21_X2 D11162 ( .B0(D11152_Y), .B1(D11153_Y), .A(D11258_Y),     .Y(D11162_Y));
KC_OAI21_X2 D11161 ( .B0(D11152_Y), .B1(D11154_Y), .A(D11258_Y),     .Y(D11161_Y));
KC_OAI21_X2 D11160 ( .B0(D11143_Y), .B1(D11152_Y), .A(D11258_Y),     .Y(D11160_Y));
KC_OAI21_X2 D11159 ( .B0(D11144_Y), .B1(D11152_Y), .A(D11258_Y),     .Y(D11159_Y));
KC_OAI21_X2 D11158 ( .B0(D11143_Y), .B1(D11148_Y), .A(D11258_Y),     .Y(D11158_Y));
KC_OAI21_X2 D11157 ( .B0(D11144_Y), .B1(D11148_Y), .A(D11258_Y),     .Y(D11157_Y));
KC_OAI21_X2 D11156 ( .B0(D11148_Y), .B1(D11154_Y), .A(D11258_Y),     .Y(D11156_Y));
KC_OAI21_X2 D11155 ( .B0(D11148_Y), .B1(D11153_Y), .A(D11258_Y),     .Y(D11155_Y));
KC_OAI21_X2 D11099 ( .B0(D11548_Y), .B1(D11566_Y), .A(D11536_Y),     .Y(D11099_Y));
KC_OAI21_X2 D11065 ( .B0(D11552_Y), .B1(D11548_Y), .A(D11536_Y),     .Y(D11065_Y));
KC_OAI21_X2 D11064 ( .B0(D11548_Y), .B1(D11565_Y), .A(D11536_Y),     .Y(D11064_Y));
KC_OAI21_X2 D10874 ( .B0(D10855_Y), .B1(D10846_Y), .A(D11256_Y),     .Y(D10874_Y));
KC_OAI21_X2 D10872 ( .B0(D10852_Y), .B1(D10862_Y), .A(D11256_Y),     .Y(D10872_Y));
KC_OAI21_X2 D10868 ( .B0(D10846_Y), .B1(D10862_Y), .A(D11256_Y),     .Y(D10868_Y));
KC_OAI21_X2 D10867 ( .B0(D10847_Y), .B1(D10852_Y), .A(D11256_Y),     .Y(D10867_Y));
KC_OAI21_X2 D10866 ( .B0(D10847_Y), .B1(D10846_Y), .A(D11256_Y),     .Y(D10866_Y));
KC_OAI21_X2 D10865 ( .B0(D10855_Y), .B1(D10852_Y), .A(D11256_Y),     .Y(D10865_Y));
KC_OAI21_X2 D10139 ( .B0(D417_Y), .B1(D10161_Y), .A(D7683_Y),     .Y(D10139_Y));
KC_OAI21_X2 D10138 ( .B0(D417_Y), .B1(D10162_Y), .A(D7683_Y),     .Y(D10138_Y));
KC_OAI21_X2 D10056 ( .B0(D10065_Y), .B1(D2122_Y), .A(D10055_Y),     .Y(D10056_Y));
KC_OAI21_X2 D9931 ( .B0(D9946_Y), .B1(D9946_Y), .A(D9927_Y),     .Y(D9931_Y));
KC_OAI21_X2 D9932 ( .B0(D9927_Y), .B1(D9926_Y), .A(D8697_Y),     .Y(D9932_Y));
KC_OAI21_X2 D9560 ( .B0(D9523_Y), .B1(D622_Y), .A(D9389_Y),     .Y(D9560_Y));
KC_OAI21_X2 D9557 ( .B0(D9511_Y), .B1(D9521_Y), .A(D9508_Y),     .Y(D9557_Y));
KC_OAI21_X2 D9445 ( .B0(D1994_Y), .B1(D9407_Y), .A(D1982_Y),     .Y(D9445_Y));
KC_OAI21_X2 D9444 ( .B0(D9400_Y), .B1(D8079_Y), .A(D9473_Y),     .Y(D9444_Y));
KC_OAI21_X2 D9317 ( .B0(D417_Y), .B1(D10159_Y), .A(D9167_Y),     .Y(D9317_Y));
KC_OAI21_X2 D9316 ( .B0(D417_Y), .B1(D7730_Y), .A(D2002_Y),     .Y(D9316_Y));
KC_OAI21_X2 D9314 ( .B0(D417_Y), .B1(D10157_Y), .A(D9167_Y),     .Y(D9314_Y));
KC_OAI21_X2 D9313 ( .B0(D417_Y), .B1(D9354_Y), .A(D434_Y),     .Y(D9313_Y));
KC_OAI21_X2 D9312 ( .B0(D417_Y), .B1(D9266_Y), .A(D9240_Y),     .Y(D9312_Y));
KC_OAI21_X2 D9311 ( .B0(D417_Y), .B1(D481_Y), .A(D434_Y), .Y(D9311_Y));
KC_OAI21_X2 D9310 ( .B0(D417_Y), .B1(D7784_Y), .A(D9240_Y),     .Y(D9310_Y));
KC_OAI21_X2 D9256 ( .B0(D417_Y), .B1(D7785_Y), .A(D9101_Y),     .Y(D9256_Y));
KC_OAI21_X2 D9253 ( .B0(D417_Y), .B1(D7713_Y), .A(D2002_Y),     .Y(D9253_Y));
KC_OAI21_X2 D9252 ( .B0(D417_Y), .B1(D10142_Y), .A(D9175_Y),     .Y(D9252_Y));
KC_OAI21_X2 D9251 ( .B0(D417_Y), .B1(D10158_Y), .A(D9180_Y),     .Y(D9251_Y));
KC_OAI21_X2 D9207 ( .B0(D7643_Y), .B1(D9113_Y), .A(D382_Y),     .Y(D9207_Y));
KC_OAI21_X2 D9206 ( .B0(D1711_Y), .B1(D9186_Y), .A(D9147_Y),     .Y(D9206_Y));
KC_OAI21_X2 D9204 ( .B0(D417_Y), .B1(D10160_Y), .A(D9175_Y),     .Y(D9204_Y));
KC_OAI21_X2 D9086 ( .B0(D8072_Y), .B1(D8970_Y), .A(D7510_Y),     .Y(D9086_Y));
KC_OAI21_X2 D9001 ( .B0(D2065_Y), .B1(D8993_Y), .A(D7430_Y),     .Y(D9001_Y));
KC_OAI21_X2 D8996 ( .B0(D9019_Q), .B1(D8970_Y), .A(D7447_Y),     .Y(D8996_Y));
KC_OAI21_X2 D8801 ( .B0(D204_Y), .B1(D8742_Y), .A(D211_Y),     .Y(D8801_Y));
KC_OAI21_X2 D8792 ( .B0(D2029_Y), .B1(D2028_Y), .A(D8797_Y),     .Y(D8792_Y));
KC_OAI21_X2 D8309 ( .B0(D1993_Y), .B1(D8297_Y), .A(D8029_Y),     .Y(D8309_Y));
KC_OAI21_X2 D8302 ( .B0(D9369_Y), .B1(D8297_Y), .A(D8029_Y),     .Y(D8302_Y));
KC_OAI21_X2 D8223 ( .B0(D8219_Y), .B1(D9545_Y), .A(D8256_Y),     .Y(D8223_Y));
KC_OAI21_X2 D8139 ( .B0(D8835_Q), .B1(D8242_Y), .A(D8099_Y),     .Y(D8139_Y));
KC_OAI21_X2 D8137 ( .B0(D8248_Q), .B1(D8120_Y), .A(D704_Q),     .Y(D8137_Y));
KC_OAI21_X2 D8136 ( .B0(D4137_Q), .B1(D9437_Y), .A(D8120_Y),     .Y(D8136_Y));
KC_OAI21_X2 D8135 ( .B0(D8836_Q), .B1(D8242_Y), .A(D8099_Y),     .Y(D8135_Y));
KC_OAI21_X2 D8130 ( .B0(D1989_Y), .B1(D9518_Y), .A(D8079_Y),     .Y(D8130_Y));
KC_OAI21_X2 D8044 ( .B0(D609_Q), .B1(D581_Y), .A(D8015_Y),     .Y(D8044_Y));
KC_OAI21_X2 D8031 ( .B0(D8002_Y), .B1(D9365_Y), .A(D8029_Y),     .Y(D8031_Y));
KC_OAI21_X2 D7961 ( .B0(D7943_Y), .B1(D7919_Y), .A(D7888_Q),     .Y(D7961_Y));
KC_OAI21_X2 D7879 ( .B0(D7872_Y), .B1(D7848_Y), .A(D7945_Y),     .Y(D7879_Y));
KC_OAI21_X2 D7878 ( .B0(D6441_Y), .B1(D7858_Y), .A(D7852_Y),     .Y(D7878_Y));
KC_OAI21_X2 D7876 ( .B0(D7848_Y), .B1(D7881_Y), .A(D1856_Y),     .Y(D7876_Y));
KC_OAI21_X2 D7874 ( .B0(D1859_Y), .B1(D7888_Q), .A(D7835_Y),     .Y(D7874_Y));
KC_OAI21_X2 D7873 ( .B0(D7839_Y), .B1(D7829_Y), .A(D7836_Y),     .Y(D7873_Y));
KC_OAI21_X2 D7711 ( .B0(D9021_Q), .B1(D2099_Y), .A(D7744_Y),     .Y(D7711_Y));
KC_OAI21_X2 D7707 ( .B0(D8953_Q), .B1(D2099_Y), .A(D7743_Y),     .Y(D7707_Y));
KC_OAI21_X2 D7705 ( .B0(D7713_Y), .B1(D6350_Q), .A(D7718_Y),     .Y(D7705_Y));
KC_OAI21_X2 D7703 ( .B0(D6328_Y), .B1(D7740_Y), .A(D404_Y),     .Y(D7703_Y));
KC_OAI21_X2 D7576 ( .B0(D7613_Y), .B1(D8970_Y), .A(D7447_Y),     .Y(D7576_Y));
KC_OAI21_X2 D7458 ( .B0(D6046_Y), .B1(D7517_Y), .A(D5936_Y),     .Y(D7458_Y));
KC_OAI21_X2 D7385 ( .B0(D5857_Y), .B1(D7323_Y), .A(D7204_Y),     .Y(D7385_Y));
KC_OAI21_X2 D7383 ( .B0(D7393_Y), .B1(D7342_Y), .A(D7317_Y),     .Y(D7383_Y));
KC_OAI21_X2 D7289 ( .B0(D7264_Y), .B1(D7265_Y), .A(D7249_Y),     .Y(D7289_Y));
KC_OAI21_X2 D7286 ( .B0(D7224_Y), .B1(D7208_Y), .A(D7249_Y),     .Y(D7286_Y));
KC_OAI21_X2 D7284 ( .B0(D7441_Y), .B1(D7236_Y), .A(D7202_Y),     .Y(D7284_Y));
KC_OAI21_X2 D7283 ( .B0(D7634_Y), .B1(D7205_Y), .A(D7222_Y),     .Y(D7283_Y));
KC_OAI21_X2 D7282 ( .B0(D7186_Y), .B1(D209_Y), .A(D7180_Y),     .Y(D7282_Y));
KC_OAI21_X2 D7281 ( .B0(D209_Y), .B1(D7204_Y), .A(D210_Y),     .Y(D7281_Y));
KC_OAI21_X2 D7280 ( .B0(D7209_Y), .B1(D8756_Y), .A(D7178_Y),     .Y(D7280_Y));
KC_OAI21_X2 D7129 ( .B0(D5658_Y), .B1(D5880_Y), .A(D7148_Q),     .Y(D7129_Y));
KC_OAI21_X2 D7128 ( .B0(D7124_Y), .B1(D5658_Y), .A(D7129_Y),     .Y(D7128_Y));
KC_OAI21_X2 D6537 ( .B0(D6553_Q), .B1(D6512_Y), .A(D6517_Y),     .Y(D6537_Y));
KC_OAI21_X2 D6459 ( .B0(D5031_Y), .B1(D1564_Y), .A(D6416_Y),     .Y(D6459_Y));
KC_OAI21_X2 D6318 ( .B0(D6319_Y), .B1(D6176_Y), .A(D6320_Y),     .Y(D6318_Y));
KC_OAI21_X2 D6070 ( .B0(D6038_Y), .B1(D6047_Y), .A(D7337_Y),     .Y(D6070_Y));
KC_OAI21_X2 D6069 ( .B0(D6006_Y), .B1(D1627_Y), .A(D5988_Y),     .Y(D6069_Y));
KC_OAI21_X2 D6067 ( .B0(D6000_Y), .B1(D5984_Y), .A(D5988_Y),     .Y(D6067_Y));
KC_OAI21_X2 D6063 ( .B0(D165_Y), .B1(D4405_Y), .A(D5956_Y),     .Y(D6063_Y));
KC_OAI21_X2 D6062 ( .B0(D4417_Y), .B1(D4412_Y), .A(D275_Y),     .Y(D6062_Y));
KC_OAI21_X2 D5928 ( .B0(D4340_Y), .B1(D5918_Y), .A(D7242_Y),     .Y(D5928_Y));
KC_OAI21_X2 D5927 ( .B0(D7232_Y), .B1(D5838_Y), .A(D177_Y),     .Y(D5927_Y));
KC_OAI21_X2 D5926 ( .B0(D4368_Y), .B1(D4326_Y), .A(D5870_Y),     .Y(D5926_Y));
KC_OAI21_X2 D5923 ( .B0(D5835_Y), .B1(D5905_Y), .A(D5851_Y),     .Y(D5923_Y));
KC_OAI21_X2 D5922 ( .B0(D243_Y), .B1(D10050_Y), .A(D6001_Y),     .Y(D5922_Y));
KC_OAI21_X2 D5921 ( .B0(D6073_Q), .B1(D5866_Y), .A(D5905_Y),     .Y(D5921_Y));
KC_OAI21_X2 D5920 ( .B0(D6071_Y), .B1(D254_Y), .A(D7461_Y),     .Y(D5920_Y));
KC_OAI21_X2 D5798 ( .B0(D6072_Y), .B1(D94_Y), .A(D5886_Y),     .Y(D5798_Y));
KC_OAI21_X2 D5797 ( .B0(D1754_Y), .B1(D218_Y), .A(D5804_Y),     .Y(D5797_Y));
KC_OAI21_X2 D5795 ( .B0(D8788_Y), .B1(D5769_Y), .A(D4193_Y),     .Y(D5795_Y));
KC_OAI21_X2 D5794 ( .B0(D5722_Y), .B1(D217_Y), .A(D5775_Y),     .Y(D5794_Y));
KC_OAI21_X2 D5182 ( .B0(D1411_Y), .B1(D3716_Y), .A(D5215_Y),     .Y(D5182_Y));
KC_OAI21_X2 D5181 ( .B0(D1413_Y), .B1(D3716_Y), .A(D5215_Y),     .Y(D5181_Y));
KC_OAI21_X2 D5071 ( .B0(D1565_Y), .B1(D3413_Y), .A(D4985_Y),     .Y(D5071_Y));
KC_OAI21_X2 D5070 ( .B0(D4868_Y), .B1(D5021_Y), .A(D3484_Q),     .Y(D5070_Y));
KC_OAI21_X2 D5069 ( .B0(D3067_Y), .B1(D3371_Y), .A(D4999_Y),     .Y(D5069_Y));
KC_OAI21_X2 D4954 ( .B0(D4940_Y), .B1(D4924_Y), .A(D4962_Y),     .Y(D4954_Y));
KC_OAI21_X2 D4953 ( .B0(D1537_Y), .B1(D4925_Y), .A(D4916_Y),     .Y(D4953_Y));
KC_OAI21_X2 D4951 ( .B0(D5009_Y), .B1(D4925_Y), .A(D4903_Y),     .Y(D4951_Y));
KC_OAI21_X2 D4798 ( .B0(D7764_Y), .B1(D7768_Y), .A(D3203_Y),     .Y(D4798_Y));
KC_OAI21_X2 D4796 ( .B0(D3361_Y), .B1(D4780_Y), .A(D4797_Y),     .Y(D4796_Y));
KC_OAI21_X2 D4715 ( .B0(D4690_Y), .B1(D4671_Y), .A(D4703_Y),     .Y(D4715_Y));
KC_OAI21_X2 D4713 ( .B0(D4682_Y), .B1(D4669_Y), .A(D4681_Y),     .Y(D4713_Y));
KC_OAI21_X2 D4625 ( .B0(D4605_Y), .B1(D4595_Y), .A(D4520_Y),     .Y(D4625_Y));
KC_OAI21_X2 D4620 ( .B0(D3114_Y), .B1(D1427_Y), .A(D3243_Y),     .Y(D4620_Y));
KC_OAI21_X2 D4619 ( .B0(D3234_Y), .B1(D3118_Y), .A(D4608_Y),     .Y(D4619_Y));
KC_OAI21_X2 D4542 ( .B0(D7739_Y), .B1(D7316_Y), .A(D7337_Y),     .Y(D4542_Y));
KC_OAI21_X2 D4464 ( .B0(D4304_Y), .B1(D4448_Y), .A(D4476_Y),     .Y(D4464_Y));
KC_OAI21_X2 D4383 ( .B0(D4436_Y), .B1(D4422_Y), .A(D5890_Y),     .Y(D4383_Y));
KC_OAI21_X2 D4382 ( .B0(D1721_Y), .B1(D293_Y), .A(D6058_Y),     .Y(D4382_Y));
KC_OAI21_X2 D4225 ( .B0(D7376_Y), .B1(D5786_Y), .A(D4202_Y),     .Y(D4225_Y));
KC_OAI21_X2 D4224 ( .B0(D4168_Y), .B1(D4187_Y), .A(D4197_Y),     .Y(D4224_Y));
KC_OAI21_X2 D4107 ( .B0(D7376_Y), .B1(D4262_Y), .A(D4098_Y),     .Y(D4107_Y));
KC_OAI21_X2 D4037 ( .B0(D4068_Y), .B1(D4088_Y), .A(D4063_Y),     .Y(D4037_Y));
KC_OAI21_X2 D4006 ( .B0(D3992_Y), .B1(D3987_Y), .A(D5558_Y),     .Y(D4006_Y));
KC_OAI21_X2 D4005 ( .B0(D3986_Y), .B1(D1445_Y), .A(D6958_Y),     .Y(D4005_Y));
KC_OAI21_X2 D4004 ( .B0(D3986_Y), .B1(D1444_Y), .A(D6958_Y),     .Y(D4004_Y));
KC_OAI21_X2 D4003 ( .B0(D3991_Y), .B1(D3986_Y), .A(D6958_Y),     .Y(D4003_Y));
KC_OAI21_X2 D4002 ( .B0(D3987_Y), .B1(D1445_Y), .A(D6958_Y),     .Y(D4002_Y));
KC_OAI21_X2 D4001 ( .B0(D3987_Y), .B1(D1444_Y), .A(D6958_Y),     .Y(D4001_Y));
KC_OAI21_X2 D4000 ( .B0(D3992_Y), .B1(D3986_Y), .A(D6958_Y),     .Y(D4000_Y));
KC_OAI21_X2 D3999 ( .B0(D3991_Y), .B1(D3987_Y), .A(D5558_Y),     .Y(D3999_Y));
KC_OAI21_X2 D3861 ( .B0(D3837_Y), .B1(D3839_Y), .A(D3862_Y),     .Y(D3861_Y));
KC_OAI21_X2 D3859 ( .B0(D1478_Y), .B1(D1504_Y), .A(D3863_Y),     .Y(D3859_Y));
KC_OAI21_X2 D3858 ( .B0(D3838_Y), .B1(D3839_Y), .A(D3862_Y),     .Y(D3858_Y));
KC_OAI21_X2 D3857 ( .B0(D3836_Y), .B1(D3851_Y), .A(D3862_Y),     .Y(D3857_Y));
KC_OAI21_X2 D3856 ( .B0(D3838_Y), .B1(D3836_Y), .A(D3862_Y),     .Y(D3856_Y));
KC_OAI21_X2 D3855 ( .B0(D3839_Y), .B1(D3851_Y), .A(D3862_Y),     .Y(D3855_Y));
KC_OAI21_X2 D3854 ( .B0(D3839_Y), .B1(D3850_Y), .A(D3862_Y),     .Y(D3854_Y));
KC_OAI21_X2 D3853 ( .B0(D3836_Y), .B1(D3850_Y), .A(D3862_Y),     .Y(D3853_Y));
KC_OAI21_X2 D3852 ( .B0(D3837_Y), .B1(D3836_Y), .A(D3862_Y),     .Y(D3852_Y));
KC_OAI21_X2 D3721 ( .B0(D3714_Y), .B1(D1413_Y), .A(D5215_Y),     .Y(D3721_Y));
KC_OAI21_X2 D3720 ( .B0(D3714_Y), .B1(D1411_Y), .A(D5215_Y),     .Y(D3720_Y));
KC_OAI21_X2 D3667 ( .B0(D1412_Y), .B1(D1411_Y), .A(D5215_Y),     .Y(D3667_Y));
KC_OAI21_X2 D3560 ( .B0(D68_Y), .B1(D3416_Y), .A(D5011_Y),     .Y(D3560_Y));
KC_OAI21_X2 D3558 ( .B0(D3528_Y), .B1(D3370_Y), .A(D3544_Y),     .Y(D3558_Y));
KC_OAI21_X2 D3556 ( .B0(D3501_Y), .B1(D3546_Y), .A(D4913_Y),     .Y(D3556_Y));
KC_OAI21_X2 D3475 ( .B0(D3599_Y), .B1(D3304_Y), .A(D3479_Y),     .Y(D3475_Y));
KC_OAI21_X2 D3473 ( .B0(D3372_Q), .B1(D4887_Y), .A(D1415_Y),     .Y(D3473_Y));
KC_OAI21_X2 D3471 ( .B0(D3599_Y), .B1(D3574_Y), .A(D3415_Y),     .Y(D3471_Y));
KC_OAI21_X2 D3470 ( .B0(D3416_Y), .B1(D3365_Y), .A(D3539_Y),     .Y(D3470_Y));
KC_OAI21_X2 D3469 ( .B0(D3437_Y), .B1(D474_Y), .A(D4960_Y),     .Y(D3469_Y));
KC_OAI21_X2 D3354 ( .B0(D4749_Y), .B1(D3340_Y), .A(D1671_Y),     .Y(D3354_Y));
KC_OAI21_X2 D3262 ( .B0(D12305_Y), .B1(D3141_Y), .A(D3248_Y),     .Y(D3262_Y));
KC_OAI21_X2 D3169 ( .B0(D3113_Y), .B1(D3119_Y), .A(D3349_Y),     .Y(D3169_Y));
KC_OAI21_X2 D3167 ( .B0(D4580_Y), .B1(D3116_Y), .A(D3137_Y),     .Y(D3167_Y));
KC_OAI21_X2 D3166 ( .B0(D3193_Y), .B1(D4607_Y), .A(D352_Y),     .Y(D3166_Y));
KC_OAI21_X2 D2979 ( .B0(D2823_Y), .B1(D2946_Y), .A(D2860_Y),     .Y(D2979_Y));
KC_OAI21_X2 D2978 ( .B0(D2823_Y), .B1(D2946_Y), .A(D2824_Y),     .Y(D2978_Y));
KC_OAI21_X2 D2976 ( .B0(D2925_Y), .B1(D2934_Y), .A(D2975_Y),     .Y(D2976_Y));
KC_OAI21_X2 D2975 ( .B0(D2934_Y), .B1(D2819_Y), .A(D2883_Q),     .Y(D2975_Y));
KC_OAI21_X2 D2974 ( .B0(D2929_Y), .B1(D2978_Y), .A(D2971_Y),     .Y(D2974_Y));
KC_OAI21_X2 D2973 ( .B0(D2922_Y), .B1(D1436_Y), .A(D299_Q),     .Y(D2973_Y));
KC_OAI21_X2 D2972 ( .B0(D2921_Y), .B1(D2935_Y), .A(D2970_Y),     .Y(D2972_Y));
KC_OAI21_X2 D2971 ( .B0(D2978_Y), .B1(D1436_Y), .A(D3003_Q),     .Y(D2971_Y));
KC_OAI21_X2 D2970 ( .B0(D2935_Y), .B1(D1436_Y), .A(D3002_Q),     .Y(D2970_Y));
KC_OAI21_X2 D2969 ( .B0(D2926_Y), .B1(D2928_Y), .A(D2968_Y),     .Y(D2969_Y));
KC_OAI21_X2 D2968 ( .B0(D2928_Y), .B1(D1436_Y), .A(D300_Q),     .Y(D2968_Y));
KC_OAI21_X2 D2967 ( .B0(D2819_Y), .B1(D2927_Y), .A(D297_Q),     .Y(D2967_Y));
KC_OAI21_X2 D2966 ( .B0(D2930_Y), .B1(D2819_Y), .A(D4485_Q),     .Y(D2966_Y));
KC_OAI21_X2 D2965 ( .B0(D2914_Y), .B1(D2922_Y), .A(D2973_Y),     .Y(D2965_Y));
KC_OAI21_X2 D2964 ( .B0(D2819_Y), .B1(D2915_Y), .A(D2999_Q),     .Y(D2964_Y));
KC_OAI21_X2 D2963 ( .B0(D2919_Y), .B1(D2920_Y), .A(D2962_Y),     .Y(D2963_Y));
KC_OAI21_X2 D2962 ( .B0(D2920_Y), .B1(D1436_Y), .A(D3001_Q),     .Y(D2962_Y));
KC_OAI21_X2 D2961 ( .B0(D1436_Y), .B1(D2918_Y), .A(D3000_Q),     .Y(D2961_Y));
KC_OAI21_X2 D2960 ( .B0(D1436_Y), .B1(D2917_Y), .A(D298_Q),     .Y(D2960_Y));
KC_OAI21_X2 D2959 ( .B0(D2907_Y), .B1(D2930_Y), .A(D2966_Y),     .Y(D2959_Y));
KC_OAI21_X2 D2958 ( .B0(D2979_Y), .B1(D1436_Y), .A(D4486_Q),     .Y(D2958_Y));
KC_OAI21_X2 D2957 ( .B0(D2906_Y), .B1(D2979_Y), .A(D2958_Y),     .Y(D2957_Y));
KC_OAI21_X2 D1 ( .B0(D2826_Y), .B1(D1459_Y), .A(D1439_Y), .Y(D1_Y));
KC_OAI21_X2 D2865 ( .B0(D2932_Y), .B1(D2939_Y), .A(D1471_Y),     .Y(D2865_Y));
KC_OAI21_X2 D2860 ( .B0(D2887_Q), .B1(D2775_Y), .A(D2857_Y),     .Y(D2860_Y));
KC_OAI21_X2 D2859 ( .B0(D2887_Q), .B1(D2778_Y), .A(D2854_Y),     .Y(D2859_Y));
KC_OAI21_X2 D2787 ( .B0(D2762_Y), .B1(D2768_Y), .A(D2766_Y),     .Y(D2787_Y));
KC_OAI21_X2 D2786 ( .B0(D2759_Y), .B1(D2770_Y), .A(D2769_Y),     .Y(D2786_Y));
KC_OAI21_X2 D2570 ( .B0(D14518_Q), .B1(D14497_Y), .A(D14503_Y),     .Y(D2570_Y));
KC_OAI21_X2 D2569 ( .B0(D749_Y), .B1(D2543_Y), .A(D751_Y),     .Y(D2569_Y));
KC_OAI21_X2 D2566 ( .B0(D2572_Q), .B1(D2529_Y), .A(D15047_Y),     .Y(D2566_Y));
KC_OAI21_X2 D2383 ( .B0(D12854_Q), .B1(D12785_Y), .A(D12777_Y),     .Y(D2383_Y));
KC_OAI21_X2 D2382 ( .B0(D12933_Y), .B1(D13010_Y), .A(D12947_Y),     .Y(D2382_Y));
KC_OAI21_X2 D2381 ( .B0(D13001_Y), .B1(D13010_Y), .A(D12947_Y),     .Y(D2381_Y));
KC_OAI21_X2 D2238 ( .B0(D10846_Y), .B1(D11305_Y), .A(D11256_Y),     .Y(D2238_Y));
KC_OAI21_X2 D2062 ( .B0(D1990_Y), .B1(D622_Y), .A(D8156_Y),     .Y(D2062_Y));
KC_OAI21_X2 D1768 ( .B0(D7538_Y), .B1(D5704_Y), .A(D5747_Y),     .Y(D1768_Y));
KC_OAI21_X2 D1624 ( .B0(D7496_Y), .B1(D7316_Y), .A(D7337_Y),     .Y(D1624_Y));
KC_OAI21_X2 D1623 ( .B0(D4568_Q), .B1(D4567_Q), .A(D1706_Y),     .Y(D1623_Y));
KC_OAI21_X2 D1622 ( .B0(D3112_Y), .B1(D1607_Y), .A(D4688_Y),     .Y(D1622_Y));
KC_OAI21_X2 D1620 ( .B0(D1411_Y), .B1(D3717_Y), .A(D5215_Y),     .Y(D1620_Y));
KC_OAI21_X2 D1477 ( .B0(D1525_Y), .B1(D2737_Y), .A(D2850_Y),     .Y(D1477_Y));
KC_OAI21_X2 D1471 ( .B0(D2939_Y), .B1(D2819_Y), .A(D265_Q),     .Y(D1471_Y));
KC_OAI21_X2 D1468 ( .B0(D3256_Y), .B1(D1426_Y), .A(D6344_Q),     .Y(D1468_Y));
KC_OAI21_X2 D1346 ( .B0(D11591_Y), .B1(D11565_Y), .A(D11536_Y),     .Y(D1346_Y));
KC_OAI21_X2 D1286 ( .B0(D11591_Y), .B1(D11566_Y), .A(D11536_Y),     .Y(D1286_Y));
KC_OAI21_X2 D1285 ( .B0(D11547_Y), .B1(D11548_Y), .A(D11536_Y),     .Y(D1285_Y));
KC_OAI21_X2 D1284 ( .B0(D11547_Y), .B1(D11591_Y), .A(D11536_Y),     .Y(D1284_Y));
KC_OAI21_X2 D1006 ( .B0(D11365_Y), .B1(D981_Y), .A(D2244_Y),     .Y(D1006_Y));
KC_OAI21_X2 D1005 ( .B0(D11358_Y), .B1(D980_Y), .A(D11386_Y),     .Y(D1005_Y));
KC_OAI21_X2 D888 ( .B0(D817_Q), .B1(D14109_Q), .A(D13985_Y),     .Y(D888_Y));
KC_OAI21_X2 D883 ( .B0(D10241_Y), .B1(D9494_Y), .A(D9584_Y),     .Y(D883_Y));
KC_OAI21_X2 D769 ( .B0(D777_Y), .B1(D14097_Y), .A(D13350_Y),     .Y(D769_Y));
KC_OAI21_X2 D653 ( .B0(D12749_Q), .B1(D822_Q), .A(D12707_Y),     .Y(D653_Y));
KC_OAI21_X2 D649 ( .B0(D8083_Y), .B1(D8088_Y), .A(D9444_Y),     .Y(D649_Y));
KC_OAI21_X2 D575 ( .B0(D1412_Y), .B1(D1413_Y), .A(D5215_Y),     .Y(D575_Y));
KC_OAI21_X2 D477 ( .B0(D3408_Y), .B1(D5038_Y), .A(D6449_Y),     .Y(D477_Y));
KC_OAI21_X2 D476 ( .B0(D1567_Y), .B1(D5020_Y), .A(D5021_Y),     .Y(D476_Y));
KC_OAI21_X2 D475 ( .B0(D5019_Y), .B1(D6438_Y), .A(D6455_Y),     .Y(D475_Y));
KC_OAI21_X2 D440 ( .B0(D3478_Y), .B1(D438_Y), .A(D4903_Y), .Y(D440_Y));
KC_OAI21_X2 D350 ( .B0(D40_Q), .B1(D8970_Y), .A(D7447_Y), .Y(D350_Y));
KC_OAI21_X2 D319 ( .B0(D7361_Y), .B1(D9058_Y), .A(D8983_Y),     .Y(D319_Y));
KC_OAI21_X2 D294 ( .B0(D276_Y), .B1(D7452_Y), .A(D7450_Y), .Y(D294_Y));
KC_OAI21_X2 D260 ( .B0(D243_Y), .B1(D293_Y), .A(D6058_Y), .Y(D260_Y));
KC_OAI21_X2 D259 ( .B0(D5909_Y), .B1(D7381_Y), .A(D5933_Y),     .Y(D259_Y));
KC_OAI21_X2 D99 ( .B0(D1413_Y), .B1(D3717_Y), .A(D5215_Y), .Y(D99_Y));
KC_BUF_X1 D16608 ( .Y(D16608_Y), .A(D16641_Y));
KC_BUF_X1 D16403 ( .Y(D16403_Y), .A(D776_Y));
KC_BUF_X1 D16377 ( .Y(D16377_Y), .A(D965_Y));
KC_BUF_X1 D16376 ( .Y(D16376_Y), .A(D965_Y));
KC_BUF_X1 D16267 ( .Y(D16267_Y), .A(D14858_Y));
KC_BUF_X1 D16195 ( .Y(D16195_Y), .A(D13186_Y));
KC_BUF_X1 D16126 ( .Y(D16126_Y), .A(D16087_Y));
KC_BUF_X1 D16121 ( .Y(D16121_Y), .A(D14574_Y));
KC_BUF_X1 D16066 ( .Y(D16066_Y), .A(D16052_Y));
KC_BUF_X1 D16016 ( .Y(D16016_Y), .A(D2525_Y));
KC_BUF_X1 D16015 ( .Y(D16015_Y), .A(D16017_Y));
KC_BUF_X1 D15927 ( .Y(D15927_Y), .A(D15699_Y));
KC_BUF_X1 D15838 ( .Y(D15838_Y), .A(D15678_Y));
KC_BUF_X1 D15774 ( .Y(D15774_Y), .A(D15576_Y));
KC_BUF_X1 D15765 ( .Y(D15765_Y), .A(D15673_Y));
KC_BUF_X1 D15652 ( .Y(D15652_Y), .A(D965_Y));
KC_BUF_X1 D15648 ( .Y(D15648_Y), .A(D15594_Y));
KC_BUF_X1 D15113 ( .Y(D15113_Y), .A(D15680_Y));
KC_BUF_X1 D14859 ( .Y(D14859_Y), .A(D940_Y));
KC_BUF_X1 D14858 ( .Y(D14858_Y), .A(D9360_Y));
KC_BUF_X1 D14856 ( .Y(D14856_Y), .A(D14799_Y));
KC_BUF_X1 D14811 ( .Y(D14811_Y), .A(D14812_Y));
KC_BUF_X1 D14810 ( .Y(D14810_Y), .A(D14779_Y));
KC_BUF_X1 D14774 ( .Y(D14774_Y), .A(D14783_Y));
KC_BUF_X1 D14773 ( .Y(D14773_Y), .A(D14782_Y));
KC_BUF_X1 D14772 ( .Y(D14772_Y), .A(D14780_Y));
KC_BUF_X1 D14771 ( .Y(D14771_Y), .A(D14781_Y));
KC_BUF_X1 D14760 ( .Y(D14760_Y), .A(D15569_Y));
KC_BUF_X1 D14759 ( .Y(D14759_Y), .A(D14778_Y));
KC_BUF_X1 D14291 ( .Y(D14291_Y), .A(D14858_Y));
KC_BUF_X1 D14288 ( .Y(D14288_Y), .A(D14858_Y));
KC_BUF_X1 D14224 ( .Y(D14224_Y), .A(D13444_Y));
KC_BUF_X1 D14057 ( .Y(D14057_Y), .A(D13394_Y));
KC_BUF_X1 D13738 ( .Y(D13738_Y), .A(D2429_Y));
KC_BUF_X1 D13242 ( .Y(D13242_Y), .A(D12280_Y));
KC_BUF_X1 D13186 ( .Y(D13186_Y), .A(D2455_Y));
KC_BUF_X1 D13185 ( .Y(D13185_Y), .A(D12280_Y));
KC_BUF_X1 D13153 ( .Y(D13153_Y), .A(D9361_Q));
KC_BUF_X1 D12901 ( .Y(D12901_Y), .A(D12280_Y));
KC_BUF_X1 D12900 ( .Y(D12900_Y), .A(D12280_Y));
KC_BUF_X1 D12898 ( .Y(D12898_Y), .A(D12280_Y));
KC_BUF_X1 D12734 ( .Y(D12734_Y), .A(D12280_Y));
KC_BUF_X1 D12662 ( .Y(D12662_Y), .A(D12280_Y));
KC_BUF_X1 D12258 ( .Y(D12258_Y), .A(D12280_Y));
KC_BUF_X1 D12182 ( .Y(D12182_Y), .A(D12144_Y));
KC_BUF_X1 D12135 ( .Y(D12135_Y), .A(D12134_Y));
KC_BUF_X1 D11438 ( .Y(D11438_Y), .A(D8267_Y));
KC_BUF_X1 D11308 ( .Y(D11308_Y), .A(D169_Y));
KC_BUF_X1 D11098 ( .Y(D11098_Y), .A(D10624_Y));
KC_BUF_X1 D10985 ( .Y(D10985_Y), .A(D8267_Y));
KC_BUF_X1 D10864 ( .Y(D10864_Y), .A(D11446_Y));
KC_BUF_X1 D10861 ( .Y(D10861_Y), .A(D1823_Y));
KC_BUF_X1 D10776 ( .Y(D10776_Y), .A(D10767_Y));
KC_BUF_X1 D10775 ( .Y(D10775_Y), .A(D10192_Y));
KC_BUF_X1 D10770 ( .Y(D10770_Y), .A(D8060_Y));
KC_BUF_X1 D10766 ( .Y(D10766_Y), .A(D9555_Y));
KC_BUF_X1 D10765 ( .Y(D10765_Y), .A(D8267_Y));
KC_BUF_X1 D10181 ( .Y(D10181_Y), .A(D1702_Y));
KC_BUF_X1 D10105 ( .Y(D10105_Y), .A(D1677_Y));
KC_BUF_X1 D9970 ( .Y(D9970_Y), .A(D10083_Y));
KC_BUF_X1 D9592 ( .Y(D9592_Y), .A(D2068_Y));
KC_BUF_X1 D9542 ( .Y(D9542_Y), .A(D2168_Q));
KC_BUF_X1 D9538 ( .Y(D9538_Y), .A(D12280_Y));
KC_BUF_X1 D9431 ( .Y(D9431_Y), .A(D8246_Q));
KC_BUF_X1 D9375 ( .Y(D9375_Y), .A(D12280_Y));
KC_BUF_X1 D9374 ( .Y(D9374_Y), .A(D12280_Y));
KC_BUF_X1 D9345 ( .Y(D9345_Y), .A(D726_Y));
KC_BUF_X1 D9249 ( .Y(D9249_Y), .A(D7660_Y));
KC_BUF_X1 D9247 ( .Y(D9247_Y), .A(D7785_Y));
KC_BUF_X1 D9246 ( .Y(D9246_Y), .A(D9223_Y));
KC_BUF_X1 D9200 ( .Y(D9200_Y), .A(D7135_Y));
KC_BUF_X1 D9193 ( .Y(D9193_Y), .A(D6360_Y));
KC_BUF_X1 D9128 ( .Y(D9128_Y), .A(D9358_Y));
KC_BUF_X1 D8786 ( .Y(D8786_Y), .A(D9010_Y));
KC_BUF_X1 D8779 ( .Y(D8779_Y), .A(D9358_Y));
KC_BUF_X1 D8774 ( .Y(D8774_Y), .A(D8892_Y));
KC_BUF_X1 D8773 ( .Y(D8773_Y), .A(D7272_Y));
KC_BUF_X1 D8685 ( .Y(D8685_Y), .A(D9949_Y));
KC_BUF_X1 D8684 ( .Y(D8684_Y), .A(D8674_Y));
KC_BUF_X1 D8683 ( .Y(D8683_Y), .A(D8712_Q));
KC_BUF_X1 D8431 ( .Y(D8431_Y), .A(D8013_Y));
KC_BUF_X1 D8430 ( .Y(D8430_Y), .A(D8013_Y));
KC_BUF_X1 D8300 ( .Y(D8300_Y), .A(D12280_Y));
KC_BUF_X1 D8212 ( .Y(D8212_Y), .A(D8013_Y));
KC_BUF_X1 D8211 ( .Y(D8211_Y), .A(D8177_Y));
KC_BUF_X1 D8210 ( .Y(D8210_Y), .A(D7990_Y));
KC_BUF_X1 D7950 ( .Y(D7950_Y), .A(D3647_Q));
KC_BUF_X1 D7775 ( .Y(D7775_Y), .A(D6209_Y));
KC_BUF_X1 D7701 ( .Y(D7701_Y), .A(D4630_Y));
KC_BUF_X1 D7641 ( .Y(D7641_Y), .A(D7609_Y));
KC_BUF_X1 D7571 ( .Y(D7571_Y), .A(D5930_Y));
KC_BUF_X1 D7446 ( .Y(D7446_Y), .A(D1963_Y));
KC_BUF_X1 D7376 ( .Y(D7376_Y), .A(D7460_Y));
KC_BUF_X1 D7361 ( .Y(D7361_Y), .A(D7460_Y));
KC_BUF_X1 D7125 ( .Y(D7125_Y), .A(D204_Y));
KC_BUF_X1 D6794 ( .Y(D6794_Y), .A(D1823_Y));
KC_BUF_X1 D6793 ( .Y(D6793_Y), .A(D6592_Y));
KC_BUF_X1 D6792 ( .Y(D6792_Y), .A(D6260_Y));
KC_BUF_X1 D6791 ( .Y(D6791_Y), .A(D6591_Y));
KC_BUF_X1 D6369 ( .Y(D6369_Y), .A(D7952_Y));
KC_BUF_X1 D6356 ( .Y(D6356_Y), .A(D6337_Y));
KC_BUF_X1 D6315 ( .Y(D6315_Y), .A(D6286_Y));
KC_BUF_X1 D6312 ( .Y(D6312_Y), .A(D3355_Y));
KC_BUF_X1 D6245 ( .Y(D6245_Y), .A(D1747_Y));
KC_BUF_X1 D6244 ( .Y(D6244_Y), .A(D6232_Y));
KC_BUF_X1 D6242 ( .Y(D6242_Y), .A(D6177_Y));
KC_BUF_X1 D6241 ( .Y(D6241_Y), .A(D6137_Y));
KC_BUF_X1 D6240 ( .Y(D6240_Y), .A(D6169_Y));
KC_BUF_X1 D6239 ( .Y(D6239_Y), .A(D3225_Y));
KC_BUF_X1 D6238 ( .Y(D6238_Y), .A(D7692_Y));
KC_BUF_X1 D6160 ( .Y(D6160_Y), .A(D16754_Y));
KC_BUF_X1 D6159 ( .Y(D6159_Y), .A(D4804_Y));
KC_BUF_X1 D6157 ( .Y(D6157_Y), .A(D8152_Y));
KC_BUF_X1 D6155 ( .Y(D6155_Y), .A(D1008_Y));
KC_BUF_X1 D6153 ( .Y(D6153_Y), .A(D6163_Y));
KC_BUF_X1 D6108 ( .Y(D6108_Y), .A(D9014_Y));
KC_BUF_X1 D6107 ( .Y(D6107_Y), .A(D4455_Y));
KC_BUF_X1 D6102 ( .Y(D6102_Y), .A(D7730_Y));
KC_BUF_X1 D6100 ( .Y(D6100_Y), .A(D6337_Y));
KC_BUF_X1 D5908 ( .Y(D5908_Y), .A(D6127_Y));
KC_BUF_X1 D5522 ( .Y(D5522_Y), .A(D9555_Y));
KC_BUF_X1 D5449 ( .Y(D5449_Y), .A(D9555_Y));
KC_BUF_X1 D5377 ( .Y(D5377_Y), .A(D5104_Y));
KC_BUF_X1 D5376 ( .Y(D5376_Y), .A(D5102_Y));
KC_BUF_X1 D5295 ( .Y(D5295_Y), .A(D5271_Y));
KC_BUF_X1 D5214 ( .Y(D5214_Y), .A(D497_Y));
KC_BUF_X1 D4940 ( .Y(D4940_Y), .A(D6448_Y));
KC_BUF_X1 D4785 ( .Y(D4785_Y), .A(D4817_Q));
KC_BUF_X1 D4702 ( .Y(D4702_Y), .A(D3210_Y));
KC_BUF_X1 D4616 ( .Y(D4616_Y), .A(D341_Y));
KC_BUF_X1 D4613 ( .Y(D4613_Y), .A(D4598_Y));
KC_BUF_X1 D4607 ( .Y(D4607_Y), .A(D6171_Y));
KC_BUF_X1 D4525 ( .Y(D4525_Y), .A(D4562_Q));
KC_BUF_X1 D4450 ( .Y(D4450_Y), .A(D1582_Y));
KC_BUF_X1 D4366 ( .Y(D4366_Y), .A(D6136_Y));
KC_BUF_X1 D4104 ( .Y(D4104_Y), .A(D4442_Y));
KC_BUF_X1 D4103 ( .Y(D4103_Y), .A(D4432_Y));
KC_BUF_X1 D3848 ( .Y(D3848_Y), .A(D5379_Y));
KC_BUF_X1 D3552 ( .Y(D3552_Y), .A(D16006_Y));
KC_BUF_X1 D3542 ( .Y(D3542_Y), .A(D7795_Y));
KC_BUF_X1 D3458 ( .Y(D3458_Y), .A(D3465_Y));
KC_BUF_X1 D3342 ( .Y(D3342_Y), .A(D12653_Y));
KC_BUF_X1 D3337 ( .Y(D3337_Y), .A(D3433_Y));
KC_BUF_X1 D3036 ( .Y(D3036_Y), .A(D6127_Y));
KC_BUF_X1 D2954 ( .Y(D2954_Y), .A(D15246_Y));
KC_BUF_X1 D2953 ( .Y(D2953_Y), .A(D6209_Y));
KC_BUF_X1 D2853 ( .Y(D2853_Y), .A(D2939_Y));
KC_BUF_X1 D2781 ( .Y(D2781_Y), .A(D2788_Y));
KC_BUF_X1 D2716 ( .Y(D2716_Y), .A(D264_Q));
KC_BUF_X1 D2627 ( .Y(D2627_Y), .A(D14858_Y));
KC_BUF_X1 D2500 ( .Y(D2500_Y), .A(D14905_Y));
KC_BUF_X1 D2277 ( .Y(D2277_Y), .A(D8267_Y));
KC_BUF_X1 D2032 ( .Y(D2032_Y), .A(D9725_Y));
KC_BUF_X1 D2030 ( .Y(D2030_Y), .A(D8700_Y));
KC_BUF_X1 D1905 ( .Y(D1905_Y), .A(D9058_Y));
KC_BUF_X1 D1900 ( .Y(D1900_Y), .A(D7937_Y));
KC_BUF_X1 D1895 ( .Y(D1895_Y), .A(D8207_Y));
KC_BUF_X1 D1745 ( .Y(D1745_Y), .A(D1694_Y));
KC_BUF_X1 D1596 ( .Y(D1596_Y), .A(D8267_Y));
KC_BUF_X1 D1454 ( .Y(D1454_Y), .A(D3104_Y));
KC_BUF_X1 D1453 ( .Y(D1453_Y), .A(D3250_Y));
KC_BUF_X1 D957 ( .Y(D957_Y), .A(D10319_Y));
KC_BUF_X1 D877 ( .Y(D877_Y), .A(D15575_Y));
KC_BUF_X1 D762 ( .Y(D762_Y), .A(D15581_Y));
KC_BUF_X1 D760 ( .Y(D760_Y), .A(D6521_Y));
KC_BUF_X1 D407 ( .Y(D407_Y), .A(D4630_Y));
KC_BUF_X1 D255 ( .Y(D255_Y), .A(D6110_Y));
KC_BUF_X1 D98 ( .Y(D98_Y), .A(D10735_Y));
KC_OAI22_X1 D16194 ( .A1(D16224_Y), .B0(D15476_Y), .B1(D16193_Y),     .A0(D15501_Y), .Y(D16194_Y));
KC_OAI22_X1 D15549 ( .A1(D15520_Y), .B0(D15424_Y), .B1(D15516_Y),     .A0(D15607_Y), .Y(D15549_Y));
KC_OAI22_X1 D15546 ( .A1(D15657_Y), .B0(D15489_Y), .B1(D15464_Y),     .A0(D2614_Y), .Y(D15546_Y));
KC_OAI22_X1 D15545 ( .A1(D2607_Y), .B0(D15473_Y), .B1(D15626_Y),     .A0(D15632_Y), .Y(D15545_Y));
KC_OAI22_X1 D15542 ( .A1(D15465_Y), .B0(D15471_Y), .B1(D15467_Y),     .A0(D14863_Y), .Y(D15542_Y));
KC_OAI22_X1 D15427 ( .A1(D15551_Y), .B0(D15357_Y), .B1(D15532_Y),     .A0(D15402_Y), .Y(D15427_Y));
KC_OAI22_X1 D15414 ( .A1(D15530_Y), .B0(D15344_Y), .B1(D15523_Y),     .A0(D15521_Y), .Y(D15414_Y));
KC_OAI22_X1 D15413 ( .A1(D15374_Y), .B0(D15366_Y), .B1(D15388_Y),     .A0(D14777_Y), .Y(D15413_Y));
KC_OAI22_X1 D14860 ( .A1(D14839_Y), .B0(D879_Y), .B1(D15617_Y),     .A0(D14830_Y), .Y(D14860_Y));
KC_OAI22_X1 D14762 ( .A1(D14728_Y), .B0(D14719_Y), .B1(D14867_Y),     .A0(D14841_Y), .Y(D14762_Y));
KC_OAI22_X1 D14660 ( .A1(D14625_Y), .B0(D15363_Y), .B1(D771_Y),     .A0(D14749_Y), .Y(D14660_Y));
KC_OAI22_X1 D14504 ( .A1(D14507_Y), .B0(D14502_Y), .B1(D14497_Y),     .A0(D14688_Q), .Y(D14504_Y));
KC_OAI22_X1 D14487 ( .A1(D14486_Y), .B0(D1376_Q), .B1(D15226_Y),     .A0(D14490_Q), .Y(D14487_Y));
KC_OAI22_X1 D14464 ( .A1(D14414_Y), .B0(D1323_Q), .B1(D14418_Y),     .A0(D14475_Q), .Y(D14464_Y));
KC_OAI22_X1 D14463 ( .A1(D14430_Y), .B0(D15213_Q), .B1(D15165_Y),     .A0(D1321_Q), .Y(D14463_Y));
KC_OAI22_X1 D14461 ( .A1(D14413_Y), .B0(D15217_Q), .B1(D15172_Y),     .A0(D13815_Q), .Y(D14461_Y));
KC_OAI22_X1 D14460 ( .A1(D14424_Y), .B0(D1325_Q), .B1(D1269_Y),     .A0(D13814_Q), .Y(D14460_Y));
KC_OAI22_X1 D14370 ( .A1(D14440_Y), .B0(D15218_Q), .B1(D15107_Y),     .A0(D13771_Q), .Y(D14370_Y));
KC_OAI22_X1 D14364 ( .A1(D13719_Y), .B0(D1232_Q), .B1(D15106_Y),     .A0(D13761_Q), .Y(D14364_Y));
KC_OAI22_X1 D14362 ( .A1(D14356_Y), .B0(D2524_Q), .B1(D14348_Y),     .A0(D14375_Q), .Y(D14362_Y));
KC_OAI22_X1 D14290 ( .A1(D14275_Y), .B0(D14295_Y), .B1(D14204_Y),     .A0(D14275_Y), .Y(D14290_Y));
KC_OAI22_X1 D14064 ( .A1(D14065_Y), .B0(D16765_Y), .B1(D14097_Y),     .A0(D2514_Y), .Y(D14064_Y));
KC_OAI22_X1 D14063 ( .A1(D14065_Y), .B0(D13983_Y), .B1(D14097_Y),     .A0(D13984_Y), .Y(D14063_Y));
KC_OAI22_X1 D14062 ( .A1(D14065_Y), .B0(D13982_Y), .B1(D14097_Y),     .A0(D13986_Y), .Y(D14062_Y));
KC_OAI22_X1 D14061 ( .A1(D14065_Y), .B0(D14086_Y), .B1(D14097_Y),     .A0(D14087_Y), .Y(D14061_Y));
KC_OAI22_X1 D14060 ( .A1(D14065_Y), .B0(D14081_Y), .B1(D14097_Y),     .A0(D14088_Y), .Y(D14060_Y));
KC_OAI22_X1 D14059 ( .A1(D14065_Y), .B0(D14002_Y), .B1(D14097_Y),     .A0(D14001_Y), .Y(D14059_Y));
KC_OAI22_X1 D14058 ( .A1(D14065_Y), .B0(D13985_Y), .B1(D14097_Y),     .A0(D14004_Y), .Y(D14058_Y));
KC_OAI22_X1 D13963 ( .A1(D14683_Y), .B0(D13941_Y), .B1(D14047_Y),     .A0(D13926_Y), .Y(D13963_Y));
KC_OAI22_X1 D13691 ( .A1(D13665_Y), .B0(D2471_Y), .B1(D6407_Y),     .A0(D2426_Y), .Y(D13691_Y));
KC_OAI22_X1 D13690 ( .A1(D13655_Y), .B0(D13610_Y), .B1(D6407_Y),     .A0(D13555_Y), .Y(D13690_Y));
KC_OAI22_X1 D13689 ( .A1(D13656_Y), .B0(D2420_Y), .B1(D6407_Y),     .A0(D13547_Y), .Y(D13689_Y));
KC_OAI22_X1 D13592 ( .A1(D13542_Y), .B0(D13555_Y), .B1(D14212_Y),     .A0(D13562_Y), .Y(D13592_Y));
KC_OAI22_X1 D13582 ( .A1(D13666_Y), .B0(D16767_Y), .B1(D6407_Y),     .A0(D13429_Y), .Y(D13582_Y));
KC_OAI22_X1 D13581 ( .A1(D14222_Y), .B0(D2421_Y), .B1(D6407_Y),     .A0(D13554_Y), .Y(D13581_Y));
KC_OAI22_X1 D13508 ( .A1(D13414_Y), .B0(D13309_Y), .B1(D13475_Y),     .A0(D13338_Y), .Y(D13508_Y));
KC_OAI22_X1 D13486 ( .A1(D13446_Y), .B0(D13445_Y), .B1(D870_Y),     .A0(D13440_Y), .Y(D13486_Y));
KC_OAI22_X1 D13366 ( .A1(D12772_Y), .B0(D13321_Y), .B1(D13319_Y),     .A0(D2448_Y), .Y(D13366_Y));
KC_OAI22_X1 D13244 ( .A1(D13224_Y), .B0(D13241_Y), .B1(D13282_Y),     .A0(D13245_Y), .Y(D13244_Y));
KC_OAI22_X1 D12822 ( .A1(D12784_Y), .B0(D12799_Y), .B1(D12696_Y),     .A0(D12808_Y), .Y(D12822_Y));
KC_OAI22_X1 D12821 ( .A1(D12702_Y), .B0(D12825_Y), .B1(D12808_Y),     .A0(D12800_Y), .Y(D12821_Y));
KC_OAI22_X1 D12818 ( .A1(D12792_Y), .B0(D12809_Y), .B1(D12807_Y),     .A0(D12808_Y), .Y(D12818_Y));
KC_OAI22_X1 D12817 ( .A1(D12791_Y), .B0(D12798_Y), .B1(D12711_Y),     .A0(D12808_Y), .Y(D12817_Y));
KC_OAI22_X1 D12730 ( .A1(D12699_Y), .B0(D12696_Y), .B1(D12325_Y),     .A0(D12784_Y), .Y(D12730_Y));
KC_OAI22_X1 D12727 ( .A1(D12699_Y), .B0(D12711_Y), .B1(D12715_Y),     .A0(D12791_Y), .Y(D12727_Y));
KC_OAI22_X1 D12726 ( .A1(D12699_Y), .B0(D12702_Y), .B1(D12248_Y),     .A0(D12825_Y), .Y(D12726_Y));
KC_OAI22_X1 D12724 ( .A1(D12699_Y), .B0(D12807_Y), .B1(D12716_Y),     .A0(D12792_Y), .Y(D12724_Y));
KC_OAI22_X1 D12664 ( .A1(D16_Y), .B0(D396_Y), .B1(D560_Y),     .A0(D6342_Y), .Y(D12664_Y));
KC_OAI22_X1 D12328 ( .A1(D12771_Y), .B0(D12321_Y), .B1(D12313_Y),     .A0(D12315_Y), .Y(D12328_Y));
KC_OAI22_X1 D12327 ( .A1(D12888_Y), .B0(D12313_Y), .B1(D12314_Y),     .A0(D12315_Y), .Y(D12327_Y));
KC_OAI22_X1 D12211 ( .A1(D12208_Y), .B0(D11657_Y), .B1(D12194_Y),     .A0(D10179_Y), .Y(D12211_Y));
KC_OAI22_X1 D11233 ( .A1(D2261_Y), .B0(D8146_Y), .B1(D11737_Y),     .A0(D10803_Y), .Y(D11233_Y));
KC_OAI22_X1 D9975 ( .A1(D8769_Y), .B0(D9972_Y), .B1(D9968_Y),     .A0(D9964_Y), .Y(D9975_Y));
KC_OAI22_X1 D9974 ( .A1(D8767_Y), .B0(D9973_Y), .B1(D216_Y),     .A0(D9963_Y), .Y(D9974_Y));
KC_OAI22_X1 D9969 ( .A1(D212_Y), .B0(D223_Y), .B1(D216_Y),     .A0(D9956_Y), .Y(D9969_Y));
KC_OAI22_X1 D9930 ( .A1(D9923_Y), .B0(D9973_Y), .B1(D9968_Y),     .A0(D9967_Y), .Y(D9930_Y));
KC_OAI22_X1 D9929 ( .A1(D9924_Y), .B0(D9971_Y), .B1(D9968_Y),     .A0(D9965_Y), .Y(D9929_Y));
KC_OAI22_X1 D9541 ( .A1(D9528_Y), .B0(D9502_Y), .B1(D9512_Y),     .A0(D9539_Y), .Y(D9541_Y));
KC_OAI22_X1 D9428 ( .A1(D8156_Y), .B0(D8148_Q), .B1(D9405_Y),     .A0(D826_Q), .Y(D9428_Y));
KC_OAI22_X1 D9203 ( .A1(D382_Y), .B0(D8971_Y), .B1(D2099_Y),     .A0(D9266_Y), .Y(D9203_Y));
KC_OAI22_X1 D9201 ( .A1(D382_Y), .B0(D9014_Y), .B1(D2099_Y),     .A0(D7713_Y), .Y(D9201_Y));
KC_OAI22_X1 D9199 ( .A1(D382_Y), .B0(D9122_Y), .B1(D2099_Y),     .A0(D10160_Y), .Y(D9199_Y));
KC_OAI22_X1 D9197 ( .A1(D382_Y), .B0(D9109_Y), .B1(D2099_Y),     .A0(D10158_Y), .Y(D9197_Y));
KC_OAI22_X1 D9196 ( .A1(D417_Y), .B0(D9122_Y), .B1(D2099_Y),     .A0(D10159_Y), .Y(D9196_Y));
KC_OAI22_X1 D9195 ( .A1(D382_Y), .B0(D9109_Y), .B1(D2099_Y),     .A0(D481_Y), .Y(D9195_Y));
KC_OAI22_X1 D9194 ( .A1(D9168_Y), .B0(D10105_Y), .B1(D407_Y),     .A0(D2120_Y), .Y(D9194_Y));
KC_OAI22_X1 D9129 ( .A1(D2099_Y), .B0(D7469_Y), .B1(D11116_Y),     .A0(D9023_Q), .Y(D9129_Y));
KC_OAI22_X1 D9079 ( .A1(D2008_Y), .B0(D7510_Y), .B1(D9033_Y),     .A0(D9228_Y), .Y(D9079_Y));
KC_OAI22_X1 D25 ( .A1(D242_Y), .B0(D338_Y), .B1(D7485_Y),     .A0(D10043_Y), .Y(D25_Y));
KC_OAI22_X1 D8995 ( .A1(D1880_Y), .B0(D7510_Y), .B1(D8985_Y),     .A0(D2027_Y), .Y(D8995_Y));
KC_OAI22_X1 D8994 ( .A1(D1907_Y), .B0(D7510_Y), .B1(D9014_Y),     .A0(D8748_Y), .Y(D8994_Y));
KC_OAI22_X1 D8988 ( .A1(D9045_Y), .B0(D8980_Y), .B1(D10044_Y),     .A0(D7361_Y), .Y(D8988_Y));
KC_OAI22_X1 D8942 ( .A1(D1907_Y), .B0(D8877_Y), .B1(D1880_Y),     .A0(D8756_Y), .Y(D8942_Y));
KC_OAI22_X1 D8939 ( .A1(D242_Y), .B0(D9057_Y), .B1(D7485_Y),     .A0(D9017_Y), .Y(D8939_Y));
KC_OAI22_X1 D8935 ( .A1(D9996_Y), .B0(D282_Y), .B1(D7485_Y),     .A0(D8949_Y), .Y(D8935_Y));
KC_OAI22_X1 D8933 ( .A1(D242_Y), .B0(D8908_Y), .B1(D7485_Y),     .A0(D8949_Y), .Y(D8933_Y));
KC_OAI22_X1 D8931 ( .A1(D242_Y), .B0(D8971_Y), .B1(D7485_Y),     .A0(D9013_Y), .Y(D8931_Y));
KC_OAI22_X1 D8928 ( .A1(D242_Y), .B0(D9109_Y), .B1(D7485_Y),     .A0(D9016_Y), .Y(D8928_Y));
KC_OAI22_X1 D8881 ( .A1(D7323_Y), .B0(D9015_Y), .B1(D5703_Y),     .A0(D7183_Y), .Y(D8881_Y));
KC_OAI22_X1 D8680 ( .A1(D8669_Y), .B0(D223_Y), .B1(D9968_Y),     .A0(D173_Y), .Y(D8680_Y));
KC_OAI22_X1 D8511 ( .A1(D8537_Y), .B0(D8550_Y), .B1(D6924_Y),     .A0(D8502_Y), .Y(D8511_Y));
KC_OAI22_X1 D8507 ( .A1(D1115_Y), .B0(D8550_Y), .B1(D1831_Y),     .A0(D8502_Y), .Y(D8507_Y));
KC_OAI22_X1 D8220 ( .A1(D9517_Y), .B0(D9510_Y), .B1(D9545_Y),     .A0(D9574_Q), .Y(D8220_Y));
KC_OAI22_X1 D8208 ( .A1(D8144_Y), .B0(D8146_Y), .B1(D8170_Y),     .A0(D6772_Y), .Y(D8208_Y));
KC_OAI22_X1 D8206 ( .A1(D895_Y), .B0(D8146_Y), .B1(D6710_Y),     .A0(D6772_Y), .Y(D8206_Y));
KC_OAI22_X1 D8205 ( .A1(D8233_Y), .B0(D8146_Y), .B1(D8187_Y),     .A0(D6772_Y), .Y(D8205_Y));
KC_OAI22_X1 D8129 ( .A1(D8161_Y), .B0(D8146_Y), .B1(D8009_Y),     .A0(D6772_Y), .Y(D8129_Y));
KC_OAI22_X1 D8126 ( .A1(D8160_Y), .B0(D8146_Y), .B1(D8110_Y),     .A0(D6772_Y), .Y(D8126_Y));
KC_OAI22_X1 D8123 ( .A1(D9535_Y), .B0(D8093_Y), .B1(D8080_Y),     .A0(D8078_Y), .Y(D8123_Y));
KC_OAI22_X1 D7865 ( .A1(D6428_Y), .B0(D7839_Y), .B1(D7862_Y),     .A0(D6438_Y), .Y(D7865_Y));
KC_OAI22_X1 D7696 ( .A1(D2099_Y), .B0(D9186_Y), .B1(D5963_Y),     .A0(D6097_Y), .Y(D7696_Y));
KC_OAI22_X1 D7645 ( .A1(D2122_Y), .B0(D7671_Y), .B1(D382_Y),     .A0(D7470_Y), .Y(D7645_Y));
KC_OAI22_X1 D7570 ( .A1(D2122_Y), .B0(D7503_Y), .B1(D1865_Y),     .A0(D1872_Y), .Y(D7570_Y));
KC_OAI22_X1 D7454 ( .A1(D287_Y), .B0(D7984_Y), .B1(D7419_Y),     .A0(D10753_Q), .Y(D7454_Y));
KC_OAI22_X1 D7366 ( .A1(D5857_Y), .B0(D214_Y), .B1(D6038_Y),     .A0(D7325_Y), .Y(D7366_Y));
KC_OAI22_X1 D7118 ( .A1(D5769_Y), .B0(D7101_Y), .B1(D7096_Y),     .A0(D7290_Y), .Y(D7118_Y));
KC_OAI22_X1 D6946 ( .A1(D6961_Y), .B0(D8550_Y), .B1(D6916_Y),     .A0(D8502_Y), .Y(D6946_Y));
KC_OAI22_X1 D6941 ( .A1(D6959_Y), .B0(D8550_Y), .B1(D6929_Y),     .A0(D8502_Y), .Y(D6941_Y));
KC_OAI22_X1 D6518 ( .A1(D492_Y), .B0(D492_Y), .B1(D1937_Y),     .A0(D493_Y), .Y(D6518_Y));
KC_OAI22_X1 D6453 ( .A1(D4863_Y), .B0(D7850_Y), .B1(D469_Y),     .A0(D1699_Y), .Y(D6453_Y));
KC_OAI22_X1 D6246 ( .A1(D1765_Y), .B0(D1765_Y), .B1(D1765_Y),     .A0(D6252_Y), .Y(D6246_Y));
KC_OAI22_X1 D6059 ( .A1(D1722_Y), .B0(D6023_Y), .B1(D5792_Y),     .A0(D4417_Y), .Y(D6059_Y));
KC_OAI22_X1 D6053 ( .A1(D7429_Y), .B0(D5745_Y), .B1(D6099_Y),     .A0(D4305_Y), .Y(D6053_Y));
KC_OAI22_X1 D6052 ( .A1(D6023_Y), .B0(D6002_Y), .B1(D4454_Y),     .A0(D5641_Y), .Y(D6052_Y));
KC_OAI22_X1 D6051 ( .A1(D6012_Y), .B0(D7427_Y), .B1(D6061_Y),     .A0(D726_Y), .Y(D6051_Y));
KC_OAI22_X1 D5913 ( .A1(D287_Y), .B0(D246_Y), .B1(D5685_Y),     .A0(D6015_Y), .Y(D5913_Y));
KC_OAI22_X1 D5911 ( .A1(D5847_Y), .B0(D5839_Y), .B1(D7324_Y),     .A0(D5836_Y), .Y(D5911_Y));
KC_OAI22_X1 D5902 ( .A1(D6005_Y), .B0(D4298_Y), .B1(D4443_Y),     .A0(D4425_Y), .Y(D5902_Y));
KC_OAI22_X1 D5791 ( .A1(D1735_Y), .B0(D5758_Y), .B1(D4205_Y),     .A0(D200_Y), .Y(D5791_Y));
KC_OAI22_X1 D5785 ( .A1(D5912_Y), .B0(D7376_Y), .B1(D5891_Y),     .A0(D7164_Y), .Y(D5785_Y));
KC_OAI22_X1 D5779 ( .A1(D1736_Y), .B0(D5647_Y), .B1(D7197_Y),     .A0(D1617_Y), .Y(D5779_Y));
KC_OAI22_X1 D5778 ( .A1(D4166_Y), .B0(D5769_Y), .B1(D211_Y),     .A0(D5693_Q), .Y(D5778_Y));
KC_OAI22_X1 D5777 ( .A1(D5721_Y), .B0(D7266_Y), .B1(D5722_Y),     .A0(D9477_Y), .Y(D5777_Y));
KC_OAI22_X1 D5776 ( .A1(D5847_Y), .B0(D5769_Y), .B1(D7227_Y),     .A0(D5763_Y), .Y(D5776_Y));
KC_OAI22_X1 D5067 ( .A1(D4865_Y), .B0(D1564_Y), .B1(D4880_Y),     .A0(D1561_Y), .Y(D5067_Y));
KC_OAI22_X1 D5065 ( .A1(D4889_Y), .B0(D4866_Y), .B1(D5043_Y),     .A0(D1564_Y), .Y(D5065_Y));
KC_OAI22_X1 D5061 ( .A1(D5004_Y), .B0(D5019_Y), .B1(D5043_Y),     .A0(D1564_Y), .Y(D5061_Y));
KC_OAI22_X1 D5060 ( .A1(D5020_Y), .B0(D3509_Y), .B1(D4882_Y),     .A0(D4900_Y), .Y(D5060_Y));
KC_OAI22_X1 D4976 ( .A1(D4891_Y), .B0(D3429_Y), .B1(D4914_Y),     .A0(D4912_Y), .Y(D4976_Y));
KC_OAI22_X1 D4948 ( .A1(D4941_Y), .B0(D3400_Y), .B1(D4906_Y),     .A0(D3373_Q), .Y(D4948_Y));
KC_OAI22_X1 D4937 ( .A1(D4972_Y), .B0(D1537_Y), .B1(D4905_Y),     .A0(D4919_Y), .Y(D4937_Y));
KC_OAI22_X1 D4934 ( .A1(D4894_Y), .B0(D4959_Y), .B1(D4881_Y),     .A0(D4892_Y), .Y(D4934_Y));
KC_OAI22_X1 D4931 ( .A1(D4922_Y), .B0(D1532_Y), .B1(D4869_Y),     .A0(D3402_Y), .Y(D4931_Y));
KC_OAI22_X1 D4929 ( .A1(D4865_Y), .B0(D1564_Y), .B1(D4882_Y),     .A0(D3499_Y), .Y(D4929_Y));
KC_OAI22_X1 D4705 ( .A1(D3229_Y), .B0(D1622_Y), .B1(D4733_Y),     .A0(D3232_Y), .Y(D4705_Y));
KC_OAI22_X1 D4400 ( .A1(D4374_Y), .B0(D4277_Y), .B1(D4349_Y),     .A0(D4097_Y), .Y(D4400_Y));
KC_OAI22_X1 D4379 ( .A1(D6034_Y), .B0(D4094_Y), .B1(D4347_Y),     .A0(D4357_Y), .Y(D4379_Y));
KC_OAI22_X1 D4376 ( .A1(D5876_Y), .B0(D4097_Y), .B1(D4347_Y),     .A0(D4306_Y), .Y(D4376_Y));
KC_OAI22_X1 D4372 ( .A1(D4324_Y), .B0(D4390_Y), .B1(D4391_Y),     .A0(D4394_Y), .Y(D4372_Y));
KC_OAI22_X1 D4367 ( .A1(D4319_Y), .B0(D4381_Y), .B1(D4273_Y),     .A0(D4312_Y), .Y(D4367_Y));
KC_OAI22_X1 D4365 ( .A1(D7100_Y), .B0(D4306_Y), .B1(D4304_Y),     .A0(D7460_Y), .Y(D4365_Y));
KC_OAI22_X1 D4364 ( .A1(D4284_Y), .B0(D4304_Y), .B1(D4397_Y),     .A0(D7512_Y), .Y(D4364_Y));
KC_OAI22_X1 D4222 ( .A1(D5847_Y), .B0(D7376_Y), .B1(D5758_Y),     .A0(D94_Y), .Y(D4222_Y));
KC_OAI22_X1 D4221 ( .A1(D4205_Y), .B0(D4440_Y), .B1(D1722_Y),     .A0(D94_Y), .Y(D4221_Y));
KC_OAI22_X1 D3554 ( .A1(D3594_Y), .B0(D4916_Y), .B1(D3405_Y),     .A0(D3400_Y), .Y(D3554_Y));
KC_OAI22_X1 D3548 ( .A1(D4881_Y), .B0(D3532_Y), .B1(D3371_Y),     .A0(D3576_Q), .Y(D3548_Y));
KC_OAI22_X1 D3546 ( .A1(D4882_Y), .B0(D3509_Y), .B1(D3521_Y),     .A0(D3599_Y), .Y(D3546_Y));
KC_OAI22_X1 D3462 ( .A1(D3516_Y), .B0(D3372_Q), .B1(D4867_Y),     .A0(D446_Q), .Y(D3462_Y));
KC_OAI22_X1 D3455 ( .A1(D3414_Y), .B0(D4895_Y), .B1(D3537_Y),     .A0(D4909_Y), .Y(D3455_Y));
KC_OAI22_X1 D3451 ( .A1(D3564_Y), .B0(D3476_Y), .B1(D3472_Y),     .A0(D3472_Y), .Y(D3451_Y));
KC_OAI22_X1 D3450 ( .A1(D3538_Y), .B0(D5044_Y), .B1(D4895_Y),     .A0(D3371_Y), .Y(D3450_Y));
KC_OAI22_X1 D3255 ( .A1(D1455_Y), .B0(D3349_Y), .B1(D1428_Y),     .A0(D4592_Y), .Y(D3255_Y));
KC_OAI22_X1 D3246 ( .A1(D3380_Y), .B0(D3225_Y), .B1(D4606_Y),     .A0(D3302_Q), .Y(D3246_Y));
KC_OAI22_X1 D2951 ( .A1(D2950_Y), .B0(D3070_Y), .B1(D2903_Y),     .A0(D2997_Y), .Y(D2951_Y));
KC_OAI22_X1 D2774 ( .A1(D2738_Y), .B0(D2739_Y), .B1(D2793_Y),     .A0(D2848_Y), .Y(D2774_Y));
KC_OAI22_X1 D2771 ( .A1(D2740_Y), .B0(D2848_Y), .B1(D2765_Y),     .A0(D2759_Y), .Y(D2771_Y));
KC_OAI22_X1 D2453 ( .A1(D12876_Y), .B0(D13473_Y), .B1(D13401_Y),     .A0(D13307_Y), .Y(D2453_Y));
KC_OAI22_X1 D2452 ( .A1(D12878_Y), .B0(D13473_Y), .B1(D13319_Y),     .A0(D2449_Y), .Y(D2452_Y));
KC_OAI22_X1 D2451 ( .A1(D13702_Y), .B0(D13309_Y), .B1(D13319_Y),     .A0(D13367_Y), .Y(D2451_Y));
KC_OAI22_X1 D2450 ( .A1(D13469_Y), .B0(D13322_Y), .B1(D13401_Y),     .A0(D2434_Y), .Y(D2450_Y));
KC_OAI22_X1 D2442 ( .A1(D14200_Y), .B0(D13622_Y), .B1(D6407_Y),     .A0(D13546_Y), .Y(D2442_Y));
KC_OAI22_X1 D2441 ( .A1(D13664_Y), .B0(D13641_Y), .B1(D6407_Y),     .A0(D13428_Y), .Y(D2441_Y));
KC_OAI22_X1 D2331 ( .A1(D12770_Y), .B0(D12313_Y), .B1(D12309_Y),     .A0(D12315_Y), .Y(D2331_Y));
KC_OAI22_X1 D2050 ( .A1(D242_Y), .B0(D9014_Y), .B1(D7485_Y),     .A0(D8950_Y), .Y(D2050_Y));
KC_OAI22_X1 D2044 ( .A1(D2099_Y), .B0(D7469_Y), .B1(D12287_Y),     .A0(D9019_Q), .Y(D2044_Y));
KC_OAI22_X1 D2040 ( .A1(D9391_Y), .B0(D1988_Y), .B1(D9401_Y),     .A0(D8084_Y), .Y(D2040_Y));
KC_OAI22_X1 D1906 ( .A1(D7324_Y), .B0(D7984_Y), .B1(D4304_Y),     .A0(D9478_Y), .Y(D1906_Y));
KC_OAI22_X1 D1753 ( .A1(D4284_Y), .B0(D7376_Y), .B1(D1714_Y),     .A0(D726_Y), .Y(D1753_Y));
KC_OAI22_X1 D1752 ( .A1(D1718_Y), .B0(D6050_Y), .B1(D213_Y),     .A0(D7295_Y), .Y(D1752_Y));
KC_OAI22_X1 D1742 ( .A1(D6960_Y), .B0(D8550_Y), .B1(D6989_Y),     .A0(D8502_Y), .Y(D1742_Y));
KC_OAI22_X1 D1616 ( .A1(D4358_Y), .B0(D4187_Y), .B1(D4374_Y),     .A0(D4354_Y), .Y(D1616_Y));
KC_OAI22_X1 D1615 ( .A1(D4374_Y), .B0(D4284_Y), .B1(D4347_Y),     .A0(D4304_Y), .Y(D1615_Y));
KC_OAI22_X1 D1605 ( .A1(D4838_Y), .B0(D4915_Y), .B1(D4748_Y),     .A0(D4925_Y), .Y(D1605_Y));
KC_OAI22_X1 D1604 ( .A1(D4910_Y), .B0(D5035_Y), .B1(D4960_Y),     .A0(D3599_Y), .Y(D1604_Y));
KC_OAI22_X1 D1603 ( .A1(D5043_Y), .B0(D1564_Y), .B1(D5020_Y),     .A0(D4882_Y), .Y(D1603_Y));
KC_OAI22_X1 D1452 ( .A1(D3393_Y), .B0(D3599_Y), .B1(D3415_Y),     .A0(D3375_Q), .Y(D1452_Y));
KC_OAI22_X1 D1449 ( .A1(D3405_Y), .B0(D5020_Y), .B1(D3537_Y),     .A0(D3527_Y), .Y(D1449_Y));
KC_OAI22_X1 D1448 ( .A1(D5044_Y), .B0(D4902_Y), .B1(D3528_Y),     .A0(D3416_Y), .Y(D1448_Y));
KC_OAI22_X1 D1102 ( .A1(D1116_Y), .B0(D8550_Y), .B1(D6931_Y),     .A0(D8502_Y), .Y(D1102_Y));
KC_OAI22_X1 D1098 ( .A1(D8536_Y), .B0(D8550_Y), .B1(D6927_Y),     .A0(D8502_Y), .Y(D1098_Y));
KC_OAI22_X1 D438 ( .A1(D4898_Y), .B0(D3415_Y), .B1(D3429_Y),     .A0(D3499_Y), .Y(D438_Y));
KC_OAI22_X1 D437 ( .A1(D6438_Y), .B0(D3423_Y), .B1(D4912_Y),     .A0(D3499_Y), .Y(D437_Y));
KC_OAI22_X1 D411 ( .A1(D5963_Y), .B0(D9115_Y), .B1(D9113_Y),     .A0(D7629_Y), .Y(D411_Y));
KC_OAI22_X1 D376 ( .A1(D7633_Y), .B0(D9122_Y), .B1(D2099_Y),     .A0(D7637_Y), .Y(D376_Y));
KC_OAI22_X1 D375 ( .A1(D382_Y), .B0(D7644_Y), .B1(D9113_Y),     .A0(D6023_Y), .Y(D375_Y));
KC_OAI22_X1 D345 ( .A1(D336_Y), .B0(D4590_Y), .B1(D4602_Y),     .A0(D3321_Y), .Y(D345_Y));
KC_OAI22_X1 D218 ( .A1(D7211_Y), .B0(D4444_Y), .B1(D7204_Y),     .A0(D203_Y), .Y(D218_Y));
KC_OAI22_X1 D92 ( .A1(D3235_Y), .B0(D1672_Y), .B1(D4580_Y),     .A0(D3117_Y), .Y(D92_Y));
KC_AOI21_X1 D16510 ( .B0(D16530_Y), .Y(D16510_Y), .A(D1343_Y),     .B1(D16485_Y));
KC_AOI21_X1 D16509 ( .B0(D16502_Y), .Y(D16509_Y), .A(D16496_Y),     .B1(D16504_Y));
KC_AOI21_X1 D16450 ( .B0(D16413_Y), .Y(D16450_Y), .A(D16407_Y),     .B1(D16464_Y));
KC_AOI21_X1 D16447 ( .B0(D15985_Y), .Y(D16447_Y), .A(D16407_Y),     .B1(D16464_Y));
KC_AOI21_X1 D16445 ( .B0(D16462_Y), .Y(D16445_Y), .A(D16407_Y),     .B1(D16420_Y));
KC_AOI21_X1 D16124 ( .B0(D16104_Y), .Y(D16124_Y), .A(D16111_Y),     .B1(D16088_Y));
KC_AOI21_X1 D16122 ( .B0(D16126_Y), .Y(D16122_Y), .A(D16155_Y),     .B1(D16102_Y));
KC_AOI21_X1 D15984 ( .B0(D14248_Y), .Y(D15984_Y), .A(D14070_Y),     .B1(D877_Y));
KC_AOI21_X1 D15983 ( .B0(D15684_Y), .Y(D15983_Y), .A(D14070_Y),     .B1(D14250_Y));
KC_AOI21_X1 D15982 ( .B0(D15684_Y), .Y(D15982_Y), .A(D14070_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15980 ( .B0(D14251_Y), .Y(D15980_Y), .A(D14062_Y),     .B1(D16381_Y));
KC_AOI21_X1 D15979 ( .B0(D15684_Y), .Y(D15979_Y), .A(D14070_Y),     .B1(D14251_Y));
KC_AOI21_X1 D15978 ( .B0(D14251_Y), .Y(D15978_Y), .A(D14070_Y),     .B1(D877_Y));
KC_AOI21_X1 D15977 ( .B0(D15927_Y), .Y(D15977_Y), .A(D14062_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15976 ( .B0(D14250_Y), .Y(D15976_Y), .A(D14070_Y),     .B1(D877_Y));
KC_AOI21_X1 D15975 ( .B0(D15999_Q), .Y(D15975_Y), .A(D15968_Y),     .B1(D15960_Y));
KC_AOI21_X1 D15931 ( .B0(D15927_Y), .Y(D15931_Y), .A(D14062_Y),     .B1(D14251_Y));
KC_AOI21_X1 D15930 ( .B0(D14250_Y), .Y(D15930_Y), .A(D14062_Y),     .B1(D16381_Y));
KC_AOI21_X1 D15929 ( .B0(D16381_Y), .Y(D15929_Y), .A(D14062_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15924 ( .B0(D877_Y), .Y(D15924_Y), .A(D14070_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15923 ( .B0(D15997_Q), .Y(D15923_Y), .A(D15891_Y),     .B1(D15896_Y));
KC_AOI21_X1 D15922 ( .B0(D1229_Q), .Y(D15922_Y), .A(D15889_Y),     .B1(D15899_Y));
KC_AOI21_X1 D15919 ( .B0(D14248_Y), .Y(D15919_Y), .A(D14062_Y),     .B1(D16381_Y));
KC_AOI21_X1 D15855 ( .B0(D14251_Y), .Y(D15855_Y), .A(D14064_Y),     .B1(D16309_Y));
KC_AOI21_X1 D15854 ( .B0(D14250_Y), .Y(D15854_Y), .A(D14064_Y),     .B1(D16309_Y));
KC_AOI21_X1 D15853 ( .B0(D16309_Y), .Y(D15853_Y), .A(D14064_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15852 ( .B0(D14248_Y), .Y(D15852_Y), .A(D14064_Y),     .B1(D16309_Y));
KC_AOI21_X1 D15845 ( .B0(D14250_Y), .Y(D15845_Y), .A(D14063_Y),     .B1(D15586_Y));
KC_AOI21_X1 D15843 ( .B0(D14248_Y), .Y(D15843_Y), .A(D14063_Y),     .B1(D15586_Y));
KC_AOI21_X1 D15842 ( .B0(D15688_Y), .Y(D15842_Y), .A(D14063_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15841 ( .B0(D15586_Y), .Y(D15841_Y), .A(D14063_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15840 ( .B0(D14251_Y), .Y(D15840_Y), .A(D14063_Y),     .B1(D15586_Y));
KC_AOI21_X1 D15839 ( .B0(D16351_Y), .Y(D15839_Y), .A(D14064_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15776 ( .B0(D15683_Y), .Y(D15776_Y), .A(D14059_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15775 ( .B0(D15587_Y), .Y(D15775_Y), .A(D14059_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15772 ( .B0(D15664_Y), .Y(D15772_Y), .A(D14061_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15771 ( .B0(D14248_Y), .Y(D15771_Y), .A(D14059_Y),     .B1(D15587_Y));
KC_AOI21_X1 D15768 ( .B0(D14251_Y), .Y(D15768_Y), .A(D14059_Y),     .B1(D15587_Y));
KC_AOI21_X1 D15767 ( .B0(D2666_Y), .Y(D15767_Y), .A(D14061_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15766 ( .B0(D14248_Y), .Y(D15766_Y), .A(D14061_Y),     .B1(D2666_Y));
KC_AOI21_X1 D15761 ( .B0(D14251_Y), .Y(D15761_Y), .A(D14061_Y),     .B1(D2666_Y));
KC_AOI21_X1 D15760 ( .B0(D14250_Y), .Y(D15760_Y), .A(D14061_Y),     .B1(D2666_Y));
KC_AOI21_X1 D15759 ( .B0(D15587_Y), .Y(D15759_Y), .A(D14059_Y),     .B1(D14250_Y));
KC_AOI21_X1 D15757 ( .B0(D15592_Y), .Y(D15757_Y), .A(D14060_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15756 ( .B0(D14248_Y), .Y(D15756_Y), .A(D14060_Y),     .B1(D15592_Y));
KC_AOI21_X1 D15753 ( .B0(D14250_Y), .Y(D15753_Y), .A(D14060_Y),     .B1(D15592_Y));
KC_AOI21_X1 D15752 ( .B0(D14251_Y), .Y(D15752_Y), .A(D14060_Y),     .B1(D15592_Y));
KC_AOI21_X1 D15750 ( .B0(D14248_Y), .Y(D15750_Y), .A(D14058_Y),     .B1(D16278_Y));
KC_AOI21_X1 D15749 ( .B0(D16278_Y), .Y(D15749_Y), .A(D14058_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15747 ( .B0(D14904_Y), .Y(D15747_Y), .A(D14060_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15658 ( .B0(D15562_Y), .Y(D15658_Y), .A(D14846_Y),     .B1(D15149_Y));
KC_AOI21_X1 D15657 ( .B0(D15562_Y), .Y(D15657_Y), .A(D2610_Y),     .B1(D14187_Y));
KC_AOI21_X1 D15559 ( .B0(D15563_Y), .Y(D15559_Y), .A(D15539_Y),     .B1(D15952_Y));
KC_AOI21_X1 D15554 ( .B0(D15563_Y), .Y(D15554_Y), .A(D15528_Y),     .B1(D2644_Y));
KC_AOI21_X1 D15551 ( .B0(D15563_Y), .Y(D15551_Y), .A(D15526_Y),     .B1(D14184_Y));
KC_AOI21_X1 D15544 ( .B0(D14719_Y), .Y(D15544_Y), .A(D15633_Y),     .B1(D2607_Y));
KC_AOI21_X1 D15543 ( .B0(D15562_Y), .Y(D15543_Y), .A(D15484_Y),     .B1(D14514_Y));
KC_AOI21_X1 D15417 ( .B0(D15363_Y), .Y(D15417_Y), .A(D15513_Y),     .B1(D15530_Y));
KC_AOI21_X1 D15412 ( .B0(D15563_Y), .Y(D15412_Y), .A(D15367_Y),     .B1(D14513_Y));
KC_AOI21_X1 D15227 ( .B0(D16008_Q), .Y(D15227_Y), .A(D15223_Y),     .B1(D15224_Y));
KC_AOI21_X1 D15207 ( .B0(D984_Y), .Y(D15207_Y), .A(D14067_Y),     .B1(D14760_Y));
KC_AOI21_X1 D15206 ( .B0(D984_Y), .Y(D15206_Y), .A(D14076_Y),     .B1(D15128_Y));
KC_AOI21_X1 D15205 ( .B0(D15993_Q), .Y(D15205_Y), .A(D15166_Y),     .B1(D15971_Y));
KC_AOI21_X1 D15203 ( .B0(D16011_Q), .Y(D15203_Y), .A(D15105_Y),     .B1(D15110_Y));
KC_AOI21_X1 D15201 ( .B0(D14247_Y), .Y(D15201_Y), .A(D14076_Y),     .B1(D15128_Y));
KC_AOI21_X1 D15200 ( .B0(D15838_Y), .Y(D15200_Y), .A(D14076_Y),     .B1(D14247_Y));
KC_AOI21_X1 D15197 ( .B0(D16012_Q), .Y(D15197_Y), .A(D1272_Y),     .B1(D15964_Y));
KC_AOI21_X1 D15193 ( .B0(D14251_Y), .Y(D15193_Y), .A(D14076_Y),     .B1(D15128_Y));
KC_AOI21_X1 D15192 ( .B0(D14251_Y), .Y(D15192_Y), .A(D14067_Y),     .B1(D14760_Y));
KC_AOI21_X1 D15190 ( .B0(D15789_Y), .Y(D15190_Y), .A(D14067_Y),     .B1(D13540_Y));
KC_AOI21_X1 D15189 ( .B0(D15838_Y), .Y(D15189_Y), .A(D14076_Y),     .B1(D13540_Y));
KC_AOI21_X1 D15186 ( .B0(D15789_Y), .Y(D15186_Y), .A(D14067_Y),     .B1(D14247_Y));
KC_AOI21_X1 D15185 ( .B0(D14247_Y), .Y(D15185_Y), .A(D14067_Y),     .B1(D14760_Y));
KC_AOI21_X1 D15121 ( .B0(D15838_Y), .Y(D15121_Y), .A(D14076_Y),     .B1(D14251_Y));
KC_AOI21_X1 D15120 ( .B0(D15789_Y), .Y(D15120_Y), .A(D14067_Y),     .B1(D14251_Y));
KC_AOI21_X1 D15119 ( .B0(D15128_Y), .Y(D15119_Y), .A(D14076_Y),     .B1(D14249_Y));
KC_AOI21_X1 D15118 ( .B0(D16009_Q), .Y(D15118_Y), .A(D15098_Y),     .B1(D15101_Y));
KC_AOI21_X1 D15115 ( .B0(D14248_Y), .Y(D15115_Y), .A(D14067_Y),     .B1(D15789_Y));
KC_AOI21_X1 D15114 ( .B0(D15927_Y), .Y(D15114_Y), .A(D14062_Y),     .B1(D14250_Y));
KC_AOI21_X1 D15066 ( .B0(D14248_Y), .Y(D15066_Y), .A(D14062_Y),     .B1(D15927_Y));
KC_AOI21_X1 D15064 ( .B0(D14248_Y), .Y(D15064_Y), .A(D14063_Y),     .B1(D15688_Y));
KC_AOI21_X1 D15063 ( .B0(D2676_Y), .Y(D15063_Y), .A(D14058_Y),     .B1(D14250_Y));
KC_AOI21_X1 D15060 ( .B0(D14248_Y), .Y(D15060_Y), .A(D14064_Y),     .B1(D16351_Y));
KC_AOI21_X1 D15057 ( .B0(D16351_Y), .Y(D15057_Y), .A(D14064_Y),     .B1(D14250_Y));
KC_AOI21_X1 D15054 ( .B0(D15688_Y), .Y(D15054_Y), .A(D14063_Y),     .B1(D14250_Y));
KC_AOI21_X1 D15052 ( .B0(D15688_Y), .Y(D15052_Y), .A(D14063_Y),     .B1(D14251_Y));
KC_AOI21_X1 D15051 ( .B0(D16351_Y), .Y(D15051_Y), .A(D14064_Y),     .B1(D14251_Y));
KC_AOI21_X1 D14974 ( .B0(D15664_Y), .Y(D14974_Y), .A(D14061_Y),     .B1(D14251_Y));
KC_AOI21_X1 D14973 ( .B0(D15664_Y), .Y(D14973_Y), .A(D14061_Y),     .B1(D14250_Y));
KC_AOI21_X1 D14971 ( .B0(D14904_Y), .Y(D14971_Y), .A(D14060_Y),     .B1(D14251_Y));
KC_AOI21_X1 D14968 ( .B0(D14904_Y), .Y(D14968_Y), .A(D14060_Y),     .B1(D14250_Y));
KC_AOI21_X1 D14863 ( .B0(D15562_Y), .Y(D14863_Y), .A(D14850_Y),     .B1(D14262_Y));
KC_AOI21_X1 D14862 ( .B0(D15562_Y), .Y(D14862_Y), .A(D14853_Y),     .B1(D15079_Y));
KC_AOI21_X1 D14777 ( .B0(D15563_Y), .Y(D14777_Y), .A(D15538_Y),     .B1(D2578_Y));
KC_AOI21_X1 D14776 ( .B0(D13988_Y), .Y(D14776_Y), .A(D13932_Y),     .B1(D14707_Y));
KC_AOI21_X1 D14671 ( .B0(D14694_Y), .Y(D14671_Y), .A(D103_Y),     .B1(D14647_Y));
KC_AOI21_X1 D14659 ( .B0(D13931_Y), .Y(D14659_Y), .A(D13934_Y),     .B1(D14744_Y));
KC_AOI21_X1 D14658 ( .B0(D14776_Y), .Y(D14658_Y), .A(D13934_Y),     .B1(D14670_Y));
KC_AOI21_X1 D14560 ( .B0(D14708_Y), .Y(D14560_Y), .A(D14531_Y),     .B1(D14541_Y));
KC_AOI21_X1 D14506 ( .B0(D2512_Y), .Y(D14506_Y), .A(D14567_Y),     .B1(D14516_Y));
KC_AOI21_X1 D14505 ( .B0(D14687_Q), .Y(D14505_Y), .A(D14504_Y),     .B1(D2545_Y));
KC_AOI21_X1 D14503 ( .B0(D12173_Y), .Y(D14503_Y), .A(D14567_Y),     .B1(D14497_Y));
KC_AOI21_X1 D14462 ( .B0(D15113_Y), .Y(D14462_Y), .A(D14071_Y),     .B1(D14247_Y));
KC_AOI21_X1 D14459 ( .B0(D15113_Y), .Y(D14459_Y), .A(D14071_Y),     .B1(D13540_Y));
KC_AOI21_X1 D14227 ( .B0(D15683_Y), .Y(D14227_Y), .A(D14059_Y),     .B1(D14220_Y));
KC_AOI21_X1 D14226 ( .B0(D14248_Y), .Y(D14226_Y), .A(D14059_Y),     .B1(D15683_Y));
KC_AOI21_X1 D14225 ( .B0(D15683_Y), .Y(D14225_Y), .A(D14059_Y),     .B1(D14250_Y));
KC_AOI21_X1 D14223 ( .B0(D14248_Y), .Y(D14223_Y), .A(D14058_Y),     .B1(D2676_Y));
KC_AOI21_X1 D14147 ( .B0(D87_Y), .Y(D14147_Y), .A(D14026_Y),     .B1(D750_Y));
KC_AOI21_X1 D14146 ( .B0(D13304_Y), .Y(D14146_Y), .A(D14026_Y),     .B1(D13291_Y));
KC_AOI21_X1 D14145 ( .B0(D13310_Y), .Y(D14145_Y), .A(D14026_Y),     .B1(D13303_Y));
KC_AOI21_X1 D14144 ( .B0(D2495_Y), .Y(D14144_Y), .A(D14026_Y),     .B1(D2437_Y));
KC_AOI21_X1 D14142 ( .B0(D13449_Y), .Y(D14142_Y), .A(D14074_Y),     .B1(D14264_Q));
KC_AOI21_X1 D14066 ( .B0(D14046_Y), .Y(D14066_Y), .A(D14676_Y),     .B1(D13941_Y));
KC_AOI21_X1 D13968 ( .B0(D13970_Y), .Y(D13968_Y), .A(D573_Y),     .B1(D14047_Y));
KC_AOI21_X1 D13793 ( .B0(D984_Y), .Y(D13793_Y), .A(D14071_Y),     .B1(D14856_Y));
KC_AOI21_X1 D13792 ( .B0(D2500_Y), .Y(D13792_Y), .A(D14068_Y),     .B1(D14247_Y));
KC_AOI21_X1 D13789 ( .B0(D2500_Y), .Y(D13789_Y), .A(D14068_Y),     .B1(D14220_Y));
KC_AOI21_X1 D13786 ( .B0(D14220_Y), .Y(D13786_Y), .A(D14068_Y),     .B1(D15648_Y));
KC_AOI21_X1 D13784 ( .B0(D14247_Y), .Y(D13784_Y), .A(D14068_Y),     .B1(D15648_Y));
KC_AOI21_X1 D13783 ( .B0(D2500_Y), .Y(D13783_Y), .A(D14068_Y),     .B1(D13540_Y));
KC_AOI21_X1 D13781 ( .B0(D984_Y), .Y(D13781_Y), .A(D14068_Y),     .B1(D15648_Y));
KC_AOI21_X1 D13780 ( .B0(D14247_Y), .Y(D13780_Y), .A(D14071_Y),     .B1(D14856_Y));
KC_AOI21_X1 D13744 ( .B0(D14220_Y), .Y(D13744_Y), .A(D14071_Y),     .B1(D14856_Y));
KC_AOI21_X1 D13740 ( .B0(D14856_Y), .Y(D13740_Y), .A(D14071_Y),     .B1(D13540_Y));
KC_AOI21_X1 D13739 ( .B0(D984_Y), .Y(D13739_Y), .A(D14068_Y),     .B1(D2500_Y));
KC_AOI21_X1 D13734 ( .B0(D15113_Y), .Y(D13734_Y), .A(D14071_Y),     .B1(D14220_Y));
KC_AOI21_X1 D13732 ( .B0(D15648_Y), .Y(D13732_Y), .A(D14068_Y),     .B1(D13540_Y));
KC_AOI21_X1 D13681 ( .B0(D14250_Y), .Y(D13681_Y), .A(D14073_Y),     .B1(D762_Y));
KC_AOI21_X1 D13680 ( .B0(D15691_Y), .Y(D13680_Y), .A(D14073_Y),     .B1(D14250_Y));
KC_AOI21_X1 D13678 ( .B0(D984_Y), .Y(D13678_Y), .A(D14073_Y),     .B1(D762_Y));
KC_AOI21_X1 D13677 ( .B0(D15691_Y), .Y(D13677_Y), .A(D14073_Y),     .B1(D13540_Y));
KC_AOI21_X1 D13676 ( .B0(D15691_Y), .Y(D13676_Y), .A(D14073_Y),     .B1(D14220_Y));
KC_AOI21_X1 D13675 ( .B0(D762_Y), .Y(D13675_Y), .A(D14073_Y),     .B1(D13540_Y));
KC_AOI21_X1 D13600 ( .B0(D13455_Y), .Y(D13600_Y), .A(D13543_Y),     .B1(D13462_Y));
KC_AOI21_X1 D13598 ( .B0(D13556_Y), .Y(D13598_Y), .A(D14074_Y),     .B1(D14243_Q));
KC_AOI21_X1 D13597 ( .B0(D13455_Y), .Y(D13597_Y), .A(D13567_Y),     .B1(D13462_Y));
KC_AOI21_X1 D13596 ( .B0(D13550_Y), .Y(D13596_Y), .A(D14074_Y),     .B1(D14244_Q));
KC_AOI21_X1 D13595 ( .B0(D13567_Y), .Y(D13595_Y), .A(D13527_Y),     .B1(D13514_Y));
KC_AOI21_X1 D13591 ( .B0(D13455_Y), .Y(D13591_Y), .A(D13548_Y),     .B1(D13462_Y));
KC_AOI21_X1 D13590 ( .B0(D2436_Y), .Y(D13590_Y), .A(D13527_Y),     .B1(D13514_Y));
KC_AOI21_X1 D13587 ( .B0(D13561_Y), .Y(D13587_Y), .A(D14074_Y),     .B1(D1066_Q));
KC_AOI21_X1 D13586 ( .B0(D13514_Y), .Y(D13586_Y), .A(D13529_Y),     .B1(D13543_Y));
KC_AOI21_X1 D13580 ( .B0(D13514_Y), .Y(D13580_Y), .A(D13529_Y),     .B1(D13548_Y));
KC_AOI21_X1 D13507 ( .B0(D13523_Y), .Y(D13507_Y), .A(D13532_Y),     .B1(D2438_Y));
KC_AOI21_X1 D13505 ( .B0(D13523_Y), .Y(D13505_Y), .A(D13535_Y),     .B1(D2435_Y));
KC_AOI21_X1 D13504 ( .B0(D13523_Y), .Y(D13504_Y), .A(D13535_Y),     .B1(D13466_Y));
KC_AOI21_X1 D13502 ( .B0(D13523_Y), .Y(D13502_Y), .A(D13532_Y),     .B1(D13458_Y));
KC_AOI21_X1 D13501 ( .B0(D13515_Q), .Y(D13501_Y), .A(D930_Q),     .B1(D12887_Y));
KC_AOI21_X1 D13497 ( .B0(D13393_Y), .Y(D13497_Y), .A(D13448_Y),     .B1(D13323_Y));
KC_AOI21_X1 D13496 ( .B0(D13455_Y), .Y(D13496_Y), .A(D13458_Y),     .B1(D13462_Y));
KC_AOI21_X1 D13490 ( .B0(D13450_Y), .Y(D13490_Y), .A(D14074_Y),     .B1(D14265_Q));
KC_AOI21_X1 D13489 ( .B0(D13455_Y), .Y(D13489_Y), .A(D2438_Y),     .B1(D13462_Y));
KC_AOI21_X1 D13485 ( .B0(D13455_Y), .Y(D13485_Y), .A(D2435_Y),     .B1(D13462_Y));
KC_AOI21_X1 D13482 ( .B0(D13422_Y), .Y(D13482_Y), .A(D14074_Y),     .B1(D14245_Q));
KC_AOI21_X1 D13371 ( .B0(D14024_Y), .Y(D13371_Y), .A(D13364_Y),     .B1(D12823_Y));
KC_AOI21_X1 D13367 ( .B0(D13329_Y), .Y(D13367_Y), .A(D13296_Y),     .B1(D13309_Y));
KC_AOI21_X1 D12963 ( .B0(D814_Q), .Y(D12963_Y), .A(D12995_Q),     .B1(D12873_Y));
KC_AOI21_X1 D12899 ( .B0(D855_Q), .Y(D12899_Y), .A(D954_Q),     .B1(D12875_Y));
KC_AOI21_X1 D12897 ( .B0(D13028_Y), .Y(D12897_Y), .A(D2398_Y),     .B1(D12878_Y));
KC_AOI21_X1 D12896 ( .B0(D13027_Y), .Y(D12896_Y), .A(D2397_Y),     .B1(D12876_Y));
KC_AOI21_X1 D12895 ( .B0(D13699_Y), .Y(D12895_Y), .A(D12933_Y),     .B1(D12772_Y));
KC_AOI21_X1 D12819 ( .B0(D12729_Y), .Y(D12819_Y), .A(D12804_Y),     .B1(D13268_Q));
KC_AOI21_X1 D12209 ( .B0(D12362_Y), .Y(D12209_Y), .A(D12276_Y),     .B1(D12801_Y));
KC_AOI21_X1 D11776 ( .B0(D10787_Y), .Y(D11776_Y), .A(D10803_Y),     .B1(D11753_Y));
KC_AOI21_X1 D11775 ( .B0(D10787_Y), .Y(D11775_Y), .A(D10803_Y),     .B1(D11770_Y));
KC_AOI21_X1 D11648 ( .B0(D10181_Y), .Y(D11648_Y), .A(D11645_Y),     .B1(D12197_Y));
KC_AOI21_X1 D11526 ( .B0(D7991_Y), .Y(D11526_Y), .A(D1936_Y),     .B1(D13058_Y));
KC_AOI21_X1 D11525 ( .B0(D7991_Y), .Y(D11525_Y), .A(D1936_Y),     .B1(D1264_Y));
KC_AOI21_X1 D11524 ( .B0(D7991_Y), .Y(D11524_Y), .A(D1936_Y),     .B1(D13072_Y));
KC_AOI21_X1 D11523 ( .B0(D7991_Y), .Y(D11523_Y), .A(D1936_Y),     .B1(D12517_Y));
KC_AOI21_X1 D11522 ( .B0(D7991_Y), .Y(D11522_Y), .A(D1936_Y),     .B1(D12022_Y));
KC_AOI21_X1 D11521 ( .B0(D7991_Y), .Y(D11521_Y), .A(D1936_Y),     .B1(D13057_Y));
KC_AOI21_X1 D11520 ( .B0(D7991_Y), .Y(D11520_Y), .A(D1936_Y),     .B1(D12538_Y));
KC_AOI21_X1 D11519 ( .B0(D7991_Y), .Y(D11519_Y), .A(D1936_Y),     .B1(D12568_Y));
KC_AOI21_X1 D11518 ( .B0(D7991_Y), .Y(D11518_Y), .A(D1936_Y),     .B1(D12570_Y));
KC_AOI21_X1 D11517 ( .B0(D7991_Y), .Y(D11517_Y), .A(D1936_Y),     .B1(D12070_Y));
KC_AOI21_X1 D11516 ( .B0(D7991_Y), .Y(D11516_Y), .A(D1936_Y),     .B1(D13103_Y));
KC_AOI21_X1 D11515 ( .B0(D7991_Y), .Y(D11515_Y), .A(D1936_Y),     .B1(D13074_Y));
KC_AOI21_X1 D11514 ( .B0(D7991_Y), .Y(D11514_Y), .A(D1936_Y),     .B1(D12537_Y));
KC_AOI21_X1 D11513 ( .B0(D7991_Y), .Y(D11513_Y), .A(D1936_Y),     .B1(D12061_Y));
KC_AOI21_X1 D11443 ( .B0(D7991_Y), .Y(D11443_Y), .A(D10748_Y),     .B1(D11428_Y));
KC_AOI21_X1 D11442 ( .B0(D8210_Y), .Y(D11442_Y), .A(D1936_Y),     .B1(D12436_Y));
KC_AOI21_X1 D11441 ( .B0(D8210_Y), .Y(D11441_Y), .A(D10748_Y),     .B1(D2269_Y));
KC_AOI21_X1 D11440 ( .B0(D7990_Y), .Y(D11440_Y), .A(D1936_Y),     .B1(D12484_Y));
KC_AOI21_X1 D11439 ( .B0(D8210_Y), .Y(D11439_Y), .A(D1936_Y),     .B1(D12489_Y));
KC_AOI21_X1 D11378 ( .B0(D8210_Y), .Y(D11378_Y), .A(D10748_Y),     .B1(D12439_Y));
KC_AOI21_X1 D11376 ( .B0(D7990_Y), .Y(D11376_Y), .A(D10748_Y),     .B1(D12491_Y));
KC_AOI21_X1 D11312 ( .B0(D10787_Y), .Y(D11312_Y), .A(D10803_Y),     .B1(D12423_Y));
KC_AOI21_X1 D11311 ( .B0(D7990_Y), .Y(D11311_Y), .A(D10748_Y),     .B1(D2276_Y));
KC_AOI21_X1 D11310 ( .B0(D10787_Y), .Y(D11310_Y), .A(D10803_Y),     .B1(D12375_Y));
KC_AOI21_X1 D11309 ( .B0(D10787_Y), .Y(D11309_Y), .A(D10803_Y),     .B1(D11878_Y));
KC_AOI21_X1 D11307 ( .B0(D10787_Y), .Y(D11307_Y), .A(D10803_Y),     .B1(D11834_Y));
KC_AOI21_X1 D11306 ( .B0(D10787_Y), .Y(D11306_Y), .A(D10803_Y),     .B1(D11837_Y));
KC_AOI21_X1 D11304 ( .B0(D8210_Y), .Y(D11304_Y), .A(D10748_Y),     .B1(D12391_Y));
KC_AOI21_X1 D11239 ( .B0(D10787_Y), .Y(D11239_Y), .A(D10803_Y),     .B1(D11218_Y));
KC_AOI21_X1 D11238 ( .B0(D10787_Y), .Y(D11238_Y), .A(D10803_Y),     .B1(D11699_Y));
KC_AOI21_X1 D11237 ( .B0(D10787_Y), .Y(D11237_Y), .A(D10803_Y),     .B1(D11697_Y));
KC_AOI21_X1 D11236 ( .B0(D10787_Y), .Y(D11236_Y), .A(D10803_Y),     .B1(D10754_Y));
KC_AOI21_X1 D11235 ( .B0(D10787_Y), .Y(D11235_Y), .A(D10803_Y),     .B1(D10675_Y));
KC_AOI21_X1 D11234 ( .B0(D10787_Y), .Y(D11234_Y), .A(D10803_Y),     .B1(D11222_Y));
KC_AOI21_X1 D11232 ( .B0(D10787_Y), .Y(D11232_Y), .A(D10803_Y),     .B1(D11214_Y));
KC_AOI21_X1 D11231 ( .B0(D10787_Y), .Y(D11231_Y), .A(D10803_Y),     .B1(D11754_Y));
KC_AOI21_X1 D10859 ( .B0(D2135_Y), .Y(D10859_Y), .A(D10849_Y),     .B1(D98_Y));
KC_AOI21_X1 D10774 ( .B0(D10787_Y), .Y(D10774_Y), .A(D10803_Y),     .B1(D10680_Y));
KC_AOI21_X1 D10773 ( .B0(D10787_Y), .Y(D10773_Y), .A(D10803_Y),     .B1(D10699_Y));
KC_AOI21_X1 D10772 ( .B0(D10787_Y), .Y(D10772_Y), .A(D10803_Y),     .B1(D10760_Y));
KC_AOI21_X1 D10769 ( .B0(D7990_Y), .Y(D10769_Y), .A(D10748_Y),     .B1(D10692_Y));
KC_AOI21_X1 D10088 ( .B0(D10074_Y), .Y(D10088_Y), .A(D10077_Y),     .B1(D10081_Y));
KC_AOI21_X1 D10054 ( .B0(D11114_Y), .Y(D10054_Y), .A(D6091_Y),     .B1(D2123_Y));
KC_AOI21_X1 D9973 ( .B0(D8702_Y), .Y(D9973_Y), .A(D201_Y),     .B1(D9961_Y));
KC_AOI21_X1 D9972 ( .B0(D9961_Y), .Y(D9972_Y), .A(D201_Y),     .B1(D9960_Y));
KC_AOI21_X1 D9971 ( .B0(D7882_Y), .Y(D9971_Y), .A(D201_Y),     .B1(D9960_Y));
KC_AOI21_X1 D9549 ( .B0(D9597_Y), .Y(D9549_Y), .A(D9548_Y),     .B1(D9219_Q));
KC_AOI21_X1 D9539 ( .B0(D2039_Y), .Y(D9539_Y), .A(D9532_Y),     .B1(D9512_Y));
KC_AOI21_X1 D9084 ( .B0(D9054_Y), .Y(D9084_Y), .A(D9061_Y),     .B1(D394_Y));
KC_AOI21_X1 D9081 ( .B0(D9054_Y), .Y(D9081_Y), .A(D9074_Y),     .B1(D9279_Q));
KC_AOI21_X1 D8941 ( .B0(D8898_Q), .Y(D8941_Y), .A(D25_Y),     .B1(D8883_Y));
KC_AOI21_X1 D8936 ( .B0(D8955_Q), .Y(D8936_Y), .A(D8928_Y),     .B1(D8901_Y));
KC_AOI21_X1 D8934 ( .B0(D8900_Y), .Y(D8934_Y), .A(D8935_Y),     .B1(D10047_Q));
KC_AOI21_X1 D8932 ( .B0(D305_Q), .Y(D8932_Y), .A(D8933_Y),     .B1(D8901_Y));
KC_AOI21_X1 D8930 ( .B0(D151_Q), .Y(D8930_Y), .A(D8931_Y),     .B1(D8901_Y));
KC_AOI21_X1 D8883 ( .B0(D5710_Y), .Y(D8883_Y), .A(D7361_Y),     .B1(D7396_Y));
KC_AOI21_X1 D8843 ( .B0(D8844_Y), .Y(D8843_Y), .A(D8780_Y),     .B1(D8791_Y));
KC_AOI21_X1 D8841 ( .B0(D8821_Q), .Y(D8841_Y), .A(D8839_Y),     .B1(D8840_Y));
KC_AOI21_X1 D8785 ( .B0(D8823_Q), .Y(D8785_Y), .A(D8765_Y),     .B1(D8833_Y));
KC_AOI21_X1 D8784 ( .B0(D205_Y), .Y(D8784_Y), .A(D9981_Q),     .B1(D212_Y));
KC_AOI21_X1 D8780 ( .B0(D8797_Y), .Y(D8780_Y), .A(D8827_Y),     .B1(D8791_Y));
KC_AOI21_X1 D8433 ( .B0(D8240_Y), .Y(D8433_Y), .A(D8502_Y),     .B1(D3916_Y));
KC_AOI21_X1 D8432 ( .B0(D8240_Y), .Y(D8432_Y), .A(D8502_Y),     .B1(D11887_Y));
KC_AOI21_X1 D8301 ( .B0(D8240_Y), .Y(D8301_Y), .A(D6772_Y),     .B1(D1552_Y));
KC_AOI21_X1 D8299 ( .B0(D8240_Y), .Y(D8299_Y), .A(D6772_Y),     .B1(D5429_Y));
KC_AOI21_X1 D8298 ( .B0(D8240_Y), .Y(D8298_Y), .A(D6772_Y),     .B1(D3923_Y));
KC_AOI21_X1 D8218 ( .B0(D8210_Y), .Y(D8218_Y), .A(D6772_Y),     .B1(D3829_Y));
KC_AOI21_X1 D8217 ( .B0(D8240_Y), .Y(D8217_Y), .A(D6772_Y),     .B1(D740_Y));
KC_AOI21_X1 D8216 ( .B0(D8210_Y), .Y(D8216_Y), .A(D6772_Y),     .B1(D3792_Y));
KC_AOI21_X1 D8214 ( .B0(D8240_Y), .Y(D8214_Y), .A(D6772_Y),     .B1(D5293_Y));
KC_AOI21_X1 D8213 ( .B0(D8210_Y), .Y(D8213_Y), .A(D6772_Y),     .B1(D6625_Y));
KC_AOI21_X1 D8209 ( .B0(D8240_Y), .Y(D8209_Y), .A(D6772_Y),     .B1(D5268_Y));
KC_AOI21_X1 D8127 ( .B0(D8210_Y), .Y(D8127_Y), .A(D6772_Y),     .B1(D6633_Y));
KC_AOI21_X1 D8124 ( .B0(D8115_Y), .Y(D8124_Y), .A(D9407_Y),     .B1(D8094_Y));
KC_AOI21_X1 D8029 ( .B0(D8073_Q), .Y(D8029_Y), .A(D8016_Y),     .B1(D7960_Y));
KC_AOI21_X1 D8028 ( .B0(D8210_Y), .Y(D8028_Y), .A(D8011_Y),     .B1(D6589_Y));
KC_AOI21_X1 D8027 ( .B0(D8210_Y), .Y(D8027_Y), .A(D8011_Y),     .B1(D5154_Y));
KC_AOI21_X1 D8026 ( .B0(D8210_Y), .Y(D8026_Y), .A(D8011_Y),     .B1(D5180_Y));
KC_AOI21_X1 D8025 ( .B0(D8210_Y), .Y(D8025_Y), .A(D8011_Y),     .B1(D5160_Y));
KC_AOI21_X1 D8024 ( .B0(D8210_Y), .Y(D8024_Y), .A(D8011_Y),     .B1(D6585_Y));
KC_AOI21_X1 D8023 ( .B0(D8210_Y), .Y(D8023_Y), .A(D8011_Y),     .B1(D5172_Y));
KC_AOI21_X1 D7951 ( .B0(D7888_Q), .Y(D7951_Y), .A(D7929_Y),     .B1(D7919_Y));
KC_AOI21_X1 D7872 ( .B0(D479_Q), .Y(D7872_Y), .A(D6441_Y),     .B1(D7856_Y));
KC_AOI21_X1 D7869 ( .B0(D7883_Q), .Y(D7869_Y), .A(D7855_Y),     .B1(D7852_Y));
KC_AOI21_X1 D7864 ( .B0(D7835_Y), .Y(D7864_Y), .A(D7833_Y),     .B1(D533_Q));
KC_AOI21_X1 D7642 ( .B0(D7627_Y), .Y(D7642_Y), .A(D6250_Y),     .B1(D7626_Y));
KC_AOI21_X1 D7569 ( .B0(D6174_Y), .Y(D7569_Y), .A(D7541_Y),     .B1(D7639_Y));
KC_AOI21_X1 D7451 ( .B0(D8153_Y), .Y(D7451_Y), .A(D8_Y), .B1(D7435_Y));
KC_AOI21_X1 D7449 ( .B0(D5867_Y), .Y(D7449_Y), .A(D7480_Q),     .B1(D7419_Y));
KC_AOI21_X1 D7367 ( .B0(D7330_Y), .Y(D7367_Y), .A(D7382_Y),     .B1(D7381_Y));
KC_AOI21_X1 D7364 ( .B0(D7263_Y), .Y(D7364_Y), .A(D5903_Y),     .B1(D7442_Y));
KC_AOI21_X1 D7276 ( .B0(D8742_Y), .Y(D7276_Y), .A(D204_Y),     .B1(D222_Y));
KC_AOI21_X1 D7127 ( .B0(D8706_Y), .Y(D7127_Y), .A(D5682_Y),     .B1(D7125_Y));
KC_AOI21_X1 D7001 ( .B0(D8466_Y), .Y(D7001_Y), .A(D8502_Y),     .B1(D7039_Y));
KC_AOI21_X1 D7000 ( .B0(D8466_Y), .Y(D7000_Y), .A(D8502_Y),     .B1(D5579_Y));
KC_AOI21_X1 D6999 ( .B0(D8466_Y), .Y(D6999_Y), .A(D8502_Y),     .B1(D5623_Y));
KC_AOI21_X1 D6998 ( .B0(D8466_Y), .Y(D6998_Y), .A(D8502_Y),     .B1(D6985_Y));
KC_AOI21_X1 D6997 ( .B0(D8466_Y), .Y(D6997_Y), .A(D8502_Y),     .B1(D7026_Y));
KC_AOI21_X1 D6996 ( .B0(D8466_Y), .Y(D6996_Y), .A(D8502_Y),     .B1(D1681_Y));
KC_AOI21_X1 D6945 ( .B0(D8466_Y), .Y(D6945_Y), .A(D8502_Y),     .B1(D5502_Y));
KC_AOI21_X1 D6884 ( .B0(D8240_Y), .Y(D6884_Y), .A(D8011_Y),     .B1(D976_Y));
KC_AOI21_X1 D6726 ( .B0(D8210_Y), .Y(D6726_Y), .A(D6772_Y),     .B1(D6725_Y));
KC_AOI21_X1 D6519 ( .B0(D6553_Q), .Y(D6519_Y), .A(D6513_Y),     .B1(D6554_Q));
KC_AOI21_X1 D6456 ( .B0(D4877_Y), .Y(D6456_Y), .A(D6437_Y),     .B1(D3408_Y));
KC_AOI21_X1 D6455 ( .B0(D4885_Y), .Y(D6455_Y), .A(D4995_Y),     .B1(D476_Y));
KC_AOI21_X1 D6450 ( .B0(D6415_Y), .Y(D6450_Y), .A(D6531_Y),     .B1(D6418_Y));
KC_AOI21_X1 D6411 ( .B0(D441_Y), .Y(D6411_Y), .A(D6365_Y),     .B1(D445_Q));
KC_AOI21_X1 D6314 ( .B0(D6298_Y), .Y(D6314_Y), .A(D6315_Y),     .B1(D6325_Y));
KC_AOI21_X1 D6243 ( .B0(D6227_Y), .Y(D6243_Y), .A(D6272_Y),     .B1(D6226_Y));
KC_AOI21_X1 D6162 ( .B0(D6184_Y), .Y(D6162_Y), .A(D6146_Y),     .B1(D6146_Y));
KC_AOI21_X1 D6105 ( .B0(D6106_Y), .Y(D6105_Y), .A(D7531_Y),     .B1(D6089_Y));
KC_AOI21_X1 D6058 ( .B0(D7295_Y), .Y(D6058_Y), .A(D6006_Y),     .B1(D4439_Y));
KC_AOI21_X1 D6050 ( .B0(D7429_Y), .Y(D6050_Y), .A(D6044_Y),     .B1(D7474_Y));
KC_AOI21_X1 D6049 ( .B0(D5869_Y), .Y(D6049_Y), .A(D1724_Y),     .B1(D1748_Y));
KC_AOI21_X1 D6042 ( .B0(D7353_Y), .Y(D6042_Y), .A(D5952_Y),     .B1(D5805_Y));
KC_AOI21_X1 D5916 ( .B0(D5684_Y), .Y(D5916_Y), .A(D7344_Y),     .B1(D5876_Y));
KC_AOI21_X1 D5915 ( .B0(D249_Y), .Y(D5915_Y), .A(D5894_Y),     .B1(D5870_Y));
KC_AOI21_X1 D5786 ( .B0(D5646_Y), .Y(D5786_Y), .A(D5788_Y),     .B1(D5798_Y));
KC_AOI21_X1 D5782 ( .B0(D5755_Y), .Y(D5782_Y), .A(D5881_Y),     .B1(D219_Y));
KC_AOI21_X1 D5059 ( .B0(D3524_Y), .Y(D5059_Y), .A(D5043_Y),     .B1(D5003_Y));
KC_AOI21_X1 D5053 ( .B0(D4999_Y), .Y(D5053_Y), .A(D5023_Y),     .B1(D4992_Y));
KC_AOI21_X1 D5050 ( .B0(D4983_Y), .Y(D5050_Y), .A(D6437_Y),     .B1(D5079_Y));
KC_AOI21_X1 D5046 ( .B0(D4983_Y), .Y(D5046_Y), .A(D6437_Y),     .B1(D5082_Y));
KC_AOI21_X1 D4944 ( .B0(D4946_Y), .Y(D4944_Y), .A(D3400_Y),     .B1(D4945_Y));
KC_AOI21_X1 D4943 ( .B0(D1537_Y), .Y(D4943_Y), .A(D4939_Y),     .B1(D4908_Y));
KC_AOI21_X1 D4936 ( .B0(D6449_Y), .Y(D4936_Y), .A(D4937_Y),     .B1(D4934_Y));
KC_AOI21_X1 D4709 ( .B0(D4694_Y), .Y(D4709_Y), .A(D371_Y),     .B1(D4572_Y));
KC_AOI21_X1 D4697 ( .B0(D4591_Y), .Y(D4697_Y), .A(D3097_Y),     .B1(D4673_Y));
KC_AOI21_X1 D4611 ( .B0(D3172_Y), .Y(D4611_Y), .A(D4591_Y),     .B1(D3250_Y));
KC_AOI21_X1 D4610 ( .B0(D4598_Y), .Y(D4610_Y), .A(D4613_Y),     .B1(D4817_Q));
KC_AOI21_X1 D4608 ( .B0(D3349_Y), .Y(D4608_Y), .A(D369_Y),     .B1(D3125_Y));
KC_AOI21_X1 D4371 ( .B0(D4173_Y), .Y(D4371_Y), .A(D6024_Y),     .B1(D4430_Y));
KC_AOI21_X1 D4219 ( .B0(D5936_Y), .Y(D4219_Y), .A(D4225_Y),     .B1(D4382_Y));
KC_AOI21_X1 D4210 ( .B0(D4136_Q), .Y(D4210_Y), .A(D5776_Y),     .B1(D1615_Y));
KC_AOI21_X1 D4033 ( .B0(D4036_Y), .Y(D4033_Y), .A(D4079_Y),     .B1(D4032_Y));
KC_AOI21_X1 D3553 ( .B0(D1570_Y), .Y(D3553_Y), .A(D3521_Y),     .B1(D3502_Y));
KC_AOI21_X1 D3543 ( .B0(D4983_Y), .Y(D3543_Y), .A(D3503_Y),     .B1(D3508_Y));
KC_AOI21_X1 D3467 ( .B0(D4897_Y), .Y(D3467_Y), .A(D3419_Y),     .B1(D3475_Y));
KC_AOI21_X1 D3464 ( .B0(D3433_Y), .Y(D3464_Y), .A(D4939_Y),     .B1(D4902_Y));
KC_AOI21_X1 D3459 ( .B0(D1537_Y), .Y(D3459_Y), .A(D3414_Y),     .B1(D3498_Y));
KC_AOI21_X1 D3454 ( .B0(D3458_Y), .Y(D3454_Y), .A(D3407_Y),     .B1(D3458_Y));
KC_AOI21_X1 D3344 ( .B0(D3343_Y), .Y(D3344_Y), .A(D1454_Y),     .B1(D3377_Y));
KC_AOI21_X1 D3340 ( .B0(D3376_Q), .Y(D3340_Y), .A(D3311_Y),     .B1(D3338_Y));
KC_AOI21_X1 D3257 ( .B0(D3267_Y), .Y(D3257_Y), .A(D3269_Y),     .B1(D4717_Y));
KC_AOI21_X1 D3241 ( .B0(D3261_Y), .Y(D3241_Y), .A(D3212_Y),     .B1(D3209_Y));
KC_AOI21_X1 D3240 ( .B0(D398_Y), .Y(D3240_Y), .A(D7641_Y),     .B1(D3218_Y));
KC_AOI21_X1 D3164 ( .B0(D4599_Y), .Y(D3164_Y), .A(D7641_Y),     .B1(D4600_Y));
KC_AOI21_X1 D3160 ( .B0(D3110_Y), .Y(D3160_Y), .A(D7641_Y),     .B1(D3102_Y));
KC_AOI21_X1 D3158 ( .B0(D3097_Y), .Y(D3158_Y), .A(D3098_Y),     .B1(D3061_Y));
KC_AOI21_X1 D3046 ( .B0(D3072_Y), .Y(D3046_Y), .A(D3031_Y),     .B1(D4512_Y));
KC_AOI21_X1 D3045 ( .B0(D4627_Y), .Y(D3045_Y), .A(D3091_Y),     .B1(D4525_Y));
KC_AOI21_X1 D2857 ( .B0(D2834_Y), .Y(D2857_Y), .A(D2761_Y),     .B1(D2820_Y));
KC_AOI21_X1 D2854 ( .B0(D2827_Y), .Y(D2854_Y), .A(D2760_Y),     .B1(D2820_Y));
KC_AOI21_X1 D2664 ( .B0(D16227_Y), .Y(D2664_Y), .A(D16260_Y),     .B1(D16263_Y));
KC_AOI21_X1 D2624 ( .B0(D14250_Y), .Y(D2624_Y), .A(D14058_Y),     .B1(D16278_Y));
KC_AOI21_X1 D2623 ( .B0(D14251_Y), .Y(D2623_Y), .A(D14058_Y),     .B1(D16278_Y));
KC_AOI21_X1 D2622 ( .B0(D2676_Y), .Y(D2622_Y), .A(D14058_Y),     .B1(D14249_Y));
KC_AOI21_X1 D2563 ( .B0(D14532_Y), .Y(D2563_Y), .A(D2545_Y),     .B1(D14499_Y));
KC_AOI21_X1 D2559 ( .B0(D14248_Y), .Y(D2559_Y), .A(D14060_Y),     .B1(D14904_Y));
KC_AOI21_X1 D2558 ( .B0(D14248_Y), .Y(D2558_Y), .A(D14061_Y),     .B1(D15664_Y));
KC_AOI21_X1 D2555 ( .B0(D2676_Y), .Y(D2555_Y), .A(D14058_Y),     .B1(D14251_Y));
KC_AOI21_X1 D2553 ( .B0(D14248_Y), .Y(D2553_Y), .A(D14076_Y),     .B1(D15838_Y));
KC_AOI21_X1 D2552 ( .B0(D14760_Y), .Y(D2552_Y), .A(D14067_Y),     .B1(D14249_Y));
KC_AOI21_X1 D2449 ( .B0(D13329_Y), .Y(D2449_Y), .A(D13296_Y),     .B1(D13473_Y));
KC_AOI21_X1 D2448 ( .B0(D13329_Y), .Y(D2448_Y), .A(D13296_Y),     .B1(D13321_Y));
KC_AOI21_X1 D2445 ( .B0(D13455_Y), .Y(D2445_Y), .A(D13466_Y),     .B1(D13462_Y));
KC_AOI21_X1 D2444 ( .B0(D2428_Y), .Y(D2444_Y), .A(D14074_Y),     .B1(D14242_Q));
KC_AOI21_X1 D2235 ( .B0(D8210_Y), .Y(D2235_Y), .A(D1936_Y),     .B1(D11947_Y));
KC_AOI21_X1 D2234 ( .B0(D8210_Y), .Y(D2234_Y), .A(D10748_Y),     .B1(D12492_Y));
KC_AOI21_X1 D2208 ( .B0(D7990_Y), .Y(D2208_Y), .A(D10748_Y),     .B1(D5339_Y));
KC_AOI21_X1 D2052 ( .B0(D8895_Q), .Y(D2052_Y), .A(D8939_Y),     .B1(D8883_Y));
KC_AOI21_X1 D2049 ( .B0(D326_Q), .Y(D2049_Y), .A(D2050_Y),     .B1(D8901_Y));
KC_AOI21_X1 D1909 ( .B0(D7360_Y), .Y(D1909_Y), .A(D7352_Y),     .B1(D7195_Y));
KC_AOI21_X1 D1903 ( .B0(D7319_Y), .Y(D1903_Y), .A(D2122_Y),     .B1(D4515_Y));
KC_AOI21_X1 D1901 ( .B0(D1859_Y), .Y(D1901_Y), .A(D1858_Y),     .B1(D7963_Y));
KC_AOI21_X1 D1896 ( .B0(D8087_Y), .Y(D1896_Y), .A(D8084_Y),     .B1(D9391_Y));
KC_AOI21_X1 D1894 ( .B0(D8406_Y), .Y(D1894_Y), .A(D6787_Y),     .B1(D8474_Y));
KC_AOI21_X1 D1893 ( .B0(D8240_Y), .Y(D1893_Y), .A(D8011_Y),     .B1(D3903_Y));
KC_AOI21_X1 D1888 ( .B0(D105_Y), .Y(D1888_Y), .A(D1966_Y),     .B1(D1827_Y));
KC_AOI21_X1 D1614 ( .B0(D4157_Y), .Y(D1614_Y), .A(D5867_Y),     .B1(D4358_Y));
KC_AOI21_X1 D1610 ( .B0(D4524_Y), .Y(D1610_Y), .A(D3243_Y),     .B1(D3030_Y));
KC_AOI21_X1 D1602 ( .B0(D3525_Y), .Y(D1602_Y), .A(D4910_Y),     .B1(D4911_Y));
KC_AOI21_X1 D1455 ( .B0(D9345_Y), .Y(D1455_Y), .A(D3098_Y),     .B1(D1428_Y));
KC_AOI21_X1 D1447 ( .B0(D3432_Y), .Y(D1447_Y), .A(D3551_Y),     .B1(D3526_Y));
KC_AOI21_X1 D1446 ( .B0(D3498_Y), .Y(D1446_Y), .A(D3406_Y),     .B1(D4960_Y));
KC_AOI21_X1 D1194 ( .B0(D7991_Y), .Y(D1194_Y), .A(D1936_Y),     .B1(D12071_Y));
KC_AOI21_X1 D1193 ( .B0(D7991_Y), .Y(D1193_Y), .A(D1936_Y),     .B1(D12004_Y));
KC_AOI21_X1 D1192 ( .B0(D14248_Y), .Y(D1192_Y), .A(D14070_Y),     .B1(D15684_Y));
KC_AOI21_X1 D1190 ( .B0(D14248_Y), .Y(D1190_Y), .A(D14071_Y),     .B1(D15113_Y));
KC_AOI21_X1 D1186 ( .B0(D8466_Y), .Y(D1186_Y), .A(D8502_Y),     .B1(D5547_Y));
KC_AOI21_X1 D1165 ( .B0(D14248_Y), .Y(D1165_Y), .A(D14073_Y),     .B1(D15691_Y));
KC_AOI21_X1 D1105 ( .B0(D14251_Y), .Y(D1105_Y), .A(D14073_Y),     .B1(D762_Y));
KC_AOI21_X1 D993 ( .B0(D8240_Y), .Y(D993_Y), .A(D8011_Y),     .B1(D5420_Y));
KC_AOI21_X1 D766 ( .B0(D10787_Y), .Y(D766_Y), .A(D10803_Y),     .B1(D11683_Y));
KC_AOI21_X1 D644 ( .B0(D14664_Y), .Y(D644_Y), .A(D16608_Y),     .B1(D13953_Y));
KC_AOI21_X1 D309 ( .B0(D1578_Y), .Y(D309_Y), .A(D4498_Y),     .B1(D4505_Y));
KC_AOI21_X1 D223 ( .B0(D7882_Y), .Y(D223_Y), .A(D201_Y), .B1(D8702_Y));
KC_AOI21_X1 D94 ( .B0(D5755_Y), .Y(D94_Y), .A(D1751_Y), .B1(D5746_Y));
KC_AOI21_X1 D91 ( .B0(D8240_Y), .Y(D91_Y), .A(D6772_Y), .B1(D5366_Y));
KC_OAI211_X1 D16518 ( .B(D16546_Y), .C0(D16547_Y), .A(D16523_Y),     .C1(D16624_Y), .Y(D16518_Y));
KC_OAI211_X1 D16123 ( .B(D16175_Y), .C0(D16124_Y), .A(D16104_Y),     .C1(D16124_Y), .Y(D16123_Y));
KC_OAI211_X1 D16069 ( .B(D16050_Y), .C0(D16051_Y), .A(D16060_Y),     .C1(D16059_Y), .Y(D16069_Y));
KC_OAI211_X1 D16004 ( .B(D16003_Y), .C0(D15228_Y), .A(D1339_Y),     .C1(D16003_Y), .Y(D16004_Y));
KC_OAI211_X1 D16002 ( .B(D15959_Y), .C0(D2471_Y), .A(D15982_Y),     .C1(D6406_Y), .Y(D16002_Y));
KC_OAI211_X1 D15981 ( .B(D15967_Y), .C0(D13610_Y), .A(D15978_Y),     .C1(D6406_Y), .Y(D15981_Y));
KC_OAI211_X1 D15974 ( .B(D15970_Y), .C0(D2471_Y), .A(D15977_Y),     .C1(D6410_Y), .Y(D15974_Y));
KC_OAI211_X1 D15973 ( .B(D15965_Y), .C0(D13641_Y), .A(D15984_Y),     .C1(D6406_Y), .Y(D15973_Y));
KC_OAI211_X1 D15972 ( .B(D15987_Y), .C0(D2421_Y), .A(D15976_Y),     .C1(D6406_Y), .Y(D15972_Y));
KC_OAI211_X1 D15928 ( .B(D15902_Y), .C0(D13641_Y), .A(D15852_Y),     .C1(D1813_Y), .Y(D15928_Y));
KC_OAI211_X1 D15926 ( .B(D15905_Y), .C0(D16767_Y), .A(D15929_Y),     .C1(D6410_Y), .Y(D15926_Y));
KC_OAI211_X1 D15925 ( .B(D15890_Y), .C0(D86_Y), .A(D15930_Y),     .C1(D6410_Y), .Y(D15925_Y));
KC_OAI211_X1 D15921 ( .B(D15878_Y), .C0(D13641_Y), .A(D15919_Y),     .C1(D6410_Y), .Y(D15921_Y));
KC_OAI211_X1 D15920 ( .B(D15090_Y), .C0(D13622_Y), .A(D15931_Y),     .C1(D6410_Y), .Y(D15920_Y));
KC_OAI211_X1 D15918 ( .B(D15914_Y), .C0(D13610_Y), .A(D15980_Y),     .C1(D6410_Y), .Y(D15918_Y));
KC_OAI211_X1 D15851 ( .B(D15906_Y), .C0(D16767_Y), .A(D15853_Y),     .C1(D1813_Y), .Y(D15851_Y));
KC_OAI211_X1 D15850 ( .B(D15907_Y), .C0(D13610_Y), .A(D15855_Y),     .C1(D1813_Y), .Y(D15850_Y));
KC_OAI211_X1 D15849 ( .B(D15824_Y), .C0(D13641_Y), .A(D15750_Y),     .C1(D813_Y), .Y(D15849_Y));
KC_OAI211_X1 D15848 ( .B(D15827_Y), .C0(D86_Y), .A(D2624_Y),     .C1(D813_Y), .Y(D15848_Y));
KC_OAI211_X1 D15847 ( .B(D15814_Y), .C0(D16767_Y), .A(D15841_Y),     .C1(D1814_Y), .Y(D15847_Y));
KC_OAI211_X1 D15846 ( .B(D15812_Y), .C0(D13641_Y), .A(D15843_Y),     .C1(D1814_Y), .Y(D15846_Y));
KC_OAI211_X1 D15844 ( .B(D15808_Y), .C0(D13610_Y), .A(D15840_Y),     .C1(D1814_Y), .Y(D15844_Y));
KC_OAI211_X1 D15837 ( .B(D15811_Y), .C0(D2471_Y), .A(D15839_Y),     .C1(D1813_Y), .Y(D15837_Y));
KC_OAI211_X1 D15836 ( .B(D15863_Y), .C0(D2471_Y), .A(D15842_Y),     .C1(D1814_Y), .Y(D15836_Y));
KC_OAI211_X1 D15773 ( .B(D15743_Y), .C0(D13641_Y), .A(D15771_Y),     .C1(D9617_Y), .Y(D15773_Y));
KC_OAI211_X1 D15770 ( .B(D15744_Y), .C0(D16767_Y), .A(D15767_Y),     .C1(D10358_Y), .Y(D15770_Y));
KC_OAI211_X1 D15769 ( .B(D987_Y), .C0(D2471_Y), .A(D15772_Y),     .C1(D10358_Y), .Y(D15769_Y));
KC_OAI211_X1 D15764 ( .B(D15724_Y), .C0(D13610_Y), .A(D15768_Y),     .C1(D9617_Y), .Y(D15764_Y));
KC_OAI211_X1 D15763 ( .B(D15741_Y), .C0(D13641_Y), .A(D15766_Y),     .C1(D10358_Y), .Y(D15763_Y));
KC_OAI211_X1 D15762 ( .B(D15727_Y), .C0(D86_Y), .A(D15760_Y),     .C1(D10358_Y), .Y(D15762_Y));
KC_OAI211_X1 D15758 ( .B(D15786_Y), .C0(D86_Y), .A(D15759_Y),     .C1(D9617_Y), .Y(D15758_Y));
KC_OAI211_X1 D15755 ( .B(D15716_Y), .C0(D13641_Y), .A(D15756_Y),     .C1(D8336_Y), .Y(D15755_Y));
KC_OAI211_X1 D15754 ( .B(D15723_Y), .C0(D16767_Y), .A(D15757_Y),     .C1(D8336_Y), .Y(D15754_Y));
KC_OAI211_X1 D15751 ( .B(D15721_Y), .C0(D13610_Y), .A(D15752_Y),     .C1(D8336_Y), .Y(D15751_Y));
KC_OAI211_X1 D15748 ( .B(D15713_Y), .C0(D86_Y), .A(D15753_Y),     .C1(D8336_Y), .Y(D15748_Y));
KC_OAI211_X1 D15746 ( .B(D15787_Y), .C0(D2471_Y), .A(D15747_Y),     .C1(D8336_Y), .Y(D15746_Y));
KC_OAI211_X1 D15709 ( .B(D15667_Y), .C0(D14862_Y), .A(D15708_Y),     .C1(D15478_Y), .Y(D15709_Y));
KC_OAI211_X1 D15662 ( .B(D15477_Y), .C0(D749_Y), .A(D15642_Y),     .C1(D15615_Y), .Y(D15662_Y));
KC_OAI211_X1 D15661 ( .B(D2635_Y), .C0(D15658_Y), .A(D15645_Y),     .C1(D2605_Y), .Y(D15661_Y));
KC_OAI211_X1 D15656 ( .B(D2634_Y), .C0(D14867_Y), .A(D15640_Y),     .C1(D15478_Y), .Y(D15656_Y));
KC_OAI211_X1 D15655 ( .B(D15705_Y), .C0(D14845_Y), .A(D15639_Y),     .C1(D2605_Y), .Y(D15655_Y));
KC_OAI211_X1 D15654 ( .B(D15625_Y), .C0(D15615_Y), .A(D15635_Y),     .C1(D15543_Y), .Y(D15654_Y));
KC_OAI211_X1 D15653 ( .B(D15666_Y), .C0(D15622_Y), .A(D15702_Y),     .C1(D15478_Y), .Y(D15653_Y));
KC_OAI211_X1 D15651 ( .B(D15638_Y), .C0(D15621_Y), .A(D15665_Y),     .C1(D15543_Y), .Y(D15651_Y));
KC_OAI211_X1 D15650 ( .B(D15631_Y), .C0(D15627_Y), .A(D873_Y),     .C1(D15543_Y), .Y(D15650_Y));
KC_OAI211_X1 D15649 ( .B(D878_Y), .C0(D15617_Y), .A(D15623_Y),     .C1(D15650_Y), .Y(D15649_Y));
KC_OAI211_X1 D15558 ( .B(D15565_Y), .C0(D15559_Y), .A(D15535_Y),     .C1(D15540_Y), .Y(D15558_Y));
KC_OAI211_X1 D15557 ( .B(D15446_Y), .C0(D771_Y), .A(D15400_Y),     .C1(D15537_Y), .Y(D15557_Y));
KC_OAI211_X1 D15556 ( .B(D15444_Y), .C0(D15527_Y), .A(D15399_Y),     .C1(D15540_Y), .Y(D15556_Y));
KC_OAI211_X1 D15553 ( .B(D15566_Y), .C0(D15554_Y), .A(D15601_Y),     .C1(D15537_Y), .Y(D15553_Y));
KC_OAI211_X1 D15552 ( .B(D15452_Y), .C0(D15512_Y), .A(D15604_Y),     .C1(D15537_Y), .Y(D15552_Y));
KC_OAI211_X1 D15548 ( .B(D15550_Y), .C0(D15516_Y), .A(D759_Y),     .C1(D15426_Y), .Y(D15548_Y));
KC_OAI211_X1 D15426 ( .B(D15342_Y), .C0(D15525_Y), .A(D15401_Y),     .C1(D15412_Y), .Y(D15426_Y));
KC_OAI211_X1 D15425 ( .B(D15403_Y), .C0(D15519_Y), .A(D15445_Y),     .C1(D15412_Y), .Y(D15425_Y));
KC_OAI211_X1 D15416 ( .B(D15369_Y), .C0(D636_Y), .A(D15358_Y),     .C1(D15518_Y), .Y(D15416_Y));
KC_OAI211_X1 D15411 ( .B(D15351_Y), .C0(D15518_Y), .A(D15360_Y),     .C1(D15412_Y), .Y(D15411_Y));
KC_OAI211_X1 D15204 ( .B(D1280_Y), .C0(D13641_Y), .A(D15206_Y),     .C1(D10191_Y), .Y(D15204_Y));
KC_OAI211_X1 D15202 ( .B(D15167_Y), .C0(D13622_Y), .A(D15120_Y),     .C1(D1964_Y), .Y(D15202_Y));
KC_OAI211_X1 D15199 ( .B(D15208_Y), .C0(D2420_Y), .A(D15200_Y),     .C1(D10191_Y), .Y(D15199_Y));
KC_OAI211_X1 D15198 ( .B(D15181_Y), .C0(D2471_Y), .A(D15190_Y),     .C1(D1964_Y), .Y(D15198_Y));
KC_OAI211_X1 D15196 ( .B(D14416_Y), .C0(D13641_Y), .A(D15207_Y),     .C1(D1964_Y), .Y(D15196_Y));
KC_OAI211_X1 D15195 ( .B(D15177_Y), .C0(D13610_Y), .A(D15193_Y),     .C1(D10191_Y), .Y(D15195_Y));
KC_OAI211_X1 D15191 ( .B(D14409_Y), .C0(D13610_Y), .A(D15192_Y),     .C1(D1964_Y), .Y(D15191_Y));
KC_OAI211_X1 D15188 ( .B(D14447_Y), .C0(D2471_Y), .A(D15189_Y),     .C1(D10191_Y), .Y(D15188_Y));
KC_OAI211_X1 D15187 ( .B(D15162_Y), .C0(D2421_Y), .A(D15201_Y),     .C1(D10191_Y), .Y(D15187_Y));
KC_OAI211_X1 D15184 ( .B(D15221_Y), .C0(D2420_Y), .A(D15186_Y),     .C1(D1964_Y), .Y(D15184_Y));
KC_OAI211_X1 D15183 ( .B(D14428_Y), .C0(D2421_Y), .A(D15185_Y),     .C1(D1964_Y), .Y(D15183_Y));
KC_OAI211_X1 D15117 ( .B(D1183_Y), .C0(D16767_Y), .A(D15119_Y),     .C1(D10191_Y), .Y(D15117_Y));
KC_OAI211_X1 D15116 ( .B(D15097_Y), .C0(D6406_Y), .A(D1192_Y),     .C1(D13619_Y), .Y(D15116_Y));
KC_OAI211_X1 D15062 ( .B(D15027_Y), .C0(D1814_Y), .A(D15064_Y),     .C1(D13619_Y), .Y(D15062_Y));
KC_OAI211_X1 D15059 ( .B(D15013_Y), .C0(D1813_Y), .A(D15060_Y),     .C1(D13619_Y), .Y(D15059_Y));
KC_OAI211_X1 D15058 ( .B(D15010_Y), .C0(D2487_Y), .A(D15057_Y),     .C1(D1813_Y), .Y(D15058_Y));
KC_OAI211_X1 D15056 ( .B(D15044_Y), .C0(D6410_Y), .A(D15066_Y),     .C1(D13619_Y), .Y(D15056_Y));
KC_OAI211_X1 D15053 ( .B(D15021_Y), .C0(D2487_Y), .A(D15054_Y),     .C1(D1814_Y), .Y(D15053_Y));
KC_OAI211_X1 D15050 ( .B(D15016_Y), .C0(D13622_Y), .A(D15051_Y),     .C1(D1813_Y), .Y(D15050_Y));
KC_OAI211_X1 D15049 ( .B(D15020_Y), .C0(D13622_Y), .A(D15052_Y),     .C1(D1814_Y), .Y(D15049_Y));
KC_OAI211_X1 D14972 ( .B(D14949_Y), .C0(D2487_Y), .A(D14225_Y),     .C1(D9617_Y), .Y(D14972_Y));
KC_OAI211_X1 D14970 ( .B(D14944_Y), .C0(D2487_Y), .A(D14973_Y),     .C1(D10358_Y), .Y(D14970_Y));
KC_OAI211_X1 D14967 ( .B(D14938_Y), .C0(D13622_Y), .A(D14974_Y),     .C1(D10358_Y), .Y(D14967_Y));
KC_OAI211_X1 D14966 ( .B(D14930_Y), .C0(D13622_Y), .A(D14971_Y),     .C1(D8336_Y), .Y(D14966_Y));
KC_OAI211_X1 D14963 ( .B(D2530_Y), .C0(D13622_Y), .A(D2555_Y),     .C1(D813_Y), .Y(D14963_Y));
KC_OAI211_X1 D14961 ( .B(D14939_Y), .C0(D2487_Y), .A(D14968_Y),     .C1(D8336_Y), .Y(D14961_Y));
KC_OAI211_X1 D14855 ( .B(D14816_Y), .C0(D8336_Y), .A(D2559_Y),     .C1(D13619_Y), .Y(D14855_Y));
KC_OAI211_X1 D14807 ( .B(D13935_Y), .C0(D2617_Y), .A(D15505_Y),     .C1(D14735_Y), .Y(D14807_Y));
KC_OAI211_X1 D14770 ( .B(D14733_Y), .C0(D14054_Y), .A(D14102_Y),     .C1(D1813_Y), .Y(D14770_Y));
KC_OAI211_X1 D14769 ( .B(D14740_Y), .C0(D14115_Y), .A(D839_Y),     .C1(D14727_Y), .Y(D14769_Y));
KC_OAI211_X1 D14768 ( .B(D14732_Y), .C0(D14054_Y), .A(D14101_Y),     .C1(D6410_Y), .Y(D14768_Y));
KC_OAI211_X1 D14767 ( .B(D14031_Y), .C0(D14115_Y), .A(D14098_Y),     .C1(D14011_Y), .Y(D14767_Y));
KC_OAI211_X1 D14766 ( .B(D14729_Y), .C0(D14054_Y), .A(D839_Y),     .C1(D10358_Y), .Y(D14766_Y));
KC_OAI211_X1 D14765 ( .B(D14739_Y), .C0(D14115_Y), .A(D838_Y),     .C1(D14726_Y), .Y(D14765_Y));
KC_OAI211_X1 D14764 ( .B(D14738_Y), .C0(D14115_Y), .A(D14101_Y),     .C1(D14809_Y), .Y(D14764_Y));
KC_OAI211_X1 D14763 ( .B(D14717_Y), .C0(D14054_Y), .A(D838_Y),     .C1(D8336_Y), .Y(D14763_Y));
KC_OAI211_X1 D14761 ( .B(D2540_Y), .C0(D14148_Y), .A(D14102_Y),     .C1(D1813_Y), .Y(D14761_Y));
KC_OAI211_X1 D14758 ( .B(D14723_Y), .C0(D2503_Y), .A(D14102_Y),     .C1(D1813_Y), .Y(D14758_Y));
KC_OAI211_X1 D14757 ( .B(D14722_Y), .C0(D2503_Y), .A(D839_Y),     .C1(D10358_Y), .Y(D14757_Y));
KC_OAI211_X1 D14756 ( .B(D14716_Y), .C0(D2503_Y), .A(D14101_Y),     .C1(D6410_Y), .Y(D14756_Y));
KC_OAI211_X1 D14755 ( .B(D14721_Y), .C0(D2503_Y), .A(D838_Y),     .C1(D8336_Y), .Y(D14755_Y));
KC_OAI211_X1 D14709 ( .B(D14678_Y), .C0(D14805_Y), .A(D14710_Y),     .C1(D15504_Y), .Y(D14709_Y));
KC_OAI211_X1 D14568 ( .B(D14595_Y), .C0(D14802_Y), .A(D14538_Y),     .C1(D12235_Q), .Y(D14568_Y));
KC_OAI211_X1 D14565 ( .B(D14566_Y), .C0(D14572_Y), .A(D14551_Y),     .C1(D14520_Q), .Y(D14565_Y));
KC_OAI211_X1 D14561 ( .B(D14593_Y), .C0(D14802_Y), .A(D14537_Y),     .C1(D12234_Q), .Y(D14561_Y));
KC_OAI211_X1 D14559 ( .B(D14598_Y), .C0(D14802_Y), .A(D14533_Y),     .C1(D12237_Q), .Y(D14559_Y));
KC_OAI211_X1 D14558 ( .B(D14554_Y), .C0(D14544_Y), .A(D14645_Y),     .C1(D14557_Y), .Y(D14558_Y));
KC_OAI211_X1 D14458 ( .B(D14450_Y), .C0(D2471_Y), .A(D14459_Y),     .C1(D10192_Y), .Y(D14458_Y));
KC_OAI211_X1 D14457 ( .B(D14402_Y), .C0(D2421_Y), .A(D13780_Y),     .C1(D10192_Y), .Y(D14457_Y));
KC_OAI211_X1 D14456 ( .B(D14398_Y), .C0(D2420_Y), .A(D14462_Y),     .C1(D10192_Y), .Y(D14456_Y));
KC_OAI211_X1 D14368 ( .B(D2480_Y), .C0(D10192_Y), .A(D1190_Y),     .C1(D13619_Y), .Y(D14368_Y));
KC_OAI211_X1 D14367 ( .B(D14330_Y), .C0(D16767_Y), .A(D2552_Y),     .C1(D1964_Y), .Y(D14367_Y));
KC_OAI211_X1 D14153 ( .B(D14178_Y), .C0(D14148_Y), .A(D14100_Y),     .C1(D1814_Y), .Y(D14153_Y));
KC_OAI211_X1 D14152 ( .B(D14012_Y), .C0(D2503_Y), .A(D14099_Y),     .C1(D9617_Y), .Y(D14152_Y));
KC_OAI211_X1 D14151 ( .B(D14140_Y), .C0(D14148_Y), .A(D14098_Y),     .C1(D813_Y), .Y(D14151_Y));
KC_OAI211_X1 D14150 ( .B(D14135_Y), .C0(D14148_Y), .A(D14099_Y),     .C1(D9617_Y), .Y(D14150_Y));
KC_OAI211_X1 D14116 ( .B(D14132_Y), .C0(D13313_Y), .A(D14029_Y),     .C1(D13321_Y), .Y(D14116_Y));
KC_OAI211_X1 D14056 ( .B(D14027_Y), .C0(D14115_Y), .A(D14099_Y),     .C1(D14016_Y), .Y(D14056_Y));
KC_OAI211_X1 D14055 ( .B(D14014_Y), .C0(D14054_Y), .A(D14098_Y),     .C1(D813_Y), .Y(D14055_Y));
KC_OAI211_X1 D14053 ( .B(D14007_Y), .C0(D14054_Y), .A(D14099_Y),     .C1(D9617_Y), .Y(D14053_Y));
KC_OAI211_X1 D14052 ( .B(D14015_Y), .C0(D14054_Y), .A(D14100_Y),     .C1(D1814_Y), .Y(D14052_Y));
KC_OAI211_X1 D14051 ( .B(D14028_Y), .C0(D14115_Y), .A(D14100_Y),     .C1(D14725_Y), .Y(D14051_Y));
KC_OAI211_X1 D14050 ( .B(D14137_Y), .C0(D13313_Y), .A(D14029_Y),     .C1(D13322_Y), .Y(D14050_Y));
KC_OAI211_X1 D14049 ( .B(D14013_Y), .C0(D2503_Y), .A(D14100_Y),     .C1(D1814_Y), .Y(D14049_Y));
KC_OAI211_X1 D14048 ( .B(D2497_Y), .C0(D2503_Y), .A(D14098_Y),     .C1(D813_Y), .Y(D14048_Y));
KC_OAI211_X1 D13967 ( .B(D13234_Y), .C0(D764_Y), .A(D13934_Y),     .C1(D13939_Y), .Y(D13967_Y));
KC_OAI211_X1 D13966 ( .B(D13969_Y), .C0(D13970_Y), .A(D13219_Y),     .C1(D13937_Y), .Y(D13966_Y));
KC_OAI211_X1 D13964 ( .B(D13234_Y), .C0(D15508_Y), .A(D13220_Y),     .C1(D13941_Y), .Y(D13964_Y));
KC_OAI211_X1 D13791 ( .B(D13795_Y), .C0(D2421_Y), .A(D13784_Y),     .C1(D463_Y), .Y(D13791_Y));
KC_OAI211_X1 D13790 ( .B(D13772_Y), .C0(D13641_Y), .A(D13781_Y),     .C1(D463_Y), .Y(D13790_Y));
KC_OAI211_X1 D13788 ( .B(D14429_Y), .C0(D2420_Y), .A(D13792_Y),     .C1(D463_Y), .Y(D13788_Y));
KC_OAI211_X1 D13785 ( .B(D13777_Y), .C0(D13610_Y), .A(D13786_Y),     .C1(D463_Y), .Y(D13785_Y));
KC_OAI211_X1 D13782 ( .B(D13773_Y), .C0(D2471_Y), .A(D13783_Y),     .C1(D463_Y), .Y(D13782_Y));
KC_OAI211_X1 D13743 ( .B(D13728_Y), .C0(D463_Y), .A(D13739_Y),     .C1(D13619_Y), .Y(D13743_Y));
KC_OAI211_X1 D13742 ( .B(D2412_Y), .C0(D462_Y), .A(D1165_Y),     .C1(D13619_Y), .Y(D13742_Y));
KC_OAI211_X1 D13737 ( .B(D13750_Y), .C0(D16767_Y), .A(D13740_Y),     .C1(D10192_Y), .Y(D13737_Y));
KC_OAI211_X1 D13735 ( .B(D13751_Y), .C0(D16767_Y), .A(D13732_Y),     .C1(D463_Y), .Y(D13735_Y));
KC_OAI211_X1 D13733 ( .B(D13713_Y), .C0(D13622_Y), .A(D13734_Y),     .C1(D10192_Y), .Y(D13733_Y));
KC_OAI211_X1 D13731 ( .B(D13714_Y), .C0(D13622_Y), .A(D13789_Y),     .C1(D463_Y), .Y(D13731_Y));
KC_OAI211_X1 D13712 ( .B(D13642_Y), .C0(D16767_Y), .A(D13675_Y),     .C1(D462_Y), .Y(D13712_Y));
KC_OAI211_X1 D13688 ( .B(D2399_Y), .C0(D13542_Y), .A(D13654_Y),     .C1(D13661_Y), .Y(D13688_Y));
KC_OAI211_X1 D13687 ( .B(D13630_Y), .C0(D13602_Y), .A(D13651_Y),     .C1(D13660_Y), .Y(D13687_Y));
KC_OAI211_X1 D13686 ( .B(D13708_Y), .C0(D13603_Y), .A(D13650_Y),     .C1(D13659_Y), .Y(D13686_Y));
KC_OAI211_X1 D13685 ( .B(D13647_Y), .C0(D13641_Y), .A(D13678_Y),     .C1(D462_Y), .Y(D13685_Y));
KC_OAI211_X1 D13684 ( .B(D13643_Y), .C0(D13622_Y), .A(D13676_Y),     .C1(D462_Y), .Y(D13684_Y));
KC_OAI211_X1 D13683 ( .B(D13701_Y), .C0(D2421_Y), .A(D13681_Y),     .C1(D462_Y), .Y(D13683_Y));
KC_OAI211_X1 D13682 ( .B(D1089_Y), .C0(D2420_Y), .A(D13680_Y),     .C1(D462_Y), .Y(D13682_Y));
KC_OAI211_X1 D13679 ( .B(D13648_Y), .C0(D2471_Y), .A(D13677_Y),     .C1(D462_Y), .Y(D13679_Y));
KC_OAI211_X1 D13674 ( .B(D13667_Y), .C0(D13610_Y), .A(D1105_Y),     .C1(D462_Y), .Y(D13674_Y));
KC_OAI211_X1 D13638 ( .B(D12956_Y), .C0(D13437_Y), .A(D13563_Y),     .C1(D13572_Y), .Y(D13638_Y));
KC_OAI211_X1 D13594 ( .B(D13576_Y), .C0(D13436_Y), .A(D13568_Y),     .C1(D13570_Y), .Y(D13594_Y));
KC_OAI211_X1 D13593 ( .B(D13004_Y), .C0(D13572_Y), .A(D13574_Y),     .C1(D13436_Y), .Y(D13593_Y));
KC_OAI211_X1 D13589 ( .B(D12953_Y), .C0(D13437_Y), .A(D13564_Y),     .C1(D13570_Y), .Y(D13589_Y));
KC_OAI211_X1 D13588 ( .B(D13393_Y), .C0(D13709_Y), .A(D13566_Y),     .C1(D12754_Q), .Y(D13588_Y));
KC_OAI211_X1 D13585 ( .B(D13543_Y), .C0(D13573_Y), .A(D2436_Y),     .C1(D13338_Y), .Y(D13585_Y));
KC_OAI211_X1 D13584 ( .B(D13548_Y), .C0(D170_Y), .A(D2436_Y),     .C1(D13338_Y), .Y(D13584_Y));
KC_OAI211_X1 D13583 ( .B(D13632_Y), .C0(D13619_Y), .A(D13425_Y),     .C1(D6407_Y), .Y(D13583_Y));
KC_OAI211_X1 D13537 ( .B(D13435_Y), .C0(D855_Q), .A(D966_Y),     .C1(D2395_Y), .Y(D13537_Y));
KC_OAI211_X1 D13533 ( .B(D13435_Y), .C0(D13515_Q), .A(D13534_Y),     .C1(D12861_Y), .Y(D13533_Y));
KC_OAI211_X1 D13500 ( .B(D13463_Y), .C0(D13436_Y), .A(D13433_Y),     .C1(D13479_Y), .Y(D13500_Y));
KC_OAI211_X1 D13495 ( .B(D13435_Y), .C0(D852_Q), .A(D13441_Y),     .C1(D2394_Y), .Y(D13495_Y));
KC_OAI211_X1 D13494 ( .B(D13453_Y), .C0(D13437_Y), .A(D13432_Y),     .C1(D13479_Y), .Y(D13494_Y));
KC_OAI211_X1 D13493 ( .B(D2438_Y), .C0(D13438_Y), .A(D2436_Y),     .C1(D13338_Y), .Y(D13493_Y));
KC_OAI211_X1 D13488 ( .B(D2436_Y), .C0(D13431_Y), .A(D13458_Y),     .C1(D13338_Y), .Y(D13488_Y));
KC_OAI211_X1 D13484 ( .B(D2435_Y), .C0(D13424_Y), .A(D2436_Y),     .C1(D13338_Y), .Y(D13484_Y));
KC_OAI211_X1 D13483 ( .B(D13426_Y), .C0(D13436_Y), .A(D13415_Y),     .C1(D13423_Y), .Y(D13483_Y));
KC_OAI211_X1 D13480 ( .B(D2424_Y), .C0(D13437_Y), .A(D2423_Y),     .C1(D13423_Y), .Y(D13480_Y));
KC_OAI211_X1 D13373 ( .B(D13385_Y), .C0(D12718_Y), .A(D13355_Y),     .C1(D12732_Y), .Y(D13373_Y));
KC_OAI211_X1 D13026 ( .B(D13053_Y), .C0(D2370_Y), .A(D13657_Y),     .C1(D2369_Y), .Y(D13026_Y));
KC_OAI211_X1 D13025 ( .B(D13000_Y), .C0(D13019_Y), .A(D13653_Y),     .C1(D13018_Y), .Y(D13025_Y));
KC_OAI211_X1 D12966 ( .B(D13435_Y), .C0(D12926_Q), .A(D13539_Y),     .C1(D12928_Y), .Y(D12966_Y));
KC_OAI211_X1 D12962 ( .B(D13435_Y), .C0(D12931_Y), .A(D13553_Y),     .C1(D814_Q), .Y(D12962_Y));
KC_OAI211_X1 D12961 ( .B(D13435_Y), .C0(D956_Q), .A(D13552_Y),     .C1(D12930_Y), .Y(D12961_Y));
KC_OAI211_X1 D12864 ( .B(D12794_Y), .C0(D783_Y), .A(D12865_Y),     .C1(D12855_Q), .Y(D12864_Y));
KC_OAI211_X1 D12765 ( .B(D13234_Y), .C0(D12718_Y), .A(D12736_Y),     .C1(D13268_Q), .Y(D12765_Y));
KC_OAI211_X1 D12728 ( .B(D12693_Y), .C0(D12719_Y), .A(D12706_Y),     .C1(D12729_Y), .Y(D12728_Y));
KC_OAI211_X1 D12242 ( .B(D12189_Y), .C0(D12196_Y), .A(D12243_Y),     .C1(D12212_Y), .Y(D12242_Y));
KC_OAI211_X1 D10519 ( .B(D10509_Q), .C0(D10407_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D10519_Y));
KC_OAI211_X1 D10491 ( .B(D10518_Y), .C0(D9746_Y), .A(D10487_Y),     .C1(D10408_Y), .Y(D10491_Y));
KC_OAI211_X1 D10490 ( .B(D10410_Y), .C0(D10407_Y), .A(D10489_Y),     .C1(D9746_Y), .Y(D10490_Y));
KC_OAI211_X1 D10489 ( .B(D10513_Q), .C0(D10408_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D10489_Y));
KC_OAI211_X1 D10488 ( .B(D1919_Y), .C0(D10994_Q), .A(D10465_Y),     .C1(D10505_Y), .Y(D10488_Y));
KC_OAI211_X1 D10484 ( .B(D9785_Q), .C0(D10455_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D10484_Y));
KC_OAI211_X1 D10482 ( .B(D10409_Y), .C0(D10388_Y), .A(D10519_Y),     .C1(D9746_Y), .Y(D10482_Y));
KC_OAI211_X1 D10481 ( .B(D1127_Q), .C0(D10389_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D10481_Y));
KC_OAI211_X1 D10480 ( .B(D2140_Y), .C0(D10389_Y), .A(D2138_Y),     .C1(D9746_Y), .Y(D10480_Y));
KC_OAI211_X1 D10477 ( .B(D10483_Y), .C0(D10453_Y), .A(D10476_Y),     .C1(D9746_Y), .Y(D10477_Y));
KC_OAI211_X1 D10476 ( .B(D1123_Q), .C0(D10454_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D10476_Y));
KC_OAI211_X1 D10475 ( .B(D116_Q), .C0(D10446_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D10475_Y));
KC_OAI211_X1 D10474 ( .B(D2157_Q), .C0(D10453_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D10474_Y));
KC_OAI211_X1 D10472 ( .B(D10478_Y), .C0(D10446_Y), .A(D10474_Y),     .C1(D9746_Y), .Y(D10472_Y));
KC_OAI211_X1 D10314 ( .B(D10252_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D10299_Q), .Y(D10314_Y));
KC_OAI211_X1 D10312 ( .B(D10251_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D10301_Q), .Y(D10312_Y));
KC_OAI211_X1 D10265 ( .B(D9428_Y), .C0(D2862_Y), .A(D2136_Y),     .C1(D10232_Y), .Y(D10265_Y));
KC_OAI211_X1 D10264 ( .B(D9428_Y), .C0(D774_Y), .A(D10258_Y),     .C1(D848_Y), .Y(D10264_Y));
KC_OAI211_X1 D10263 ( .B(D10255_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D10294_Q), .Y(D10263_Y));
KC_OAI211_X1 D10262 ( .B(D10254_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D10311_Q), .Y(D10262_Y));
KC_OAI211_X1 D10261 ( .B(D10250_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D10303_Q), .Y(D10261_Y));
KC_OAI211_X1 D10260 ( .B(D10249_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D10302_Q), .Y(D10260_Y));
KC_OAI211_X1 D10259 ( .B(D10256_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D825_Q), .Y(D10259_Y));
KC_OAI211_X1 D10238 ( .B(D10199_Y), .C0(D9414_Y), .A(D9483_Y),     .C1(D9530_Y), .Y(D10238_Y));
KC_OAI211_X1 D10237 ( .B(D10230_Y), .C0(D9424_Y), .A(D9483_Y),     .C1(D9530_Y), .Y(D10237_Y));
KC_OAI211_X1 D10236 ( .B(D10257_Y), .C0(D9406_Y), .A(D9483_Y),     .C1(D9530_Y), .Y(D10236_Y));
KC_OAI211_X1 D10203 ( .B(D2169_Y), .C0(D10196_Y), .A(D9483_Y),     .C1(D9530_Y), .Y(D10203_Y));
KC_OAI211_X1 D10202 ( .B(D10198_Y), .C0(D9415_Y), .A(D9483_Y),     .C1(D9530_Y), .Y(D10202_Y));
KC_OAI211_X1 D10092 ( .B(D5966_Y), .C0(D11623_Y), .A(D11114_Y),     .C1(D10629_Y), .Y(D10092_Y));
KC_OAI211_X1 D10042 ( .B(D8878_Y), .C0(D10039_Y), .A(D2017_Y),     .C1(D7407_Y), .Y(D10042_Y));
KC_OAI211_X1 D10041 ( .B(D10036_Y), .C0(D7407_Y), .A(D10046_Y),     .C1(D9016_Y), .Y(D10041_Y));
KC_OAI211_X1 D10040 ( .B(D2049_Y), .C0(D7407_Y), .A(D279_Y),     .C1(D10044_Y), .Y(D10040_Y));
KC_OAI211_X1 D10025 ( .B(D10015_Y), .C0(D7407_Y), .A(D10030_Y),     .C1(D8950_Y), .Y(D10025_Y));
KC_OAI211_X1 D10024 ( .B(D8932_Y), .C0(D7407_Y), .A(D10018_Y),     .C1(D9017_Y), .Y(D10024_Y));
KC_OAI211_X1 D10023 ( .B(D10010_Y), .C0(D10027_Y), .A(D10012_Y),     .C1(D242_Y), .Y(D10023_Y));
KC_OAI211_X1 D10022 ( .B(D10013_Y), .C0(D7407_Y), .A(D2163_Y),     .C1(D9013_Y), .Y(D10022_Y));
KC_OAI211_X1 D10004 ( .B(D9993_Y), .C0(D10027_Y), .A(D250_Y),     .C1(D9996_Y), .Y(D10004_Y));
KC_OAI211_X1 D10003 ( .B(D9988_Y), .C0(D10028_Y), .A(D9997_Y),     .C1(D9996_Y), .Y(D10003_Y));
KC_OAI211_X1 D9797 ( .B(D9790_Q), .C0(D9738_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D9797_Y));
KC_OAI211_X1 D9796 ( .B(D9756_Y), .C0(D9743_Y), .A(D9764_Y),     .C1(D8550_Y), .Y(D9796_Y));
KC_OAI211_X1 D9769 ( .B(D9839_Q), .C0(D1978_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D9769_Y));
KC_OAI211_X1 D9768 ( .B(D9789_Q), .C0(D9728_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D9768_Y));
KC_OAI211_X1 D9767 ( .B(D2033_Y), .C0(D9737_Y), .A(D1166_Y),     .C1(D8550_Y), .Y(D9767_Y));
KC_OAI211_X1 D9766 ( .B(D2079_Q), .C0(D9648_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D9766_Y));
KC_OAI211_X1 D9765 ( .B(D9793_Q), .C0(D9735_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D9765_Y));
KC_OAI211_X1 D9764 ( .B(D1131_Q), .C0(D9737_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D9764_Y));
KC_OAI211_X1 D9763 ( .B(D9759_Y), .C0(D9739_Y), .A(D9760_Y),     .C1(D9746_Y), .Y(D9763_Y));
KC_OAI211_X1 D9762 ( .B(D9758_Y), .C0(D9738_Y), .A(D9761_Y),     .C1(D9746_Y), .Y(D9762_Y));
KC_OAI211_X1 D9761 ( .B(D9792_Q), .C0(D9739_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D9761_Y));
KC_OAI211_X1 D9760 ( .B(D9791_Q), .C0(D9743_Y), .A(D8534_Y),     .C1(D8363_Y), .Y(D9760_Y));
KC_OAI211_X1 D9757 ( .B(D9753_Y), .C0(D9735_Y), .A(D9797_Y),     .C1(D8550_Y), .Y(D9757_Y));
KC_OAI211_X1 D9724 ( .B(D9786_Q), .C0(D9646_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D9724_Y));
KC_OAI211_X1 D9723 ( .B(D9689_Y), .C0(D9644_Y), .A(D2036_Y),     .C1(D9746_Y), .Y(D9723_Y));
KC_OAI211_X1 D9686 ( .B(D9691_Y), .C0(D9647_Y), .A(D9724_Y),     .C1(D9746_Y), .Y(D9686_Y));
KC_OAI211_X1 D9685 ( .B(D9690_Y), .C0(D9646_Y), .A(D2111_Y),     .C1(D9746_Y), .Y(D9685_Y));
KC_OAI211_X1 D9684 ( .B(D9704_Q), .C0(D9644_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D9684_Y));
KC_OAI211_X1 D9548 ( .B(D9572_Y), .C0(D9219_Q), .A(D9571_Y),     .C1(D9597_Y), .Y(D9548_Y));
KC_OAI211_X1 D9438 ( .B(D8137_Y), .C0(D9417_Y), .A(D9412_Y),     .C1(D9486_Y), .Y(D9438_Y));
KC_OAI211_X1 D9433 ( .B(D2116_Y), .C0(D9422_Y), .A(D9483_Y),     .C1(D9530_Y), .Y(D9433_Y));
KC_OAI211_X1 D9430 ( .B(D9397_Y), .C0(D622_Y), .A(D8086_Y),     .C1(D9402_Y), .Y(D9430_Y));
KC_OAI211_X1 D9429 ( .B(D10245_Y), .C0(D9423_Y), .A(D9483_Y),     .C1(D9530_Y), .Y(D9429_Y));
KC_OAI211_X1 D9427 ( .B(D8156_Y), .C0(D9401_Y), .A(D9392_Y),     .C1(D9582_Q), .Y(D9427_Y));
KC_OAI211_X1 D9202 ( .B(D9183_Y), .C0(D9186_Y), .A(D9305_Y),     .C1(D9108_Y), .Y(D9202_Y));
KC_OAI211_X1 D9198 ( .B(D9304_Y), .C0(D7680_Y), .A(D9307_Y),     .C1(D9186_Y), .Y(D9198_Y));
KC_OAI211_X1 D9127 ( .B(D9152_Y), .C0(D9108_Y), .A(D9100_Y),     .C1(D9147_Y), .Y(D9127_Y));
KC_OAI211_X1 D9083 ( .B(D7539_Y), .C0(D7510_Y), .A(D9037_Y),     .C1(D9056_Y), .Y(D9083_Y));
KC_OAI211_X1 D9082 ( .B(D9094_Y), .C0(D9017_Y), .A(D9043_Y),     .C1(D5703_Y), .Y(D9082_Y));
KC_OAI211_X1 D9080 ( .B(D382_Y), .C0(D5704_Y), .A(D354_Q),     .C1(D9109_Y), .Y(D9080_Y));
KC_OAI211_X1 D9078 ( .B(D382_Y), .C0(D5704_Y), .A(D10058_Q),     .C1(D9122_Y), .Y(D9078_Y));
KC_OAI211_X1 D8993 ( .B(D8984_Y), .C0(D9109_Y), .A(D9031_Y),     .C1(D7510_Y), .Y(D8993_Y));
KC_OAI211_X1 D8940 ( .B(D8936_Y), .C0(D8851_Y), .A(D8854_Y),     .C1(D8949_Y), .Y(D8940_Y));
KC_OAI211_X1 D8929 ( .B(D7458_Y), .C0(D2086_Y), .A(D8967_Y),     .C1(D8980_Y), .Y(D8929_Y));
KC_OAI211_X1 D8884 ( .B(D8879_Y), .C0(D10027_Y), .A(D8905_Y),     .C1(D7407_Y), .Y(D8884_Y));
KC_OAI211_X1 D8880 ( .B(D2052_Y), .C0(D8851_Y), .A(D8855_Y),     .C1(D8950_Y), .Y(D8880_Y));
KC_OAI211_X1 D8777 ( .B(D9476_Y), .C0(D8876_Y), .A(D9480_Y),     .C1(D8747_Y), .Y(D8777_Y));
KC_OAI211_X1 D8682 ( .B(D8770_Y), .C0(D8746_Y), .A(D8668_Y),     .C1(D8667_Y), .Y(D8682_Y));
KC_OAI211_X1 D8681 ( .B(D205_Y), .C0(D9941_Q), .A(D9923_Y),     .C1(D175_Y), .Y(D8681_Y));
KC_OAI211_X1 D8566 ( .B(D8568_Y), .C0(D8559_Y), .A(D8518_Y),     .C1(D8550_Y), .Y(D8566_Y));
KC_OAI211_X1 D8521 ( .B(D8547_Q), .C0(D8487_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D8521_Y));
KC_OAI211_X1 D8520 ( .B(D8549_Q), .C0(D8485_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D8520_Y));
KC_OAI211_X1 D8519 ( .B(D8595_Q), .C0(D8559_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D8519_Y));
KC_OAI211_X1 D8518 ( .B(D8539_Q), .C0(D8484_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D8518_Y));
KC_OAI211_X1 D8516 ( .B(D8517_Y), .C0(D8421_Y), .A(D8512_Y),     .C1(D8550_Y), .Y(D8516_Y));
KC_OAI211_X1 D8515 ( .B(D8543_Q), .C0(D9683_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D8515_Y));
KC_OAI211_X1 D8514 ( .B(D8513_Y), .C0(D9683_Y), .A(D1889_Y),     .C1(D8550_Y), .Y(D8514_Y));
KC_OAI211_X1 D8512 ( .B(D8544_Q), .C0(D8420_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D8512_Y));
KC_OAI211_X1 D8509 ( .B(D8510_Y), .C0(D8487_Y), .A(D8520_Y),     .C1(D8550_Y), .Y(D8509_Y));
KC_OAI211_X1 D8506 ( .B(D8508_Y), .C0(D8484_Y), .A(D8521_Y),     .C1(D8550_Y), .Y(D8506_Y));
KC_OAI211_X1 D8438 ( .B(D8475_Y), .C0(D1914_S), .A(D7928_Y),     .C1(D8387_Y), .Y(D8438_Y));
KC_OAI211_X1 D8437 ( .B(D7928_Y), .C0(D8397_Y), .A(D8412_Y),     .C1(D8457_Y), .Y(D8437_Y));
KC_OAI211_X1 D8436 ( .B(D1837_Y), .C0(D8419_Y), .A(D8388_Y),     .C1(D8369_Y), .Y(D8436_Y));
KC_OAI211_X1 D8435 ( .B(D8436_Y), .C0(D8386_Y), .A(D8406_Y),     .C1(D8388_Y), .Y(D8435_Y));
KC_OAI211_X1 D8434 ( .B(D7928_Y), .C0(D8376_Y), .A(D8385_Y),     .C1(D8435_Y), .Y(D8434_Y));
KC_OAI211_X1 D8429 ( .B(D1928_Q), .C0(D6864_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D8429_Y));
KC_OAI211_X1 D8428 ( .B(D8534_Y), .C0(D8421_Y), .A(D8545_Q),     .C1(D8542_Y), .Y(D8428_Y));
KC_OAI211_X1 D8427 ( .B(D8458_Q), .C0(D9647_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D8427_Y));
KC_OAI211_X1 D7904 ( .B(D7877_Y), .C0(D1855_Y), .A(D7905_Y),     .C1(D7888_Q), .Y(D7904_Y));
KC_OAI211_X1 D7868 ( .B(D7834_Y), .C0(D469_Y), .A(D1744_Y),     .C1(D7858_Y), .Y(D7868_Y));
KC_OAI211_X1 D7863 ( .B(D7864_Y), .C0(D7831_Y), .A(D7953_Y),     .C1(D7888_Q), .Y(D7863_Y));
KC_OAI211_X1 D7695 ( .B(D9180_Y), .C0(D7620_Y), .A(D9164_Y),     .C1(D7684_Y), .Y(D7695_Y));
KC_OAI211_X1 D7694 ( .B(D9175_Y), .C0(D7620_Y), .A(D9164_Y),     .C1(D9115_Y), .Y(D7694_Y));
KC_OAI211_X1 D7646 ( .B(D9130_Y), .C0(D9146_Y), .A(D9125_Y),     .C1(D9151_Y), .Y(D7646_Y));
KC_OAI211_X1 D7511 ( .B(D2009_Y), .C0(D282_Y), .A(D7493_Y),     .C1(D7510_Y), .Y(D7511_Y));
KC_OAI211_X1 D7448 ( .B(D8853_Y), .C0(D1867_Y), .A(D278_Y),     .C1(D7361_Y), .Y(D7448_Y));
KC_OAI211_X1 D7410 ( .B(D7364_Y), .C0(D4434_Y), .A(D7411_Y),     .C1(D10057_Y), .Y(D7410_Y));
KC_OAI211_X1 D7408 ( .B(D7332_Y), .C0(D7328_Y), .A(D75_Y),     .C1(D7538_Y), .Y(D7408_Y));
KC_OAI211_X1 D7379 ( .B(D1881_Y), .C0(D287_Y), .A(D1969_Y),     .C1(D7346_Y), .Y(D7379_Y));
KC_OAI211_X1 D7378 ( .B(D7100_Y), .C0(D2892_Y), .A(D7357_Y),     .C1(D7359_Y), .Y(D7378_Y));
KC_OAI211_X1 D7373 ( .B(D5866_Y), .C0(D7338_Y), .A(D7364_Y),     .C1(D5857_Y), .Y(D7373_Y));
KC_OAI211_X1 D7369 ( .B(D7328_Y), .C0(D214_Y), .A(D75_Y), .C1(D1581_Y),     .Y(D7369_Y));
KC_OAI211_X1 D7363 ( .B(D7365_Y), .C0(D6027_Y), .A(D7143_Y),     .C1(D6038_Y), .Y(D7363_Y));
KC_OAI211_X1 D7278 ( .B(D5804_Y), .C0(D7245_Y), .A(D7170_Y),     .C1(D7267_Y), .Y(D7278_Y));
KC_OAI211_X1 D7277 ( .B(D7261_Y), .C0(D7163_Y), .A(D7259_Y),     .C1(D7260_Y), .Y(D7277_Y));
KC_OAI211_X1 D7275 ( .B(D7238_Y), .C0(D202_Y), .A(D7237_Y),     .C1(D8756_Y), .Y(D7275_Y));
KC_OAI211_X1 D7272 ( .B(D4199_Y), .C0(D7306_Y), .A(D7223_Y),     .C1(D7376_Y), .Y(D7272_Y));
KC_OAI211_X1 D7270 ( .B(D7271_Y), .C0(D5703_Y), .A(D76_Y),     .C1(D5866_Y), .Y(D7270_Y));
KC_OAI211_X1 D7269 ( .B(D2053_Y), .C0(D8877_Y), .A(D234_Y),     .C1(D8776_Y), .Y(D7269_Y));
KC_OAI211_X1 D7265 ( .B(D7215_Y), .C0(D8744_Y), .A(D7182_Y),     .C1(D7268_Y), .Y(D7265_Y));
KC_OAI211_X1 D7122 ( .B(D7289_Y), .C0(D7096_Y), .A(D7259_Y),     .C1(D7099_Y), .Y(D7122_Y));
KC_OAI211_X1 D7121 ( .B(D7278_Y), .C0(D7096_Y), .A(D7105_Y),     .C1(D7107_Y), .Y(D7121_Y));
KC_OAI211_X1 D6879 ( .B(D6842_Y), .C0(D6843_Y), .A(D6842_Y),     .C1(D8371_Y), .Y(D6879_Y));
KC_OAI211_X1 D6458 ( .B(D477_Y), .C0(D1564_Y), .A(D5073_Y),     .C1(D6446_Y), .Y(D6458_Y));
KC_OAI211_X1 D6454 ( .B(D5071_Y), .C0(D5031_Y), .A(D6455_Y),     .C1(D4865_Y), .Y(D6454_Y));
KC_OAI211_X1 D6313 ( .B(D428_Y), .C0(D6294_Y), .A(D6312_Y),     .C1(D6340_Y), .Y(D6313_Y));
KC_OAI211_X1 D6310 ( .B(D6289_Y), .C0(D3325_Y), .A(D4655_Y),     .C1(D4682_Y), .Y(D6310_Y));
KC_OAI211_X1 D6309 ( .B(D4659_Y), .C0(D3325_Y), .A(D400_Y),     .C1(D4666_Y), .Y(D6309_Y));
KC_OAI211_X1 D6237 ( .B(D6241_Y), .C0(D9264_Y), .A(D6249_Y),     .C1(D6220_Y), .Y(D6237_Y));
KC_OAI211_X1 D6161 ( .B(D6168_Y), .C0(D6172_Y), .A(D6205_Y),     .C1(D6166_Y), .Y(D6161_Y));
KC_OAI211_X1 D6156 ( .B(D6159_Y), .C0(D6155_Y), .A(D6155_Y),     .C1(D6181_Y), .Y(D6156_Y));
KC_OAI211_X1 D6056 ( .B(D6004_Y), .C0(D5641_Y), .A(D6049_Y),     .C1(D6020_Y), .Y(D6056_Y));
KC_OAI211_X1 D6055 ( .B(D5996_Y), .C0(D6016_Y), .A(D6022_Y),     .C1(D214_Y), .Y(D6055_Y));
KC_OAI211_X1 D6041 ( .B(D8313_Q), .C0(D4409_Y), .A(D4149_Q),     .C1(D165_Y), .Y(D6041_Y));
KC_OAI211_X1 D5919 ( .B(D5879_Y), .C0(D5888_Y), .A(D1909_Y),     .C1(D5944_Y), .Y(D5919_Y));
KC_OAI211_X1 D5914 ( .B(D7351_Y), .C0(D4284_Y), .A(D5912_Y),     .C1(D5859_Y), .Y(D5914_Y));
KC_OAI211_X1 D5910 ( .B(D7372_Y), .C0(D5830_Y), .A(D7100_Y),     .C1(D4295_Y), .Y(D5910_Y));
KC_OAI211_X1 D5906 ( .B(D5948_Y), .C0(D213_Y), .A(D5898_Y),     .C1(D5925_Y), .Y(D5906_Y));
KC_OAI211_X1 D5901 ( .B(D5832_Y), .C0(D5905_Y), .A(D5831_Y),     .C1(D5852_Y), .Y(D5901_Y));
KC_OAI211_X1 D5900 ( .B(D5672_Y), .C0(D1872_Y), .A(D7391_Q),     .C1(D1739_Y), .Y(D5900_Y));
KC_OAI211_X1 D5897 ( .B(D5830_Y), .C0(D6030_Y), .A(D5900_Y),     .C1(D726_Y), .Y(D5897_Y));
KC_OAI211_X1 D5896 ( .B(D7329_Y), .C0(D4447_Y), .A(D213_Y),     .C1(D5763_Y), .Y(D5896_Y));
KC_OAI211_X1 D5895 ( .B(D7371_Y), .C0(D5763_Y), .A(D1585_Y),     .C1(D1735_Y), .Y(D5895_Y));
KC_OAI211_X1 D5790 ( .B(D5723_Y), .C0(D7294_Y), .A(D5770_Y),     .C1(D7211_Y), .Y(D5790_Y));
KC_OAI211_X1 D5784 ( .B(D5739_Y), .C0(D5734_Y), .A(D5740_Y),     .C1(D7376_Y), .Y(D5784_Y));
KC_OAI211_X1 D5781 ( .B(D7262_Y), .C0(D5912_Y), .A(D5818_Y),     .C1(D5866_Y), .Y(D5781_Y));
KC_OAI211_X1 D5780 ( .B(D210_Y), .C0(D5876_Y), .A(D5884_Y),     .C1(D5729_Y), .Y(D5780_Y));
KC_OAI211_X1 D5774 ( .B(D5942_Y), .C0(D5825_Y), .A(D5711_Y),     .C1(D5693_Q), .Y(D5774_Y));
KC_OAI211_X1 D5094 ( .B(D470_Y), .C0(D5003_Y), .A(D5095_Y),     .C1(D5023_Y), .Y(D5094_Y));
KC_OAI211_X1 D5064 ( .B(D5062_Y), .C0(D4912_Y), .A(D4997_Y),     .C1(D5044_Y), .Y(D5064_Y));
KC_OAI211_X1 D5063 ( .B(D5025_Y), .C0(D4925_Y), .A(D5070_Y),     .C1(D3530_Y), .Y(D5063_Y));
KC_OAI211_X1 D5056 ( .B(D5005_Y), .C0(D3371_Y), .A(D4881_Y),     .C1(D1565_Y), .Y(D5056_Y));
KC_OAI211_X1 D5055 ( .B(D5066_Y), .C0(D4865_Y), .A(D5007_Y),     .C1(D4880_Y), .Y(D5055_Y));
KC_OAI211_X1 D5049 ( .B(D5077_Y), .C0(D1564_Y), .A(D4997_Y),     .C1(D3498_Y), .Y(D5049_Y));
KC_OAI211_X1 D5048 ( .B(D5047_Y), .C0(D4865_Y), .A(D5054_Y),     .C1(D4999_Y), .Y(D5048_Y));
KC_OAI211_X1 D4947 ( .B(D4960_Y), .C0(D1605_Y), .A(D4926_Y),     .C1(D4890_Y), .Y(D4947_Y));
KC_OAI211_X1 D4942 ( .B(D4956_Y), .C0(D4923_Y), .A(D4974_Y),     .C1(D4959_Y), .Y(D4942_Y));
KC_OAI211_X1 D4939 ( .B(D5018_Y), .C0(D4915_Y), .A(D4936_Y),     .C1(D4904_Y), .Y(D4939_Y));
KC_OAI211_X1 D4928 ( .B(D3599_Y), .C0(D4875_Y), .A(D4874_Y),     .C1(D4913_Y), .Y(D4928_Y));
KC_OAI211_X1 D4927 ( .B(D4878_Y), .C0(D3470_Y), .A(D5034_Y),     .C1(D4860_Y), .Y(D4927_Y));
KC_OAI211_X1 D4786 ( .B(D4697_Y), .C0(D4767_Y), .A(D4760_Y),     .C1(D3325_Y), .Y(D4786_Y));
KC_OAI211_X1 D4784 ( .B(D4755_Y), .C0(D2086_Y), .A(D4655_Y),     .C1(D3325_Y), .Y(D4784_Y));
KC_OAI211_X1 D4782 ( .B(D4949_Y), .C0(D4805_Y), .A(D1569_Y),     .C1(D4750_Y), .Y(D4782_Y));
KC_OAI211_X1 D4738 ( .B(D4689_Y), .C0(D4693_Y), .A(D4739_Y),     .C1(D4580_Y), .Y(D4738_Y));
KC_OAI211_X1 D4708 ( .B(D4694_Y), .C0(D4695_Y), .A(D4638_Q),     .C1(D4575_Y), .Y(D4708_Y));
KC_OAI211_X1 D4707 ( .B(D4578_Y), .C0(D4572_Y), .A(D4638_Q),     .C1(D3097_Y), .Y(D4707_Y));
KC_OAI211_X1 D4704 ( .B(D4685_Y), .C0(D1622_Y), .A(D3294_Y),     .C1(D4731_Y), .Y(D4704_Y));
KC_OAI211_X1 D4615 ( .B(D4605_Y), .C0(D4504_Y), .A(D4520_Y),     .C1(D4622_Y), .Y(D4615_Y));
KC_OAI211_X1 D4458 ( .B(D5834_Y), .C0(D4280_Y), .A(D7311_Y),     .C1(D1581_Y), .Y(D4458_Y));
KC_OAI211_X1 D4378 ( .B(D1587_Y), .C0(D4323_Y), .A(D4344_Y),     .C1(D4436_Y), .Y(D4378_Y));
KC_OAI211_X1 D4375 ( .B(D4334_Y), .C0(D5868_Y), .A(D4346_Y),     .C1(D1592_Y), .Y(D4375_Y));
KC_OAI211_X1 D4370 ( .B(D4383_Y), .C0(D4315_Y), .A(D5793_Y),     .C1(D4349_Y), .Y(D4370_Y));
KC_OAI211_X1 D4269 ( .B(D4182_Y), .C0(D1722_Y), .A(D5751_Y),     .C1(D4294_Y), .Y(D4269_Y));
KC_OAI211_X1 D4223 ( .B(D4161_Y), .C0(D5766_Y), .A(D5765_Y),     .C1(D7376_Y), .Y(D4223_Y));
KC_OAI211_X1 D4220 ( .B(D4153_Y), .C0(D4374_Y), .A(D4344_Y),     .C1(D5649_Y), .Y(D4220_Y));
KC_OAI211_X1 D4218 ( .B(D4160_Y), .C0(D1722_Y), .A(D5751_Y),     .C1(D4421_Y), .Y(D4218_Y));
KC_OAI211_X1 D4215 ( .B(D4181_Y), .C0(D4374_Y), .A(D4352_Y),     .C1(D4173_Y), .Y(D4215_Y));
KC_OAI211_X1 D4214 ( .B(D1670_Y), .C0(D4304_Y), .A(D4175_Y),     .C1(D1589_Y), .Y(D4214_Y));
KC_OAI211_X1 D4213 ( .B(D4184_Y), .C0(D1732_Y), .A(D7221_Y),     .C1(D1629_Y), .Y(D4213_Y));
KC_OAI211_X1 D4209 ( .B(D5759_Y), .C0(D4219_Y), .A(D4155_Y),     .C1(D235_Y), .Y(D4209_Y));
KC_OAI211_X1 D3551 ( .B(D3539_Y), .C0(D3538_Y), .A(D3401_Y),     .C1(D3576_Q), .Y(D3551_Y));
KC_OAI211_X1 D3550 ( .B(D3536_Y), .C0(D4925_Y), .A(D4915_Y),     .C1(D3576_Q), .Y(D3550_Y));
KC_OAI211_X1 D3549 ( .B(D4881_Y), .C0(D3538_Y), .A(D3535_Y),     .C1(D3499_Y), .Y(D3549_Y));
KC_OAI211_X1 D3547 ( .B(D1450_Y), .C0(D3519_Y), .A(D3541_Y),     .C1(D3423_Y), .Y(D3547_Y));
KC_OAI211_X1 D3491 ( .B(D4977_Y), .C0(D3494_Y), .A(D3492_Y),     .C1(D3484_Q), .Y(D3491_Y));
KC_OAI211_X1 D3468 ( .B(D3445_Y), .C0(D3416_Y), .A(D3444_Y),     .C1(D3493_Y), .Y(D3468_Y));
KC_OAI211_X1 D3466 ( .B(D3485_Y), .C0(D4925_Y), .A(D4943_Y),     .C1(D3434_Y), .Y(D3466_Y));
KC_OAI211_X1 D3463 ( .B(D3422_Y), .C0(D3520_Y), .A(D3539_Y),     .C1(D3438_Y), .Y(D3463_Y));
KC_OAI211_X1 D3461 ( .B(D3538_Y), .C0(D3447_Y), .A(D3418_Y),     .C1(D3428_Y), .Y(D3461_Y));
KC_OAI211_X1 D3457 ( .B(D1450_Y), .C0(D3428_Y), .A(D3486_Y),     .C1(D3539_Y), .Y(D3457_Y));
KC_OAI211_X1 D3456 ( .B(D4889_Y), .C0(D4926_Y), .A(D3465_Y),     .C1(D3428_Y), .Y(D3456_Y));
KC_OAI211_X1 D3159 ( .B(D3137_Y), .C0(D1429_Y), .A(D3183_Y),     .C1(D3252_Y), .Y(D3159_Y));
KC_OAI211_X1 D3044 ( .B(D3027_Y), .C0(D3021_Y), .A(D39_Y),     .C1(D3027_Y), .Y(D3044_Y));
KC_OAI211_X1 D2950 ( .B(D2903_Y), .C0(D2904_Y), .A(D2997_Y),     .C1(D2952_Y), .Y(D2950_Y));
KC_OAI211_X1 D2779 ( .B(D2766_Y), .C0(D2741_Y), .A(D2769_Y),     .C1(D2762_Y), .Y(D2779_Y));
KC_OAI211_X1 D2776 ( .B(D2793_Y), .C0(D2744_Y), .A(D2748_Y),     .C1(D2838_Y), .Y(D2776_Y));
KC_OAI211_X1 D2772 ( .B(D2901_Y), .C0(D2895_Y), .A(D2783_Y),     .C1(D2901_Y), .Y(D2772_Y));
KC_OAI211_X1 D2626 ( .B(D2602_Y), .C0(D16767_Y), .A(D15775_Y),     .C1(D9617_Y), .Y(D2626_Y));
KC_OAI211_X1 D2625 ( .B(D2601_Y), .C0(D13610_Y), .A(D2623_Y),     .C1(D813_Y), .Y(D2625_Y));
KC_OAI211_X1 D2621 ( .B(D1093_Y), .C0(D2471_Y), .A(D2622_Y),     .C1(D813_Y), .Y(D2621_Y));
KC_OAI211_X1 D2620 ( .B(D2598_Y), .C0(D16767_Y), .A(D15749_Y),     .C1(D813_Y), .Y(D2620_Y));
KC_OAI211_X1 D2619 ( .B(D2597_Y), .C0(D86_Y), .A(D15854_Y),     .C1(D1813_Y), .Y(D2619_Y));
KC_OAI211_X1 D2562 ( .B(D14724_Y), .C0(D14148_Y), .A(D14101_Y),     .C1(D6410_Y), .Y(D2562_Y));
KC_OAI211_X1 D2561 ( .B(D2542_Y), .C0(D14148_Y), .A(D839_Y),     .C1(D10358_Y), .Y(D2561_Y));
KC_OAI211_X1 D2560 ( .B(D2541_Y), .C0(D14148_Y), .A(D838_Y),     .C1(D8336_Y), .Y(D2560_Y));
KC_OAI211_X1 D2557 ( .B(D2532_Y), .C0(D10358_Y), .A(D2558_Y),     .C1(D13619_Y), .Y(D2557_Y));
KC_OAI211_X1 D2556 ( .B(D14953_Y), .C0(D2471_Y), .A(D15776_Y),     .C1(D9617_Y), .Y(D2556_Y));
KC_OAI211_X1 D2554 ( .B(D2531_Y), .C0(D2487_Y), .A(D15063_Y),     .C1(D813_Y), .Y(D2554_Y));
KC_OAI211_X1 D2551 ( .B(D15073_Y), .C0(D2487_Y), .A(D15114_Y),     .C1(D6410_Y), .Y(D2551_Y));
KC_OAI211_X1 D2550 ( .B(D14347_Y), .C0(D10191_Y), .A(D2553_Y),     .C1(D13619_Y), .Y(D2550_Y));
KC_OAI211_X1 D2549 ( .B(D15173_Y), .C0(D13622_Y), .A(D15121_Y),     .C1(D10191_Y), .Y(D2549_Y));
KC_OAI211_X1 D2502 ( .B(D14134_Y), .C0(D13313_Y), .A(D14029_Y),     .C1(D13473_Y), .Y(D2502_Y));
KC_OAI211_X1 D2443 ( .B(D13466_Y), .C0(D2422_Y), .A(D2436_Y),     .C1(D13338_Y), .Y(D2443_Y));
KC_OAI211_X1 D2440 ( .B(D13631_Y), .C0(D13541_Y), .A(D13658_Y),     .C1(D2415_Y), .Y(D2440_Y));
KC_OAI211_X1 D2439 ( .B(D13776_Y), .C0(D13610_Y), .A(D13744_Y),     .C1(D10192_Y), .Y(D2439_Y));
KC_OAI211_X1 D2380 ( .B(D13435_Y), .C0(D929_Q), .A(D13538_Y),     .C1(D12929_Y), .Y(D2380_Y));
KC_OAI211_X1 D2379 ( .B(D2312_Y), .C0(D12661_Y), .A(D2343_Y),     .C1(D161_Y), .Y(D2379_Y));
KC_OAI211_X1 D2143 ( .B(D10253_Y), .C0(D1990_Y), .A(D9483_Y),     .C1(D10296_Q), .Y(D2143_Y));
KC_OAI211_X1 D2142 ( .B(D2124_Y), .C0(D7407_Y), .A(D10029_Y),     .C1(D8949_Y), .Y(D2142_Y));
KC_OAI211_X1 D2141 ( .B(D8930_Y), .C0(D7407_Y), .A(D10014_Y),     .C1(D10043_Y), .Y(D2141_Y));
KC_OAI211_X1 D2138 ( .B(D10508_Q), .C0(D10388_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D2138_Y));
KC_OAI211_X1 D2111 ( .B(D9787_Q), .C0(D9642_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D2111_Y));
KC_OAI211_X1 D2051 ( .B(D8941_Y), .C0(D8851_Y), .A(D8857_Y),     .C1(D9016_Y), .Y(D2051_Y));
KC_OAI211_X1 D2048 ( .B(D9001_Y), .C0(D8904_Y), .A(D74_Y),     .C1(D8980_Y), .Y(D2048_Y));
KC_OAI211_X1 D2047 ( .B(D9097_Y), .C0(D8948_Y), .A(D8964_Y),     .C1(D5703_Y), .Y(D2047_Y));
KC_OAI211_X1 D2046 ( .B(D9098_Y), .C0(D8973_Y), .A(D2013_Y),     .C1(D5703_Y), .Y(D2046_Y));
KC_OAI211_X1 D2039 ( .B(D9432_Y), .C0(D1897_Y), .A(D9388_Y),     .C1(D1989_Y), .Y(D2039_Y));
KC_OAI211_X1 D2037 ( .B(D9687_Y), .C0(D9640_Y), .A(D2035_Y),     .C1(D9746_Y), .Y(D2037_Y));
KC_OAI211_X1 D2036 ( .B(D9788_Q), .C0(D9640_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D2036_Y));
KC_OAI211_X1 D2035 ( .B(D9784_Q), .C0(D9641_Y), .A(D1919_Y),     .C1(D8542_Y), .Y(D2035_Y));
KC_OAI211_X1 D2034 ( .B(D9688_Y), .C0(D9642_Y), .A(D9766_Y),     .C1(D9746_Y), .Y(D2034_Y));
KC_OAI211_X1 D2031 ( .B(D9770_Y), .C0(D1978_Y), .A(D9768_Y),     .C1(D8550_Y), .Y(D2031_Y));
KC_OAI211_X1 D1908 ( .B(D1884_Y), .C0(D7271_Y), .A(D1909_Y),     .C1(D7201_Y), .Y(D1908_Y));
KC_OAI211_X1 D1898 ( .B(D8163_Y), .C0(D8146_Y), .A(D8157_Y),     .C1(D8006_Y), .Y(D1898_Y));
KC_OAI211_X1 D1891 ( .B(D8534_Y), .C0(D8377_Y), .A(D8361_Y),     .C1(D8360_Y), .Y(D1891_Y));
KC_OAI211_X1 D1890 ( .B(D1892_Y), .C0(D6864_Y), .A(D8428_Y),     .C1(D8550_Y), .Y(D1890_Y));
KC_OAI211_X1 D1889 ( .B(D1929_Q), .C0(D8423_Y), .A(D1919_Y),     .C1(D8363_Y), .Y(D1889_Y));
KC_OAI211_X1 D1820 ( .B(D1853_Y), .C0(D1821_Y), .A(D168_Y),     .C1(D471_Y), .Y(D1820_Y));
KC_OAI211_X1 D1816 ( .B(D7300_Y), .C0(D5874_Y), .A(D1734_Y),     .C1(D7419_Y), .Y(D1816_Y));
KC_OAI211_X1 D1754 ( .B(D5939_Y), .C0(D5747_Y), .A(D206_Y),     .C1(D5994_Y), .Y(D1754_Y));
KC_OAI211_X1 D1751 ( .B(D1720_Y), .C0(D5792_Y), .A(D5899_Y),     .C1(D6020_Y), .Y(D1751_Y));
KC_OAI211_X1 D1750 ( .B(D1715_Y), .C0(D6010_Y), .A(D6019_Y),     .C1(D5726_Y), .Y(D1750_Y));
KC_OAI211_X1 D1748 ( .B(D6065_Y), .C0(D7499_Y), .A(D239_Q),     .C1(D5969_Y), .Y(D1748_Y));
KC_OAI211_X1 D1613 ( .B(D4154_Y), .C0(D4292_Y), .A(D1588_Y),     .C1(D6034_Y), .Y(D1613_Y));
KC_OAI211_X1 D1609 ( .B(D4612_Y), .C0(D4524_Y), .A(D1431_Y),     .C1(D4595_Y), .Y(D1609_Y));
KC_OAI211_X1 D1608 ( .B(D1575_Y), .C0(D4504_Y), .A(D4502_Y),     .C1(D3169_Y), .Y(D1608_Y));
KC_OAI211_X1 D1601 ( .B(D1414_Y), .C0(D5032_Y), .A(D5034_Y),     .C1(D4914_Y), .Y(D1601_Y));
KC_OAI211_X1 D1600 ( .B(D433_Y), .C0(D4960_Y), .A(D4859_Y),     .C1(D1558_Y), .Y(D1600_Y));
KC_OAI211_X1 D1451 ( .B(D3371_Y), .C0(D3303_Y), .A(D1537_Y),     .C1(D1570_Y), .Y(D1451_Y));
KC_OAI211_X1 D1283 ( .B(D14411_Y), .C0(D13641_Y), .A(D13793_Y),     .C1(D10192_Y), .Y(D1283_Y));
KC_OAI211_X1 D1282 ( .B(D15222_Y), .C0(D2420_Y), .A(D15983_Y),     .C1(D6406_Y), .Y(D1282_Y));
KC_OAI211_X1 D1191 ( .B(D14346_Y), .C0(D1964_Y), .A(D15115_Y),     .C1(D13619_Y), .Y(D1191_Y));
KC_OAI211_X1 D1189 ( .B(D15903_Y), .C0(D16767_Y), .A(D15924_Y),     .C1(D6406_Y), .Y(D1189_Y));
KC_OAI211_X1 D1187 ( .B(D8567_Y), .C0(D9830_Y), .A(D8519_Y),     .C1(D8550_Y), .Y(D1187_Y));
KC_OAI211_X1 D1166 ( .B(D1212_Q), .C0(D9830_Y), .A(D8534_Y),     .C1(D8542_Y), .Y(D1166_Y));
KC_OAI211_X1 D1164 ( .B(D13707_Y), .C0(D13011_Y), .A(D13652_Y),     .C1(D13016_Y), .Y(D1164_Y));
KC_OAI211_X1 D1106 ( .B(D15864_Y), .C0(D86_Y), .A(D15845_Y),     .C1(D1814_Y), .Y(D1106_Y));
KC_OAI211_X1 D1103 ( .B(D9754_Y), .C0(D8420_Y), .A(D9765_Y),     .C1(D9746_Y), .Y(D1103_Y));
KC_OAI211_X1 D1101 ( .B(D1104_Y), .C0(D10454_Y), .A(D10484_Y),     .C1(D9746_Y), .Y(D1101_Y));
KC_OAI211_X1 D1100 ( .B(D990_Y), .C0(D10455_Y), .A(D9684_Y),     .C1(D9746_Y), .Y(D1100_Y));
KC_OAI211_X1 D1099 ( .B(D2038_Y), .C0(D9641_Y), .A(D8515_Y),     .C1(D8550_Y), .Y(D1099_Y));
KC_OAI211_X1 D1097 ( .B(D10473_Y), .C0(D9728_Y), .A(D10475_Y),     .C1(D9746_Y), .Y(D1097_Y));
KC_OAI211_X1 D1096 ( .B(D9755_Y), .C0(D8485_Y), .A(D9769_Y),     .C1(D8550_Y), .Y(D1096_Y));
KC_OAI211_X1 D1078 ( .B(D991_Y), .C0(D8423_Y), .A(D8427_Y),     .C1(D9746_Y), .Y(D1078_Y));
KC_OAI211_X1 D998 ( .B(D14950_Y), .C0(D13622_Y), .A(D14227_Y),     .C1(D9617_Y), .Y(D998_Y));
KC_OAI211_X1 D996 ( .B(D15738_Y), .C0(D13610_Y), .A(D15761_Y),     .C1(D10358_Y), .Y(D996_Y));
KC_OAI211_X1 D994 ( .B(D14918_Y), .C0(D813_Y), .A(D14223_Y),     .C1(D13619_Y), .Y(D994_Y));
KC_OAI211_X1 D876 ( .B(D13435_Y), .C0(D146_Q), .A(D13417_Y),     .C1(D12932_Y), .Y(D876_Y));
KC_OAI211_X1 D761 ( .B(D836_Q), .C0(D9524_Y), .A(D9540_Y),     .C1(D9516_Y), .Y(D761_Y));
KC_OAI211_X1 D642 ( .B(D9401_Y), .C0(D9421_Y), .A(D8085_Y),     .C1(D9402_Y), .Y(D642_Y));
KC_OAI211_X1 D574 ( .B(D15321_Y), .C0(D570_Y), .A(D568_Y),     .C1(D15295_Y), .Y(D574_Y));
KC_OAI211_X1 D491 ( .B(D3400_Y), .C0(D5004_Y), .A(D5091_Y),     .C1(D3525_Y), .Y(D491_Y));
KC_OAI211_X1 D474 ( .B(D5019_Y), .C0(D3574_Y), .A(D3521_Y),     .C1(D3420_Y), .Y(D474_Y));
KC_OAI211_X1 D473 ( .B(D5005_Y), .C0(D3520_Y), .A(D4992_Y),     .C1(D3502_Y), .Y(D473_Y));
KC_OAI211_X1 D472 ( .B(D7825_Y), .C0(D6427_Y), .A(D6424_Y),     .C1(D6425_Y), .Y(D472_Y));
KC_OAI211_X1 D439 ( .B(D4949_Y), .C0(D4951_Y), .A(D4901_Y),     .C1(D6376_Q), .Y(D439_Y));
KC_OAI211_X1 D410 ( .B(D4759_Y), .C0(D4768_Y), .A(D4746_Y),     .C1(D3325_Y), .Y(D410_Y));
KC_OAI211_X1 D409 ( .B(D4697_Y), .C0(D4762_Y), .A(D4751_Y),     .C1(D3325_Y), .Y(D409_Y));
KC_OAI211_X1 D408 ( .B(D3394_Y), .C0(D4922_Y), .A(D1671_Y),     .C1(D5005_Y), .Y(D408_Y));
KC_OAI211_X1 D313 ( .B(D8907_Y), .C0(D9016_Y), .A(D8966_Y),     .C1(D8980_Y), .Y(D313_Y));
KC_OAI211_X1 D311 ( .B(D8907_Y), .C0(D8972_Y), .A(D8968_Y),     .C1(D8980_Y), .Y(D311_Y));
KC_OAI211_X1 D292 ( .B(D8934_Y), .C0(D7407_Y), .A(D10016_Y),     .C1(D8948_Y), .Y(D292_Y));
KC_OAI211_X1 D258 ( .B(D10001_Y), .C0(D10000_Y), .A(D8906_Y),     .C1(D7407_Y), .Y(D258_Y));
KC_OAI211_X1 D256 ( .B(D9991_Y), .C0(D10028_Y), .A(D248_Y),     .C1(D242_Y), .Y(D256_Y));
KC_OAI211_X1 D254 ( .B(D288_Y), .C0(D7319_Y), .A(D7326_Y), .C1(D214_Y),     .Y(D254_Y));
KC_OAI211_X1 D221 ( .B(D5942_Y), .C0(D5721_Y), .A(D4200_Y),     .C1(D7294_Y), .Y(D221_Y));
KC_OAI211_X1 D198 ( .B(D5643_Y), .C0(D4257_Y), .A(D4146_Y),     .C1(D7376_Y), .Y(D198_Y));
KC_OAI211_X1 D184 ( .B(D4216_Y), .C0(D4263_Y), .A(D178_Y),     .C1(D7376_Y), .Y(D184_Y));
KC_OAI211_X1 D183 ( .B(D8669_Y), .C0(D205_Y), .A(D8746_Y),     .C1(D9941_Q), .Y(D183_Y));
KC_OAI211_X1 D97 ( .B(D2534_Y), .C0(D13619_Y), .A(D14226_Y),     .C1(D9617_Y), .Y(D97_Y));
KC_OAI211_X1 D96 ( .B(D14927_Y), .C0(D1111_Y), .A(D15813_Y),     .C1(D16765_Y), .Y(D96_Y));
KC_OAI211_X1 D95 ( .B(D15108_Y), .C0(D13622_Y), .A(D15979_Y),     .C1(D6406_Y), .Y(D95_Y));
KC_OAI211_X1 D93 ( .B(D6011_Y), .C0(D1721_Y), .A(D6010_Y),     .C1(D6068_Y), .Y(D93_Y));
KC_OAI211_X1 D90 ( .B(D2139_Y), .C0(D9648_Y), .A(D10481_Y),     .C1(D9746_Y), .Y(D90_Y));
KC_OAI31_X1 D16529 ( .B2(D1385_Q), .B1(D16771_Y), .B0(D16545_Y),     .Y(D16529_Y), .A(D16612_Y));
KC_OAI31_X1 D16496 ( .B2(D1344_Y), .B1(D16507_Y), .B0(D16517_Y),     .Y(D16496_Y), .A(D16382_Y));
KC_OAI31_X1 D16491 ( .B2(D14651_Y), .B1(D13988_Y), .B0(D16490_Y),     .Y(D16491_Y), .A(D16492_Y));
KC_OAI31_X1 D16407 ( .B2(D16428_Y), .B1(D16437_Y), .B0(D16427_Y),     .Y(D16407_Y), .A(D16382_Y));
KC_OAI31_X1 D16260 ( .B2(D2662_Y), .B1(D16253_Y), .B0(D2661_Y),     .Y(D16260_Y), .A(D16382_Y));
KC_OAI31_X1 D16246 ( .B2(D16264_Y), .B1(D16253_Y), .B0(D16270_Y),     .Y(D16246_Y), .A(D16255_Y));
KC_OAI31_X1 D15813 ( .B2(D2678_Q), .B1(D16364_Q), .B0(D2633_Y),     .Y(D15813_Y), .A(D16765_Y));
KC_OAI31_X1 D15635 ( .B2(D15480_Y), .B1(D15466_Y), .B0(D15633_Y),     .Y(D15635_Y), .A(D15636_Y));
KC_OAI31_X1 D15360 ( .B2(D15359_Y), .B1(D15361_Y), .B0(D15513_Y),     .Y(D15360_Y), .A(D15461_Y));
KC_OAI31_X1 D15180 ( .B2(D1270_Y), .B1(D15164_Y), .B0(D14085_Y),     .Y(D15180_Y), .A(D15194_Y));
KC_OAI31_X1 D15095 ( .B2(D15881_Y), .B1(D15099_Y), .B0(D13982_Y),     .Y(D15095_Y), .A(D15112_Y));
KC_OAI31_X1 D15038 ( .B2(D15822_Y), .B1(D15032_Y), .B0(D13983_Y),     .Y(D15038_Y), .A(D15065_Y));
KC_OAI31_X1 D14960 ( .B2(D14959_Y), .B1(D2537_Y), .B0(D14086_Y),     .Y(D14960_Y), .A(D14977_Y));
KC_OAI31_X1 D14927 ( .B2(D16318_Q), .B1(D16315_Q), .B0(D14969_Y),     .Y(D14927_Y), .A(D14081_Y));
KC_OAI31_X1 D14851 ( .B2(D818_Q), .B1(D853_Q), .B0(D14718_Y),     .Y(D14851_Y), .A(D14864_Y));
KC_OAI31_X1 D14844 ( .B2(D14787_Q), .B1(D14789_Q), .B0(D14877_Q),     .Y(D14844_Y), .A(D13982_Y));
KC_OAI31_X1 D14837 ( .B2(D14817_Y), .B1(D2538_Y), .B0(D14002_Y),     .Y(D14837_Y), .A(D14857_Y));
KC_OAI31_X1 D14754 ( .B2(D14676_Y), .B1(D14664_Y), .B0(D13968_Y),     .Y(D14754_Y), .A(D14748_Y));
KC_OAI31_X1 D14546 ( .B2(D2574_Q), .B1(D14547_Y), .B0(D14572_Y),     .Y(D14546_Y), .A(D14550_Y));
KC_OAI31_X1 D14478 ( .B2(D14479_Y), .B1(D13804_Q), .B0(D14481_Y),     .Y(D14478_Y), .A(D14482_Y));
KC_OAI31_X1 D14452 ( .B2(D14451_Y), .B1(D13811_Q), .B0(D13774_Y),     .Y(D14452_Y), .A(D14448_Y));
KC_OAI31_X1 D14445 ( .B2(D14443_Y), .B1(D13809_Q), .B0(D13779_Y),     .Y(D14445_Y), .A(D14442_Y));
KC_OAI31_X1 D14400 ( .B2(D14399_Y), .B1(D13807_Q), .B0(D14455_Y),     .Y(D14400_Y), .A(D14401_Y));
KC_OAI31_X1 D14359 ( .B2(D14358_Y), .B1(D13760_Q), .B0(D13717_Y),     .Y(D14359_Y), .A(D14433_Y));
KC_OAI31_X1 D14355 ( .B2(D14435_Y), .B1(D14356_Y), .B0(D14090_Y),     .Y(D14355_Y), .A(D14369_Y));
KC_OAI31_X1 D14354 ( .B2(D14352_Y), .B1(D13764_Q), .B0(D13729_Y),     .Y(D14354_Y), .A(D14345_Y));
KC_OAI31_X1 D14342 ( .B2(D15171_Y), .B1(D14348_Y), .B0(D14089_Y),     .Y(D14342_Y), .A(D14366_Y));
KC_OAI31_X1 D14341 ( .B2(D14444_Y), .B1(D14343_Y), .B0(D14082_Y),     .Y(D14341_Y), .A(D14361_Y));
KC_OAI31_X1 D14205 ( .B2(D14264_Q), .B1(D14242_Q), .B0(D14233_Y),     .Y(D14205_Y), .A(D13391_Y));
KC_OAI31_X1 D14136 ( .B2(D14093_Q), .B1(D14092_Q), .B0(D14030_Y),     .Y(D14136_Y), .A(D14149_Y));
KC_OAI31_X1 D14122 ( .B2(D14120_Y), .B1(D14127_Y), .B0(D777_Y),     .Y(D14122_Y), .A(D14143_Y));
KC_OAI31_X1 D13934 ( .B2(D13932_Y), .B1(D13963_Y), .B0(D14618_Y),     .Y(D13934_Y), .A(D13234_Y));
KC_OAI31_X1 D13890 ( .B2(D13918_Q), .B1(D13860_Q), .B0(D606_Y),     .Y(D13890_Y), .A(D13196_Q));
KC_OAI31_X1 D13726 ( .B2(D14334_Y), .B1(D13762_Q), .B0(D13716_Y),     .Y(D13726_Y), .A(D14332_Y));
KC_OAI31_X1 D13669 ( .B2(D13644_Y), .B1(D2414_Y), .B0(D778_Y),     .Y(D13669_Y), .A(D13692_Y));
KC_OAI31_X1 D13444 ( .B2(D13439_Y), .B1(D13447_Y), .B0(D13409_Y),     .Y(D13444_Y), .A(D13428_Y));
KC_OAI31_X1 D13406 ( .B2(D12241_Y), .B1(D2343_Y), .B0(D13309_Y),     .Y(D13406_Y), .A(D13329_Y));
KC_OAI31_X1 D13364 ( .B2(D13255_Y), .B1(D13342_Y), .B0(D13362_Y),     .Y(D13364_Y), .A(D13234_Y));
KC_OAI31_X1 D13307 ( .B2(D12241_Y), .B1(D2343_Y), .B0(D13473_Y),     .Y(D13307_Y), .A(D13329_Y));
KC_OAI31_X1 D13300 ( .B2(D12241_Y), .B1(D2343_Y), .B0(D13321_Y),     .Y(D13300_Y), .A(D13329_Y));
KC_OAI31_X1 D12892 ( .B2(D12897_Y), .B1(D12896_Y), .B0(D12871_Y),     .Y(D12892_Y), .A(D12904_Y));
KC_OAI31_X1 D12886 ( .B2(D12926_Q), .B1(D855_Q), .B0(D12880_Y),     .Y(D12886_Y), .A(D12801_Y));
KC_OAI31_X1 D12790 ( .B2(D12826_Y), .B1(D12789_Y), .B0(D12350_Q),     .Y(D12790_Y), .A(D12845_Y));
KC_OAI31_X1 D12722 ( .B2(D2353_Y), .B1(D12759_Q), .B0(D12658_Y),     .Y(D12722_Y), .A(D840_Y));
KC_OAI31_X1 D12208 ( .B2(D11657_Y), .B1(D6281_Y), .B0(D4747_Y),     .Y(D12208_Y), .A(D12194_Y));
KC_OAI31_X1 D12134 ( .B2(D495_Y), .B1(D496_Y), .B0(D12625_Y),     .Y(D12134_Y), .A(D3284_Y));
KC_OAI31_X1 D12029 ( .B2(D12059_Y), .B1(D1246_Q), .B0(D8551_Y),     .Y(D12029_Y), .A(D1173_Y));
KC_OAI31_X1 D12005 ( .B2(D12006_Y), .B1(D12042_Q), .B0(D8551_Y),     .Y(D12005_Y), .A(D1171_Y));
KC_OAI31_X1 D11999 ( .B2(D12000_Y), .B1(D12043_Q), .B0(D8551_Y),     .Y(D11999_Y), .A(D1175_Y));
KC_OAI31_X1 D11903 ( .B2(D11322_Y), .B1(D11358_Y), .B0(D11476_Y),     .Y(D11903_Y), .A(D11386_Y));
KC_OAI31_X1 D11893 ( .B2(D11322_Y), .B1(D11365_Y), .B0(D11476_Y),     .Y(D11893_Y), .A(D11386_Y));
KC_OAI31_X1 D11710 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11153_Y),     .Y(D11710_Y), .A(D11258_Y));
KC_OAI31_X1 D11700 ( .B2(D11322_Y), .B1(D11153_Y), .B0(D11476_Y),     .Y(D11700_Y), .A(D11258_Y));
KC_OAI31_X1 D11592 ( .B2(D2243_Y), .B1(D11549_Y), .B0(D11476_Y),     .Y(D11592_Y), .A(D11535_Y));
KC_OAI31_X1 D11562 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11547_Y),     .Y(D11562_Y), .A(D11536_Y));
KC_OAI31_X1 D11561 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11549_Y),     .Y(D11561_Y), .A(D11535_Y));
KC_OAI31_X1 D11560 ( .B2(D2243_Y), .B1(D11564_Y), .B0(D11476_Y),     .Y(D11560_Y), .A(D11535_Y));
KC_OAI31_X1 D11559 ( .B2(D2243_Y), .B1(D11547_Y), .B0(D11505_Y),     .Y(D11559_Y), .A(D11536_Y));
KC_OAI31_X1 D11558 ( .B2(D2243_Y), .B1(D11563_Y), .B0(D11476_Y),     .Y(D11558_Y), .A(D11535_Y));
KC_OAI31_X1 D11557 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11564_Y),     .Y(D11557_Y), .A(D11535_Y));
KC_OAI31_X1 D11556 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11563_Y),     .Y(D11556_Y), .A(D11535_Y));
KC_OAI31_X1 D11555 ( .B2(D2243_Y), .B1(D11554_Y), .B0(D11476_Y),     .Y(D11555_Y), .A(D11535_Y));
KC_OAI31_X1 D11545 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11554_Y),     .Y(D11545_Y), .A(D11535_Y));
KC_OAI31_X1 D11544 ( .B2(D2243_Y), .B1(D11552_Y), .B0(D11505_Y),     .Y(D11544_Y), .A(D11536_Y));
KC_OAI31_X1 D11512 ( .B2(D11494_Y), .B1(D1224_Q), .B0(D8551_Y),     .Y(D11512_Y), .A(D11480_Y));
KC_OAI31_X1 D11511 ( .B2(D11479_Y), .B1(D1219_Q), .B0(D8551_Y),     .Y(D11511_Y), .A(D11495_Y));
KC_OAI31_X1 D11510 ( .B2(D11491_Y), .B1(D131_Q), .B0(D8551_Y),     .Y(D11510_Y), .A(D11482_Y));
KC_OAI31_X1 D11509 ( .B2(D11499_Y), .B1(D11537_Q), .B0(D8551_Y),     .Y(D11509_Y), .A(D11497_Y));
KC_OAI31_X1 D11508 ( .B2(D11484_Y), .B1(D11538_Q), .B0(D8551_Y),     .Y(D11508_Y), .A(D11489_Y));
KC_OAI31_X1 D11507 ( .B2(D11488_Y), .B1(D11542_Q), .B0(D8551_Y),     .Y(D11507_Y), .A(D11485_Y));
KC_OAI31_X1 D11506 ( .B2(D11493_Y), .B1(D11539_Q), .B0(D8551_Y),     .Y(D11506_Y), .A(D11496_Y));
KC_OAI31_X1 D11503 ( .B2(D11504_Y), .B1(D2249_Q), .B0(D8551_Y),     .Y(D11503_Y), .A(D11501_Y));
KC_OAI31_X1 D11502 ( .B2(D11490_Y), .B1(D2251_Q), .B0(D8551_Y),     .Y(D11502_Y), .A(D11500_Y));
KC_OAI31_X1 D11487 ( .B2(D11483_Y), .B1(D11543_Q), .B0(D8551_Y),     .Y(D11487_Y), .A(D11498_Y));
KC_OAI31_X1 D11486 ( .B2(D11481_Y), .B1(D1218_Q), .B0(D8551_Y),     .Y(D11486_Y), .A(D11015_Y));
KC_OAI31_X1 D11437 ( .B2(D11419_Y), .B1(D11466_Q), .B0(D11259_Y),     .Y(D11437_Y), .A(D11423_Y));
KC_OAI31_X1 D11436 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11379_Y),     .Y(D11436_Y), .A(D11386_Y));
KC_OAI31_X1 D11435 ( .B2(D11431_Y), .B1(D11468_Q), .B0(D11259_Y),     .Y(D11435_Y), .A(D11433_Y));
KC_OAI31_X1 D11430 ( .B2(D11432_Y), .B1(D2253_Q), .B0(D11259_Y),     .Y(D11430_Y), .A(D11434_Y));
KC_OAI31_X1 D11424 ( .B2(D11426_Y), .B1(D11469_Q), .B0(D11259_Y),     .Y(D11424_Y), .A(D11422_Y));
KC_OAI31_X1 D11420 ( .B2(D11425_Y), .B1(D11475_Q), .B0(D11259_Y),     .Y(D11420_Y), .A(D11429_Y));
KC_OAI31_X1 D11375 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11365_Y),     .Y(D11375_Y), .A(D11386_Y));
KC_OAI31_X1 D11374 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11358_Y),     .Y(D11374_Y), .A(D11386_Y));
KC_OAI31_X1 D11373 ( .B2(D11372_Y), .B1(D11389_Q), .B0(D10770_Y),     .Y(D11373_Y), .A(D2231_Y));
KC_OAI31_X1 D11369 ( .B2(D11322_Y), .B1(D11377_Y), .B0(D11476_Y),     .Y(D11369_Y), .A(D11386_Y));
KC_OAI31_X1 D11364 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11377_Y),     .Y(D11364_Y), .A(D11386_Y));
KC_OAI31_X1 D11357 ( .B2(D11366_Y), .B1(D11340_Q), .B0(D11259_Y),     .Y(D11357_Y), .A(D11356_Y));
KC_OAI31_X1 D11353 ( .B2(D11322_Y), .B1(D11379_Y), .B0(D11476_Y),     .Y(D11353_Y), .A(D11386_Y));
KC_OAI31_X1 D11352 ( .B2(D11354_Y), .B1(D11392_Q), .B0(D11259_Y),     .Y(D11352_Y), .A(D11351_Y));
KC_OAI31_X1 D11303 ( .B2(D11308_Y), .B1(D11305_Y), .B0(D11476_Y),     .Y(D11303_Y), .A(D11256_Y));
KC_OAI31_X1 D11300 ( .B2(D11297_Y), .B1(D11325_Q), .B0(D11259_Y),     .Y(D11300_Y), .A(D11290_Y));
KC_OAI31_X1 D11299 ( .B2(D11302_Y), .B1(D11327_Q), .B0(D11259_Y),     .Y(D11299_Y), .A(D11301_Y));
KC_OAI31_X1 D11294 ( .B2(D11295_Y), .B1(D11342_Q), .B0(D11259_Y),     .Y(D11294_Y), .A(D11298_Y));
KC_OAI31_X1 D11293 ( .B2(D10861_Y), .B1(D11308_Y), .B0(D11305_Y),     .Y(D11293_Y), .A(D11256_Y));
KC_OAI31_X1 D11292 ( .B2(D11296_Y), .B1(D11329_Q), .B0(D11259_Y),     .Y(D11292_Y), .A(D11289_Y));
KC_OAI31_X1 D11286 ( .B2(D11287_Y), .B1(D11326_Q), .B0(D11259_Y),     .Y(D11286_Y), .A(D11284_Y));
KC_OAI31_X1 D11285 ( .B2(D11288_Y), .B1(D11341_Q), .B0(D11259_Y),     .Y(D11285_Y), .A(D11291_Y));
KC_OAI31_X1 D11230 ( .B2(D11209_Y), .B1(D11262_Q), .B0(D11259_Y),     .Y(D11230_Y), .A(D11206_Y));
KC_OAI31_X1 D11229 ( .B2(D11204_Y), .B1(D11263_Q), .B0(D10770_Y),     .Y(D11229_Y), .A(D11198_Y));
KC_OAI31_X1 D11202 ( .B2(D746_Y), .B1(D11261_Q), .B0(D11259_Y),     .Y(D11202_Y), .A(D11207_Y));
KC_OAI31_X1 D11201 ( .B2(D11210_Y), .B1(D11265_Q), .B0(D11259_Y),     .Y(D11201_Y), .A(D11208_Y));
KC_OAI31_X1 D11199 ( .B2(D11205_Y), .B1(D11264_Q), .B0(D10770_Y),     .Y(D11199_Y), .A(D11203_Y));
KC_OAI31_X1 D11197 ( .B2(D744_Y), .B1(D2256_Q), .B0(D11259_Y),     .Y(D11197_Y), .A(D11195_Y));
KC_OAI31_X1 D11196 ( .B2(D11738_Y), .B1(D136_Q), .B0(D11259_Y),     .Y(D11196_Y), .A(D11736_Y));
KC_OAI31_X1 D11193 ( .B2(D11200_Y), .B1(D797_Q), .B0(D10770_Y),     .Y(D11193_Y), .A(D745_Y));
KC_OAI31_X1 D11190 ( .B2(D11259_Y), .B1(D11260_Q), .B0(D11737_Y),     .Y(D11190_Y), .A(D742_Y));
KC_OAI31_X1 D11188 ( .B2(D11194_Y), .B1(D135_Q), .B0(D10770_Y),     .Y(D11188_Y), .A(D2232_Y));
KC_OAI31_X1 D11151 ( .B2(D11322_Y), .B1(D11143_Y), .B0(D11476_Y),     .Y(D11151_Y), .A(D11258_Y));
KC_OAI31_X1 D11150 ( .B2(D11322_Y), .B1(D11144_Y), .B0(D11476_Y),     .Y(D11150_Y), .A(D11258_Y));
KC_OAI31_X1 D11149 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11154_Y),     .Y(D11149_Y), .A(D11258_Y));
KC_OAI31_X1 D11147 ( .B2(D11322_Y), .B1(D11154_Y), .B0(D11476_Y),     .Y(D11147_Y), .A(D11258_Y));
KC_OAI31_X1 D11142 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11144_Y),     .Y(D11142_Y), .A(D11258_Y));
KC_OAI31_X1 D11062 ( .B2(D2243_Y), .B1(D11566_Y), .B0(D11505_Y),     .Y(D11062_Y), .A(D11536_Y));
KC_OAI31_X1 D10981 ( .B2(D10980_Y), .B1(D2250_Q), .B0(D8551_Y),     .Y(D10981_Y), .A(D10979_Y));
KC_OAI31_X1 D10857 ( .B2(D10861_Y), .B1(D11308_Y), .B0(D10862_Y),     .Y(D10857_Y), .A(D11256_Y));
KC_OAI31_X1 D10853 ( .B2(D10861_Y), .B1(D11308_Y), .B0(D10847_Y),     .Y(D10853_Y), .A(D11256_Y));
KC_OAI31_X1 D10851 ( .B2(D11308_Y), .B1(D10855_Y), .B0(D11476_Y),     .Y(D10851_Y), .A(D11256_Y));
KC_OAI31_X1 D10850 ( .B2(D11308_Y), .B1(D10862_Y), .B0(D11476_Y),     .Y(D10850_Y), .A(D11256_Y));
KC_OAI31_X1 D10848 ( .B2(D11308_Y), .B1(D10847_Y), .B0(D11476_Y),     .Y(D10848_Y), .A(D11256_Y));
KC_OAI31_X1 D10844 ( .B2(D10861_Y), .B1(D11308_Y), .B0(D10855_Y),     .Y(D10844_Y), .A(D11256_Y));
KC_OAI31_X1 D10740 ( .B2(D10744_Y), .B1(D10792_Q), .B0(D10770_Y),     .Y(D10740_Y), .A(D10738_Y));
KC_OAI31_X1 D10739 ( .B2(D2205_Y), .B1(D10789_Q), .B0(D10770_Y),     .Y(D10739_Y), .A(D10733_Y));
KC_OAI31_X1 D10731 ( .B2(D2204_Y), .B1(D10793_Q), .B0(D10770_Y),     .Y(D10731_Y), .A(D10736_Y));
KC_OAI31_X1 D10180 ( .B2(D10177_Y), .B1(D11657_Y), .B0(D11655_Y),     .Y(D10180_Y), .A(D11660_Y));
KC_OAI31_X1 D10053 ( .B2(D11114_Y), .B1(D2122_Y), .B0(D2123_Y),     .Y(D10053_Y), .A(D9080_Y));
KC_OAI31_X1 D9537 ( .B2(D9577_Q), .B1(D9597_Y), .B0(D9543_Y),     .Y(D9537_Y), .A(D9587_Y));
KC_OAI31_X1 D9520 ( .B2(D9536_Y), .B1(D9597_Y), .B0(D9547_Y),     .Y(D9520_Y), .A(D9545_Y));
KC_OAI31_X1 D9500 ( .B2(D9579_Q), .B1(D9499_Y), .B0(D9501_Y),     .Y(D9500_Y), .A(D9588_Y));
KC_OAI31_X1 D9495 ( .B2(D2061_Y), .B1(D9672_Y), .B0(D9672_Y),     .Y(D9495_Y), .A(D2108_Y));
KC_OAI31_X1 D9426 ( .B2(D9473_Y), .B1(D9396_Y), .B0(D9407_Y),     .Y(D9426_Y), .A(D649_Y));
KC_OAI31_X1 D9404 ( .B2(D9413_Y), .B1(D9550_Y), .B0(D7655_Y),     .Y(D9404_Y), .A(D9399_Y));
KC_OAI31_X1 D9403 ( .B2(D9395_Y), .B1(D9431_Y), .B0(D9470_Q),     .Y(D9403_Y), .A(D9485_Y));
KC_OAI31_X1 D9397 ( .B2(D1987_Y), .B1(D8083_Y), .B0(D9442_Y),     .Y(D9397_Y), .A(D9444_Y));
KC_OAI31_X1 D9373 ( .B2(D9383_Y), .B1(D9383_Y), .B0(D9383_Y),     .Y(D9373_Y), .A(D9376_Y));
KC_OAI31_X1 D9126 ( .B2(D12305_Y), .B1(D7624_Y), .B0(D382_Y),     .Y(D9126_Y), .A(D9110_Y));
KC_OAI31_X1 D9077 ( .B2(D8061_Y), .B1(D8970_Y), .B0(D8971_Y),     .Y(D9077_Y), .A(D9048_Y));
KC_OAI31_X1 D9076 ( .B2(D8067_Y), .B1(D8970_Y), .B0(D9122_Y),     .Y(D9076_Y), .A(D9051_Y));
KC_OAI31_X1 D9075 ( .B2(D8065_Y), .B1(D8970_Y), .B0(D338_Y),     .Y(D9075_Y), .A(D9046_Y));
KC_OAI31_X1 D9074 ( .B2(D8066_Y), .B1(D8970_Y), .B0(D9109_Y),     .Y(D9074_Y), .A(D9035_Y));
KC_OAI31_X1 D9069 ( .B2(D8071_Y), .B1(D8970_Y), .B0(D9057_Y),     .Y(D9069_Y), .A(D9060_Y));
KC_OAI31_X1 D9061 ( .B2(D8070_Y), .B1(D8970_Y), .B0(D8985_Y),     .Y(D9061_Y), .A(D9049_Y));
KC_OAI31_X1 D9055 ( .B2(D615_Y), .B1(D8970_Y), .B0(D9056_Y),     .Y(D9055_Y), .A(D9096_Y));
KC_OAI31_X1 D8987 ( .B2(D9024_Y), .B1(D7490_Y), .B0(D2014_Y),     .Y(D8987_Y), .A(D58_Y));
KC_OAI31_X1 D8755 ( .B2(D8816_Y), .B1(D8774_Y), .B0(D8805_Y),     .Y(D8755_Y), .A(D8794_Y));
KC_OAI31_X1 D8674 ( .B2(D2030_Y), .B1(D8685_Y), .B0(D1977_Y),     .Y(D8674_Y), .A(D2058_Y));
KC_OAI31_X1 D8565 ( .B2(D8561_Y), .B1(D1927_Q), .B0(D8551_Y),     .Y(D8565_Y), .A(D8562_Y));
KC_OAI31_X1 D8557 ( .B2(D8558_Y), .B1(D8594_Q), .B0(D8551_Y),     .Y(D8557_Y), .A(D8560_Y));
KC_OAI31_X1 D8505 ( .B2(D8551_Y), .B1(D8538_Q), .B0(D1831_Y),     .Y(D8505_Y), .A(D1830_Y));
KC_OAI31_X1 D8426 ( .B2(D8362_Y), .B1(D11390_Q), .B0(D10770_Y),     .Y(D8426_Y), .A(D8469_Y));
KC_OAI31_X1 D8425 ( .B2(D1928_Q), .B1(D8500_Y), .B0(D6864_Y),     .Y(D8425_Y), .A(D8429_Y));
KC_OAI31_X1 D8411 ( .B2(D6873_Y), .B1(D1779_Q), .B0(D10770_Y),     .Y(D8411_Y), .A(D6870_Y));
KC_OAI31_X1 D8402 ( .B2(D8404_Y), .B1(D1930_Q), .B0(D10770_Y),     .Y(D8402_Y), .A(D975_Y));
KC_OAI31_X1 D8287 ( .B2(D6768_Y), .B1(D8463_Q), .B0(D10770_Y),     .Y(D8287_Y), .A(D8284_Y));
KC_OAI31_X1 D8203 ( .B2(D8082_Y), .B1(D796_Q), .B0(D8060_Y),     .Y(D8203_Y), .A(D8197_Y));
KC_OAI31_X1 D8179 ( .B2(D8060_Y), .B1(D784_Q), .B0(D6710_Y),     .Y(D8179_Y), .A(D734_Y));
KC_OAI31_X1 D8178 ( .B2(D8060_Y), .B1(D8238_Q), .B0(D8187_Y),     .Y(D8178_Y), .A(D8180_Y));
KC_OAI31_X1 D8169 ( .B2(D10770_Y), .B1(D785_Q), .B0(D8170_Y),     .Y(D8169_Y), .A(D8168_Y));
KC_OAI31_X1 D8122 ( .B2(D8060_Y), .B1(D676_Q), .B0(D8009_Y),     .Y(D8122_Y), .A(D1842_Y));
KC_OAI31_X1 D8114 ( .B2(D8060_Y), .B1(D672_Q), .B0(D8110_Y),     .Y(D8114_Y), .A(D8119_Y));
KC_OAI31_X1 D8101 ( .B2(D8077_Y), .B1(D9413_Y), .B0(D9407_Y),     .Y(D8101_Y), .A(D8100_Y));
KC_OAI31_X1 D8090 ( .B2(D8088_Y), .B1(D8083_Y), .B0(D8124_Y),     .Y(D8090_Y), .A(D9444_Y));
KC_OAI31_X1 D8022 ( .B2(D8000_Y), .B1(D8054_Q), .B0(D8060_Y),     .Y(D8022_Y), .A(D7995_Y));
KC_OAI31_X1 D8021 ( .B2(D7999_Y), .B1(D8053_Q), .B0(D8060_Y),     .Y(D8021_Y), .A(D8010_Y));
KC_OAI31_X1 D8014 ( .B2(D7994_Y), .B1(D8052_Q), .B0(D8060_Y),     .Y(D8014_Y), .A(D8012_Y));
KC_OAI31_X1 D7998 ( .B2(D8006_Y), .B1(D8055_Q), .B0(D8060_Y),     .Y(D7998_Y), .A(D7996_Y));
KC_OAI31_X1 D7997 ( .B2(D8008_Y), .B1(D669_Q), .B0(D8060_Y),     .Y(D7997_Y), .A(D8004_Y));
KC_OAI31_X1 D7440 ( .B2(D7433_Y), .B1(D7437_Y), .B0(D7350_Y),     .Y(D7440_Y), .A(D1878_Y));
KC_OAI31_X1 D7351 ( .B2(D7349_Y), .B1(D7397_Y), .B0(D7379_Y),     .Y(D7351_Y), .A(D5804_Y));
KC_OAI31_X1 D7350 ( .B2(D7634_Y), .B1(D7199_Y), .B0(D7214_Y),     .Y(D7350_Y), .A(D7372_Y));
KC_OAI31_X1 D7262 ( .B2(D5940_Y), .B1(D7287_Y), .B0(D7190_Y),     .Y(D7262_Y), .A(D5804_Y));
KC_OAI31_X1 D7261 ( .B2(D8801_Y), .B1(D7297_Y), .B0(D7275_Y),     .Y(D7261_Y), .A(D7249_Y));
KC_OAI31_X1 D7244 ( .B2(D7181_Y), .B1(D7187_Y), .B0(D7297_Y),     .Y(D7244_Y), .A(D7249_Y));
KC_OAI31_X1 D7235 ( .B2(D7276_Y), .B1(D7169_Y), .B0(D7174_Y),     .Y(D7235_Y), .A(D7249_Y));
KC_OAI31_X1 D7196 ( .B2(D7276_Y), .B1(D7226_Y), .B0(D7284_Y),     .Y(D7196_Y), .A(D7234_Y));
KC_OAI31_X1 D7168 ( .B2(D9480_Y), .B1(D9481_Y), .B0(D7178_Y),     .Y(D7168_Y), .A(D9475_Y));
KC_OAI31_X1 D7103 ( .B2(D6333_Y), .B1(D7120_Y), .B0(D7104_Y),     .Y(D7103_Y), .A(D7119_Y));
KC_OAI31_X1 D7094 ( .B2(D7137_Y), .B1(D189_Y), .B0(D7123_Y),     .Y(D7094_Y), .A(D7296_Y));
KC_OAI31_X1 D6995 ( .B2(D8500_Y), .B1(D1774_Q), .B0(D6989_Y),     .Y(D6995_Y), .A(D6990_Y));
KC_OAI31_X1 D6994 ( .B2(D6992_Y), .B1(D7005_Q), .B0(D8500_Y),     .Y(D6994_Y), .A(D6987_Y));
KC_OAI31_X1 D6993 ( .B2(D6986_Y), .B1(D7008_Q), .B0(D8500_Y),     .Y(D6993_Y), .A(D7017_Y));
KC_OAI31_X1 D6940 ( .B2(D8500_Y), .B1(D6970_Q), .B0(D6916_Y),     .Y(D6940_Y), .A(D6914_Y));
KC_OAI31_X1 D6939 ( .B2(D8500_Y), .B1(D1126_Q), .B0(D6931_Y),     .Y(D6939_Y), .A(D6933_Y));
KC_OAI31_X1 D6790 ( .B2(D5387_Y), .B1(D6780_Y), .B0(D3881_Y),     .Y(D6790_Y), .A(D5391_Y));
KC_OAI31_X1 D6779 ( .B2(D6777_Y), .B1(D3881_Y), .B0(D6780_Y),     .Y(D6779_Y), .A(D5391_Y));
KC_OAI31_X1 D6778 ( .B2(D3881_Y), .B1(D6784_Y), .B0(D6777_Y),     .Y(D6778_Y), .A(D5391_Y));
KC_OAI31_X1 D6776 ( .B2(D5387_Y), .B1(D3881_Y), .B0(D6784_Y),     .Y(D6776_Y), .A(D5391_Y));
KC_OAI31_X1 D6775 ( .B2(D6794_Y), .B1(D5387_Y), .B0(D6780_Y),     .Y(D6775_Y), .A(D5391_Y));
KC_OAI31_X1 D6774 ( .B2(D6794_Y), .B1(D5387_Y), .B0(D6784_Y),     .Y(D6774_Y), .A(D5391_Y));
KC_OAI31_X1 D6771 ( .B2(D6765_Y), .B1(D6829_Q), .B0(D10770_Y),     .Y(D6771_Y), .A(D8276_Y));
KC_OAI31_X1 D6764 ( .B2(D6767_Y), .B1(D6825_Q), .B0(D10770_Y),     .Y(D6764_Y), .A(D66_Y));
KC_OAI31_X1 D6718 ( .B2(D6720_Y), .B1(D6750_Q), .B0(D8060_Y),     .Y(D6718_Y), .A(D6706_Y));
KC_OAI31_X1 D6713 ( .B2(D8193_Y), .B1(D6754_Q), .B0(D8060_Y),     .Y(D6713_Y), .A(D736_Y));
KC_OAI31_X1 D6429 ( .B2(D6479_Y), .B1(D5017_Y), .B0(D6454_Y),     .Y(D6429_Y), .A(D7935_Y));
KC_OAI31_X1 D6428 ( .B2(D5038_Y), .B1(D4996_Y), .B0(D6430_Y),     .Y(D6428_Y), .A(D7935_Y));
KC_OAI31_X1 D6415 ( .B2(D6418_Y), .B1(D4959_Y), .B0(D6477_Y),     .Y(D6415_Y), .A(D6422_Y));
KC_OAI31_X1 D6151 ( .B2(D6182_Y), .B1(D6117_Y), .B0(D6253_Y),     .Y(D6151_Y), .A(D6202_Y));
KC_OAI31_X1 D6148 ( .B2(D6205_Y), .B1(D6149_Y), .B0(D6149_Y),     .Y(D6148_Y), .A(D56_Y));
KC_OAI31_X1 D6134 ( .B2(D7657_Y), .B1(D378_Y), .B0(D6137_Y),     .Y(D6134_Y), .A(D6153_Y));
KC_OAI31_X1 D6099 ( .B2(D13171_Y), .B1(D9268_Y), .B0(D7750_Y),     .Y(D6099_Y), .A(D6098_Y));
KC_OAI31_X1 D5894 ( .B2(D5868_Y), .B1(D6024_Y), .B0(D5888_Y),     .Y(D5894_Y), .A(D7337_Y));
KC_OAI31_X1 D5893 ( .B2(D7470_Y), .B1(D5918_Y), .B0(D5928_Y),     .Y(D5893_Y), .A(D5850_Y));
KC_OAI31_X1 D5883 ( .B2(D5867_Y), .B1(D5651_Y), .B0(D4316_Y),     .Y(D5883_Y), .A(D1731_Y));
KC_OAI31_X1 D5873 ( .B2(D4343_Y), .B1(D5867_Y), .B0(D5876_Y),     .Y(D5873_Y), .A(D1969_Y));
KC_OAI31_X1 D5709 ( .B2(D1614_Y), .B1(D5719_Y), .B0(D5791_Y),     .Y(D5709_Y), .A(D5804_Y));
KC_OAI31_X1 D5708 ( .B2(D5717_Y), .B1(D7281_Y), .B0(D5720_Y),     .Y(D5708_Y), .A(D5804_Y));
KC_OAI31_X1 D5650 ( .B2(D5688_Q), .B1(D5880_Y), .B0(D5655_Y),     .Y(D5650_Y), .A(D5804_Y));
KC_OAI31_X1 D5039 ( .B2(D1415_Y), .B1(D1565_Y), .B0(D5040_Y),     .Y(D5039_Y), .A(D4885_Y));
KC_OAI31_X1 D5010 ( .B2(D3364_Y), .B1(D5023_Y), .B0(D5020_Y),     .Y(D5010_Y), .A(D5018_Y));
KC_OAI31_X1 D4997 ( .B2(D5002_Y), .B1(D3446_Y), .B0(D4868_Y),     .Y(D4997_Y), .A(D3484_Q));
KC_OAI31_X1 D4878 ( .B2(D4897_Y), .B1(D4871_Y), .B0(D4876_Y),     .Y(D4878_Y), .A(D4887_Y));
KC_OAI31_X1 D4781 ( .B2(D4819_Q), .B1(D3383_Q), .B0(D3385_Q),     .Y(D4781_Y), .A(D4826_Q));
KC_OAI31_X1 D4780 ( .B2(D4814_Y), .B1(D4813_Y), .B0(D4812_Y),     .Y(D4780_Y), .A(D4758_Y));
KC_OAI31_X1 D4761 ( .B2(D4768_Y), .B1(D4767_Y), .B0(D4762_Y),     .Y(D4761_Y), .A(D4811_Y));
KC_OAI31_X1 D4680 ( .B2(D4683_Y), .B1(D1622_Y), .B0(D4671_Y),     .Y(D4680_Y), .A(D1571_Y));
KC_OAI31_X1 D4445 ( .B2(D4414_Y), .B1(D4441_Y), .B0(D4280_Y),     .Y(D4445_Y), .A(D4303_Y));
KC_OAI31_X1 D4433 ( .B2(D6025_Y), .B1(D5834_Y), .B0(D5772_Y),     .Y(D4433_Y), .A(D4426_Y));
KC_OAI31_X1 D4432 ( .B2(D6025_Y), .B1(D5834_Y), .B0(D5772_Y),     .Y(D4432_Y), .A(D4426_Y));
KC_OAI31_X1 D4362 ( .B2(D4290_Y), .B1(D4371_Y), .B0(D4275_Y),     .Y(D4362_Y), .A(D5936_Y));
KC_OAI31_X1 D4314 ( .B2(D4277_Y), .B1(D5876_Y), .B0(D5888_Y),     .Y(D4314_Y), .A(D4287_Y));
KC_OAI31_X1 D4278 ( .B2(D213_Y), .B1(D4446_Y), .B0(D7474_Y),     .Y(D4278_Y), .A(D1591_Y));
KC_OAI31_X1 D4208 ( .B2(D4339_Y), .B1(D4304_Y), .B0(D1592_Y),     .Y(D4208_Y), .A(D4216_Y));
KC_OAI31_X1 D3998 ( .B2(D6794_Y), .B1(D169_Y), .B0(D1445_Y),     .Y(D3998_Y), .A(D6958_Y));
KC_OAI31_X1 D3997 ( .B2(D169_Y), .B1(D3992_Y), .B0(D3881_Y),     .Y(D3997_Y), .A(D5558_Y));
KC_OAI31_X1 D3996 ( .B2(D169_Y), .B1(D1445_Y), .B0(D3881_Y),     .Y(D3996_Y), .A(D6958_Y));
KC_OAI31_X1 D3995 ( .B2(D169_Y), .B1(D1444_Y), .B0(D3881_Y),     .Y(D3995_Y), .A(D5558_Y));
KC_OAI31_X1 D3994 ( .B2(D169_Y), .B1(D3991_Y), .B0(D3881_Y),     .Y(D3994_Y), .A(D5558_Y));
KC_OAI31_X1 D3990 ( .B2(D6794_Y), .B1(D169_Y), .B0(D3991_Y),     .Y(D3990_Y), .A(D6958_Y));
KC_OAI31_X1 D3989 ( .B2(D6794_Y), .B1(D169_Y), .B0(D1444_Y),     .Y(D3989_Y), .A(D6958_Y));
KC_OAI31_X1 D3988 ( .B2(D6794_Y), .B1(D169_Y), .B0(D3992_Y),     .Y(D3988_Y), .A(D6958_Y));
KC_OAI31_X1 D3847 ( .B2(D6794_Y), .B1(D5387_Y), .B0(D3850_Y),     .Y(D3847_Y), .A(D3862_Y));
KC_OAI31_X1 D3846 ( .B2(D6794_Y), .B1(D5387_Y), .B0(D3838_Y),     .Y(D3846_Y), .A(D3862_Y));
KC_OAI31_X1 D3844 ( .B2(D5387_Y), .B1(D3850_Y), .B0(D3881_Y),     .Y(D3844_Y), .A(D3862_Y));
KC_OAI31_X1 D3843 ( .B2(D5387_Y), .B1(D3837_Y), .B0(D3881_Y),     .Y(D3843_Y), .A(D3862_Y));
KC_OAI31_X1 D3842 ( .B2(D6794_Y), .B1(D5387_Y), .B0(D3837_Y),     .Y(D3842_Y), .A(D3862_Y));
KC_OAI31_X1 D3835 ( .B2(D6794_Y), .B1(D5387_Y), .B0(D3851_Y),     .Y(D3835_Y), .A(D3862_Y));
KC_OAI31_X1 D3832 ( .B2(D5387_Y), .B1(D3838_Y), .B0(D3881_Y),     .Y(D3832_Y), .A(D3862_Y));
KC_OAI31_X1 D3709 ( .B2(D6794_Y), .B1(D11308_Y), .B0(D3717_Y),     .Y(D3709_Y), .A(D5215_Y));
KC_OAI31_X1 D3715 ( .B2(D11308_Y), .B1(D3714_Y), .B0(D3881_Y),     .Y(D3715_Y), .A(D5215_Y));
KC_OAI31_X1 D3710 ( .B2(D11308_Y), .B1(D3717_Y), .B0(D3881_Y),     .Y(D3710_Y), .A(D5215_Y));
KC_OAI31_X1 D3708 ( .B2(D6794_Y), .B1(D11308_Y), .B0(D3714_Y),     .Y(D3708_Y), .A(D5215_Y));
KC_OAI31_X1 D3658 ( .B2(D6794_Y), .B1(D11308_Y), .B0(D3716_Y),     .Y(D3658_Y), .A(D5215_Y));
KC_OAI31_X1 D3657 ( .B2(D11308_Y), .B1(D1412_Y), .B0(D3881_Y),     .Y(D3657_Y), .A(D5215_Y));
KC_OAI31_X1 D3656 ( .B2(D11308_Y), .B1(D3716_Y), .B0(D3881_Y),     .Y(D3656_Y), .A(D5215_Y));
KC_OAI31_X1 D3655 ( .B2(D6794_Y), .B1(D11308_Y), .B0(D1412_Y),     .Y(D3655_Y), .A(D5215_Y));
KC_OAI31_X1 D3541 ( .B2(D3400_Y), .B1(D3501_Y), .B0(D3548_Y),     .Y(D3541_Y), .A(D491_Y));
KC_OAI31_X1 D3536 ( .B2(D3388_Q), .B1(D3509_Y), .B0(D3574_Y),     .Y(D3536_Y), .A(D3499_Y));
KC_OAI31_X1 D3500 ( .B2(D5047_Y), .B1(D3634_Y), .B0(D3542_Y),     .Y(D3500_Y), .A(D3510_Y));
KC_OAI31_X1 D3449 ( .B2(D3388_Q), .B1(D3439_Y), .B0(D3475_Y),     .Y(D3449_Y), .A(D3429_Y));
KC_OAI31_X1 D3404 ( .B2(D3498_Y), .B1(D4911_Y), .B0(D3502_Y),     .Y(D3404_Y), .A(D3415_Y));
KC_OAI31_X1 D3403 ( .B2(D5012_Y), .B1(D3437_Y), .B0(D3404_Y),     .Y(D3403_Y), .A(D4887_Y));
KC_OAI31_X1 D3335 ( .B2(D3321_Y), .B1(D3398_Y), .B0(D1424_Y),     .Y(D3335_Y), .A(D4764_Y));
KC_OAI31_X1 D3334 ( .B2(D405_Y), .B1(D3361_Y), .B0(D3361_Y),     .Y(D3334_Y), .A(D4797_Y));
KC_OAI31_X1 D3220 ( .B2(D371_Y), .B1(D3277_Y), .B0(D3248_Y),     .Y(D3220_Y), .A(D3251_Y));
KC_OAI31_X1 D3217 ( .B2(D3204_Y), .B1(D3204_Y), .B0(D3204_Y),     .Y(D3217_Y), .A(D1469_Y));
KC_OAI31_X1 D3154 ( .B2(D3136_Y), .B1(D1457_Y), .B0(D3151_Y),     .Y(D3154_Y), .A(D1623_Y));
KC_OAI31_X1 D3153 ( .B2(D3127_Y), .B1(D4575_Y), .B0(D3096_Y),     .Y(D3153_Y), .A(D3095_Y));
KC_OAI31_X1 D3035 ( .B2(D3050_Y), .B1(D1771_Y), .B0(D3050_Y),     .Y(D3035_Y), .A(D3011_Y));
KC_OAI31_X1 D3009 ( .B2(D1516_Q), .B1(D3016_Y), .B0(D3013_Y),     .Y(D3009_Y), .A(D3030_Y));
KC_OAI31_X1 D2949 ( .B2(D2908_Y), .B1(D1489_Y), .B0(D2927_Y),     .Y(D2949_Y), .A(D2967_Y));
KC_OAI31_X1 D2913 ( .B2(D2988_Y), .B1(D2916_Y), .B0(D2918_Y),     .Y(D2913_Y), .A(D2961_Y));
KC_OAI31_X1 D2912 ( .B2(D2908_Y), .B1(D2988_Y), .B0(D2915_Y),     .Y(D2912_Y), .A(D2964_Y));
KC_OAI31_X1 D2909 ( .B2(D15_Y), .B1(D5_Y), .B0(D3008_Y), .Y(D2909_Y),     .A(D582_Y));
KC_OAI31_X1 D2905 ( .B2(D1489_Y), .B1(D2916_Y), .B0(D2917_Y),     .Y(D2905_Y), .A(D2960_Y));
KC_OAI31_X1 D2824 ( .B2(D2750_Y), .B1(D2826_Y), .B0(D2775_Y),     .Y(D2824_Y), .A(D2857_Y));
KC_OAI31_X1 D2763 ( .B2(D2799_Q), .B1(D2798_Q), .B0(D2845_Y),     .Y(D2763_Y), .A(D2813_Y));
KC_OAI31_X1 D2377 ( .B2(D12757_Y), .B1(D12720_Y), .B0(D12195_Y),     .Y(D2377_Y), .A(D13257_Y));
KC_OAI31_X1 D2364 ( .B2(D2361_Y), .B1(D12757_Y), .B0(D12195_Y),     .Y(D2364_Y), .A(D13257_Y));
KC_OAI31_X1 D2233 ( .B2(D11192_Y), .B1(D10790_Q), .B0(D10770_Y),     .Y(D2233_Y), .A(D11189_Y));
KC_OAI31_X1 D2203 ( .B2(D10858_Y), .B1(D2221_Q), .B0(D10770_Y),     .Y(D2203_Y), .A(D2201_Y));
KC_OAI31_X1 D1884 ( .B2(D1886_Y), .B1(D7179_Y), .B0(D7283_Y),     .Y(D1884_Y), .A(D7194_Y));
KC_OAI31_X1 D1741 ( .B2(D6234_Y), .B1(D6245_Y), .B0(D6252_Y),     .Y(D1741_Y), .A(D6246_Y));
KC_OAI31_X1 D1730 ( .B2(D4351_Y), .B1(D1754_Y), .B0(D7191_Y),     .Y(D1730_Y), .A(D5804_Y));
KC_OAI31_X1 D1729 ( .B2(D5913_Y), .B1(D5731_Y), .B0(D5796_Y),     .Y(D1729_Y), .A(D5804_Y));
KC_OAI31_X1 D1594 ( .B2(D1586_Y), .B1(D6_Y), .B0(D4442_Y), .Y(D1594_Y),     .A(D1591_Y));
KC_OAI31_X1 D1593 ( .B2(D5827_Y), .B1(D4513_Y), .B0(D4481_Y),     .Y(D1593_Y), .A(D4514_Y));
KC_OAI31_X1 D1443 ( .B2(D3477_Y), .B1(D3509_Y), .B0(D1446_Y),     .Y(D1443_Y), .A(D3452_Y));
KC_OAI31_X1 D1338 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11566_Y),     .Y(D1338_Y), .A(D11536_Y));
KC_OAI31_X1 D1267 ( .B2(D1823_Y), .B1(D2243_Y), .B0(D11565_Y),     .Y(D1267_Y), .A(D11536_Y));
KC_OAI31_X1 D1184 ( .B2(D13715_Y), .B1(D13729_Y), .B0(D13987_Y),     .Y(D1184_Y), .A(D13741_Y));
KC_OAI31_X1 D1176 ( .B2(D11492_Y), .B1(D8589_Q), .B0(D8551_Y),     .Y(D1176_Y), .A(D1172_Y));
KC_OAI31_X1 D985 ( .B2(D1049_Y), .B1(D14021_Y), .B0(D1155_Q),     .Y(D985_Y), .A(D14965_Y));
KC_OAI31_X1 D983 ( .B2(D8477_Y), .B1(D903_Q), .B0(D10770_Y),     .Y(D983_Y), .A(D6875_Y));
KC_OAI31_X1 D960 ( .B2(D6781_Y), .B1(D6826_Q), .B0(D10770_Y),     .Y(D960_Y), .A(D8285_Y));
KC_OAI31_X1 D869 ( .B2(D6788_Y), .B1(D6744_Q), .B0(D8060_Y),     .Y(D869_Y), .A(D8349_Y));
KC_OAI31_X1 D868 ( .B2(D11842_Y), .B1(D11859_Q), .B0(D11259_Y),     .Y(D868_Y), .A(D867_Y));
KC_OAI31_X1 D862 ( .B2(D6794_Y), .B1(D6777_Y), .B0(D6780_Y),     .Y(D862_Y), .A(D5391_Y));
KC_OAI31_X1 D861 ( .B2(D5387_Y), .B1(D3851_Y), .B0(D3881_Y),     .Y(D861_Y), .A(D3862_Y));
KC_OAI31_X1 D860 ( .B2(D6794_Y), .B1(D6777_Y), .B0(D6784_Y),     .Y(D860_Y), .A(D5391_Y));
KC_OAI31_X1 D743 ( .B2(D10741_Y), .B1(D10791_Q), .B0(D10770_Y),     .Y(D743_Y), .A(D10737_Y));
KC_OAI31_X1 D738 ( .B2(D6711_Y), .B1(D789_Q), .B0(D8060_Y), .Y(D738_Y),     .A(D8196_Y));
KC_OAI31_X1 D631 ( .B2(D10861_Y), .B1(D11322_Y), .B0(D11143_Y),     .Y(D631_Y), .A(D11258_Y));
KC_OAI31_X1 D561 ( .B2(D9371_Y), .B1(D2042_Y), .B0(D9365_Y),     .Y(D561_Y), .A(D8029_Y));
KC_OAI31_X1 D553 ( .B2(D12202_Y), .B1(D392_Y), .B0(D6287_Y),     .Y(D553_Y), .A(D11655_Y));
KC_OAI31_X1 D253 ( .B2(D7349_Y), .B1(D7366_Y), .B0(D5924_Y),     .Y(D253_Y), .A(D7319_Y));
KC_OAI31_X1 D217 ( .B2(D5973_Y), .B1(D1735_Y), .B0(D219_Y), .Y(D217_Y),     .A(D1591_Y));
KC_OAI31_X1 D78 ( .B2(D2230_Y), .B1(D11541_Q), .B0(D8551_Y), .Y(D78_Y),     .A(D2180_Y));
KC_AOI31_X1 D16560 ( .B0(D1381_Q), .B1(D16539_Y), .B2(D16528_Y),     .Y(D16560_Y), .A(D16541_Y));
KC_AOI31_X1 D16527 ( .B0(D16512_Y), .B1(D16501_Y), .B2(D16506_Y),     .Y(D16527_Y), .A(D16496_Y));
KC_AOI31_X1 D16526 ( .B0(D16512_Y), .B1(D16503_Y), .B2(D16494_Y),     .Y(D16526_Y), .A(D16496_Y));
KC_AOI31_X1 D16440 ( .B0(D16470_Q), .B1(D1324_Q), .B2(D16456_Y),     .Y(D16440_Y), .A(D16372_Y));
KC_AOI31_X1 D16420 ( .B0(D16419_Y), .B1(D16414_Y), .B2(D16443_Y),     .Y(D16420_Y), .A(D16421_Y));
KC_AOI31_X1 D16410 ( .B0(D16459_Q), .B1(D16441_Y), .B2(D16444_Y),     .Y(D16410_Y), .A(D1281_Y));
KC_AOI31_X1 D16409 ( .B0(D16411_Y), .B1(D16461_Y), .B2(D1273_Y),     .Y(D16409_Y), .A(D16407_Y));
KC_AOI31_X1 D16406 ( .B0(D16453_Y), .B1(D16429_Y), .B2(D16460_Y),     .Y(D16406_Y), .A(D16407_Y));
KC_AOI31_X1 D16262 ( .B0(D16252_Y), .B1(D2657_Y), .B2(D16227_Y),     .Y(D16262_Y), .A(D16260_Y));
KC_AOI31_X1 D16258 ( .B0(D2657_Y), .B1(D16283_Y), .B2(D16299_Y),     .Y(D16258_Y), .A(D16260_Y));
KC_AOI31_X1 D16252 ( .B0(D16289_Q), .B1(D16281_Y), .B2(D15630_Y),     .Y(D16252_Y), .A(D16269_Y));
KC_AOI31_X1 D15462 ( .B0(D14813_Y), .B1(D2604_Y), .B2(D9085_Y),     .Y(D15462_Y), .A(D15593_Y));
KC_AOI31_X1 D15340 ( .B0(D15522_Y), .B1(D15349_Y), .B2(D8902_Y),     .Y(D15340_Y), .A(D15458_Y));
KC_AOI31_X1 D15281 ( .B0(D16088_Y), .B1(D15282_Y), .B2(D15290_Y),     .Y(D15281_Y), .A(D2629_Y));
KC_AOI31_X1 D14848 ( .B0(D14788_Q), .B1(D14789_Q), .B2(D14787_Q),     .Y(D14848_Y), .A(D13982_Y));
KC_AOI31_X1 D14617 ( .B0(D640_Y), .B1(D14648_Y), .B2(D14744_Y),     .Y(D14617_Y), .A(D13934_Y));
KC_AOI31_X1 D14616 ( .B0(D14686_Q), .B1(D647_Y), .B2(D14622_Y),     .Y(D14616_Y), .A(D14663_Y));
KC_AOI31_X1 D14613 ( .B0(D14715_Y), .B1(D644_Y), .B2(D14614_Y),     .Y(D14613_Y), .A(D13934_Y));
KC_AOI31_X1 D14612 ( .B0(D13931_Y), .B1(D640_Y), .B2(D644_Y),     .Y(D14612_Y), .A(D13934_Y));
KC_AOI31_X1 D14611 ( .B0(D14776_Y), .B1(D14715_Y), .B2(D14669_Y),     .Y(D14611_Y), .A(D13934_Y));
KC_AOI31_X1 D14123 ( .B0(D14837_Y), .B1(D14292_Y), .B2(D14124_Y),     .Y(D14123_Y), .A(D14047_Y));
KC_AOI31_X1 D13931 ( .B0(D573_Y), .B1(D13930_Y), .B2(D13936_Y),     .Y(D13931_Y), .A(D13972_Y));
KC_AOI31_X1 D13562 ( .B0(D12951_Y), .B1(D14196_Q), .B2(D12955_Y),     .Y(D13562_Y), .A(D12905_Y));
KC_AOI31_X1 D13452 ( .B0(D13468_Y), .B1(D12887_Y), .B2(D852_Q),     .Y(D13452_Y), .A(D13461_Y));
KC_AOI31_X1 D13351 ( .B0(D12694_Y), .B1(D14024_Y), .B2(D12797_Y),     .Y(D13351_Y), .A(D13364_Y));
KC_AOI31_X1 D13341 ( .B0(D12694_Y), .B1(D844_Y), .B2(D13372_Y),     .Y(D13341_Y), .A(D13364_Y));
KC_AOI31_X1 D13223 ( .B0(D13220_Y), .B1(D13225_Y), .B2(D13228_Y),     .Y(D13223_Y), .A(D12751_Y));
KC_AOI31_X1 D12796 ( .B0(D12820_Y), .B1(D12786_Y), .B2(D12864_Y),     .Y(D12796_Y), .A(D13392_Y));
KC_AOI31_X1 D12723 ( .B0(D13220_Y), .B1(D12718_Y), .B2(D13227_Y),     .Y(D12723_Y), .A(D12751_Y));
KC_AOI31_X1 D12709 ( .B0(D12719_Y), .B1(D13220_Y), .B2(D13228_Y),     .Y(D12709_Y), .A(D12751_Y));
KC_AOI31_X1 D12203 ( .B0(D10177_Y), .B1(D11657_Y), .B2(D11677_Y),     .Y(D12203_Y), .A(D1954_Y));
KC_AOI31_X1 D9531 ( .B0(D9576_Q), .B1(D9526_Y), .B2(D9521_Y),     .Y(D9531_Y), .A(D826_Q));
KC_AOI31_X1 D9416 ( .B0(D625_Y), .B1(D9486_Y), .B2(D9425_Y),     .Y(D9416_Y), .A(D7153_Y));
KC_AOI31_X1 D9172 ( .B0(D9221_Q), .B1(D9220_Q), .B2(D9174_Y),     .Y(D9172_Y), .A(D4526_Y));
KC_AOI31_X1 D9123 ( .B0(D9136_Y), .B1(D383_Y), .B2(D9121_Y),     .Y(D9123_Y), .A(D15450_Y));
KC_AOI31_X1 D9073 ( .B0(D9084_Y), .B1(D9053_Y), .B2(D7560_Y),     .Y(D9073_Y), .A(D7361_Y));
KC_AOI31_X1 D9070 ( .B0(D9081_Y), .B1(D9065_Y), .B2(D7540_Y),     .Y(D9070_Y), .A(D7361_Y));
KC_AOI31_X1 D9047 ( .B0(D340_Y), .B1(D9039_Y), .B2(D7552_Y),     .Y(D9047_Y), .A(D7361_Y));
KC_AOI31_X1 D9042 ( .B0(D9034_Y), .B1(D9124_Y), .B2(D9038_Y),     .Y(D9042_Y), .A(D7361_Y));
KC_AOI31_X1 D8406 ( .B0(D8405_Y), .B1(D8384_Y), .B2(D8414_Y),     .Y(D8406_Y), .A(D8476_Y));
KC_AOI31_X1 D8283 ( .B0(D8282_Y), .B1(D8282_Y), .B2(D8282_Y),     .Y(D8283_Y), .A(D8338_Y));
KC_AOI31_X1 D8085 ( .B0(D8087_Y), .B1(D9407_Y), .B2(D8242_Y),     .Y(D8085_Y), .A(D8084_Y));
KC_AOI31_X1 D7914 ( .B0(D1901_Y), .B1(D7912_Y), .B2(D7940_Y),     .Y(D7914_Y), .A(D6431_Y));
KC_AOI31_X1 D7687 ( .B0(D7681_Y), .B1(D7697_Y), .B2(D7728_Y),     .Y(D7687_Y), .A(D6027_Y));
KC_AOI31_X1 D7637 ( .B0(D5966_Y), .B1(D7319_Y), .B2(D4515_Y),     .Y(D7637_Y), .A(D7632_Y));
KC_AOI31_X1 D7634 ( .B0(D386_Q), .B1(D385_Q), .B2(D7633_Y),     .Y(D7634_Y), .A(D7496_Y));
KC_AOI31_X1 D7624 ( .B0(D7689_Y), .B1(D7678_Y), .B2(D6095_Y),     .Y(D7624_Y), .A(D386_Q));
KC_AOI31_X1 D7509 ( .B0(D7506_Y), .B1(D7634_Y), .B2(D1871_Y),     .Y(D7509_Y), .A(D8971_Y));
KC_AOI31_X1 D7502 ( .B0(D7506_Y), .B1(D275_Y), .B2(D7634_Y),     .Y(D7502_Y), .A(D282_Y));
KC_AOI31_X1 D7497 ( .B0(D6090_Y), .B1(D6026_Y), .B2(D6075_Y),     .Y(D7497_Y), .A(D9147_Y));
KC_AOI31_X1 D7424 ( .B0(D179_Y), .B1(D6061_Y), .B2(D6021_Y),     .Y(D7424_Y), .A(D285_Y));
KC_AOI31_X1 D7415 ( .B0(D726_Y), .B1(D5978_Y), .B2(D1962_Y),     .Y(D7415_Y), .A(D7475_Q));
KC_AOI31_X1 D7220 ( .B0(D7205_Y), .B1(D8752_Y), .B2(D7228_Y),     .Y(D7220_Y), .A(D7303_Y));
KC_AOI31_X1 D7219 ( .B0(D7188_Y), .B1(D7209_Y), .B2(D7172_Y),     .Y(D7219_Y), .A(D7301_Y));
KC_AOI31_X1 D7207 ( .B0(D7309_Y), .B1(D7175_Y), .B2(D7236_Y),     .Y(D7207_Y), .A(D7212_Y));
KC_AOI31_X1 D7200 ( .B0(D7206_Y), .B1(D8776_Y), .B2(D2053_Y),     .Y(D7200_Y), .A(D7201_Y));
KC_AOI31_X1 D7165 ( .B0(D9475_Y), .B1(D9481_Y), .B2(D7180_Y),     .Y(D7165_Y), .A(D6024_Y));
KC_AOI31_X1 D6836 ( .B0(D6889_Y), .B1(D8456_Y), .B2(D6880_Y),     .Y(D6836_Y), .A(D6843_Y));
KC_AOI31_X1 D6434 ( .B0(D5026_Y), .B1(D5030_Y), .B2(D6443_Y),     .Y(D6434_Y), .A(D6427_Y));
KC_AOI31_X1 D6233 ( .B0(D6252_Y), .B1(D1705_Y), .B2(D1705_Y),     .Y(D6233_Y), .A(D6245_Y));
KC_AOI31_X1 D6226 ( .B0(D6229_Y), .B1(D6283_Y), .B2(D6283_Y),     .Y(D6226_Y), .A(D6279_Y));
KC_AOI31_X1 D26 ( .B0(D6039_Y), .B1(D1712_Y), .B2(D6098_Y), .Y(D26_Y),     .A(D8995_Y));
KC_AOI31_X1 D6087 ( .B0(D6115_Y), .B1(D16143_Y), .B2(D7531_Y),     .Y(D6087_Y), .A(D6089_Y));
KC_AOI31_X1 D5960 ( .B0(D5955_Y), .B1(D6045_Y), .B2(D6063_Y),     .Y(D5960_Y), .A(D5972_Y));
KC_AOI31_X1 D5959 ( .B0(D6002_Y), .B1(D5987_Y), .B2(D1710_Y),     .Y(D5959_Y), .A(D6091_Y));
KC_AOI31_X1 D5878 ( .B0(D5877_Y), .B1(D5684_Y), .B2(D7984_Y),     .Y(D5878_Y), .A(D5644_Y));
KC_AOI31_X1 D5773 ( .B0(D5968_Y), .B1(D7242_Y), .B2(D7092_Y),     .Y(D5773_Y), .A(D5661_Y));
KC_AOI31_X1 D5772 ( .B0(D5686_Q), .B1(D7257_Y), .B2(D5773_Y),     .Y(D5772_Y), .A(D5650_Y));
KC_AOI31_X1 D5716 ( .B0(D5749_Y), .B1(D5727_Y), .B2(D5761_Y),     .Y(D5716_Y), .A(D7376_Y));
KC_AOI31_X1 D5342 ( .B0(D5295_Y), .B1(D5360_Y), .B2(D5369_Y),     .Y(D5342_Y), .A(D5383_Y));
KC_AOI31_X1 D5035 ( .B0(D1567_Y), .B1(D3576_Q), .B2(D4925_Y),     .Y(D5035_Y), .A(D1602_Y));
KC_AOI31_X1 D5034 ( .B0(D3576_Q), .B1(D4887_Y), .B2(D5037_Y),     .Y(D5034_Y), .A(D3410_Y));
KC_AOI31_X1 D5024 ( .B0(D5011_Y), .B1(D5032_Y), .B2(D5031_Y),     .Y(D5024_Y), .A(D5023_Y));
KC_AOI31_X1 D5013 ( .B0(D4897_Y), .B1(D3446_Y), .B2(D1563_Y),     .Y(D5013_Y), .A(D5074_Y));
KC_AOI31_X1 D5007 ( .B0(D3446_Y), .B1(D1563_Y), .B2(D4911_Y),     .Y(D5007_Y), .A(D5024_Y));
KC_AOI31_X1 D5006 ( .B0(D5009_Y), .B1(D4903_Y), .B2(D3576_Q),     .Y(D5006_Y), .A(D5064_Y));
KC_AOI31_X1 D4919 ( .B0(D3498_Y), .B1(D3388_Q), .B2(D4918_Y),     .Y(D4919_Y), .A(D4975_Y));
KC_AOI31_X1 D4904 ( .B0(D4877_Y), .B1(D3426_Y), .B2(D4964_Y),     .Y(D4904_Y), .A(D4944_Y));
KC_AOI31_X1 D4899 ( .B0(D4920_Y), .B1(D4952_Y), .B2(D4886_Y),     .Y(D4899_Y), .A(D4970_Y));
KC_AOI31_X1 D4884 ( .B0(D4883_Y), .B1(D4874_Y), .B2(D3431_Y),     .Y(D4884_Y), .A(D3456_Y));
KC_AOI31_X1 D4861 ( .B0(D4862_Y), .B1(D4935_Y), .B2(D3469_Y),     .Y(D4861_Y), .A(D4869_Y));
KC_AOI31_X1 D4860 ( .B0(D3498_Y), .B1(D4913_Y), .B2(D4867_Y),     .Y(D4860_Y), .A(D1604_Y));
KC_AOI31_X1 D4764 ( .B0(D9345_Y), .B1(D369_Y), .B2(D7818_Y),     .Y(D4764_Y), .A(D413_Y));
KC_AOI31_X1 D4750 ( .B0(D1567_Y), .B1(D4926_Y), .B2(D4960_Y),     .Y(D4750_Y), .A(D1568_Y));
KC_AOI31_X1 D4749 ( .B0(D1567_Y), .B1(D4920_Y), .B2(D4926_Y),     .Y(D4749_Y), .A(D1568_Y));
KC_AOI31_X1 D4654 ( .B0(D4712_Y), .B1(D4701_Y), .B2(D4701_Y),     .Y(D4654_Y), .A(D4701_Y));
KC_AOI31_X1 D4599 ( .B0(D4640_Q), .B1(D4591_Y), .B2(D4503_Y),     .Y(D4599_Y), .A(D4603_Y));
KC_AOI31_X1 D4596 ( .B0(D4681_Y), .B1(D4622_Y), .B2(D4611_Y),     .Y(D4596_Y), .A(D4504_Y));
KC_AOI31_X1 D4436 ( .B0(D4150_Y), .B1(D4427_Y), .B2(D4416_Y),     .Y(D4436_Y), .A(D4457_Y));
KC_AOI31_X1 D4351 ( .B0(D4336_Y), .B1(D4334_Y), .B2(D4342_Y),     .Y(D4351_Y), .A(D5867_Y));
KC_AOI31_X1 D4331 ( .B0(D4339_Y), .B1(D4316_Y), .B2(D4325_Y),     .Y(D4331_Y), .A(D4349_Y));
KC_AOI31_X1 D3440 ( .B0(D3441_Y), .B1(D4947_Y), .B2(D440_Y),     .Y(D3440_Y), .A(D4939_Y));
KC_AOI31_X1 D3424 ( .B0(D3423_Y), .B1(D3414_Y), .B2(D3427_Y),     .Y(D3424_Y), .A(D4899_Y));
KC_AOI31_X1 D3412 ( .B0(D4887_Y), .B1(D3498_Y), .B2(D3462_Y),     .Y(D3412_Y), .A(D3413_Y));
KC_AOI31_X1 D3411 ( .B0(D4889_Y), .B1(D3460_Y), .B2(D4888_Y),     .Y(D3411_Y), .A(D1537_Y));
KC_AOI31_X1 D3328 ( .B0(D4774_Y), .B1(D3241_Y), .B2(D3333_Y),     .Y(D3328_Y), .A(D7641_Y));
KC_AOI31_X1 D3316 ( .B0(D3397_Y), .B1(D4744_Y), .B2(D12135_Y),     .Y(D3316_Y), .A(D7641_Y));
KC_AOI31_X1 D3235 ( .B0(D3184_Q), .B1(D3349_Y), .B2(D3256_Y),     .Y(D3235_Y), .A(D3231_Y));
KC_AOI31_X1 D3227 ( .B0(D1456_Y), .B1(D3230_Y), .B2(D3253_Y),     .Y(D3227_Y), .A(D3284_Y));
KC_AOI31_X1 D3216 ( .B0(D3300_Y), .B1(D3243_Y), .B2(D3214_Y),     .Y(D3216_Y), .A(D7641_Y));
KC_AOI31_X1 D3210 ( .B0(D3211_Y), .B1(D12135_Y), .B2(D4710_Y),     .Y(D3210_Y), .A(D7641_Y));
KC_AOI31_X1 D3147 ( .B0(D4599_Y), .B1(D3018_Y), .B2(D366_Y),     .Y(D3147_Y), .A(D7641_Y));
KC_AOI31_X1 D3115 ( .B0(D3110_Y), .B1(D3197_Y), .B2(D3124_Y),     .Y(D3115_Y), .A(D7641_Y));
KC_AOI31_X1 D3109 ( .B0(D3106_Y), .B1(D3116_Y), .B2(D3114_Y),     .Y(D3109_Y), .A(D7641_Y));
KC_AOI31_X1 D3099 ( .B0(D3117_Y), .B1(D3103_Y), .B2(D4573_Y),     .Y(D3099_Y), .A(D7641_Y));
KC_AOI31_X1 D3032 ( .B0(D4525_Y), .B1(D3091_Y), .B2(D4627_Y),     .Y(D3032_Y), .A(D3045_Y));
KC_AOI31_X1 D2655 ( .B0(D16101_Y), .B1(D2675_Y), .B2(D16085_Y),     .Y(D2655_Y), .A(D16127_Y));
KC_AOI31_X1 D2411 ( .B0(D14477_Y), .B1(D13787_Y), .B2(D15220_Y),     .Y(D2411_Y), .A(D13668_Y));
KC_AOI31_X1 D2003 ( .B0(D407_Y), .B1(D10105_Y), .B2(D9193_Y),     .Y(D2003_Y), .A(D9194_Y));
KC_AOI31_X1 D1714 ( .B0(D5646_Y), .B1(D6072_Y), .B2(D5886_Y),     .Y(D1714_Y), .A(D7454_Y));
KC_AOI31_X1 D1707 ( .B0(D6092_Y), .B1(D5964_Y), .B2(D1749_Y),     .Y(D1707_Y), .A(D4284_Y));
KC_AOI31_X1 D1703 ( .B0(D1766_Y), .B1(D6234_Y), .B2(D6234_Y),     .Y(D1703_Y), .A(D1790_Y));
KC_AOI31_X1 D1575 ( .B0(D4595_Y), .B1(D4503_Y), .B2(D3243_Y),     .Y(D1575_Y), .A(D50_Y));
KC_AOI31_X1 D1538 ( .B0(D4091_Y), .B1(D2716_Y), .B2(D4106_Y),     .Y(D1538_Y), .A(D1653_Y));
KC_AOI31_X1 D1417 ( .B0(D3265_Y), .B1(D3266_Y), .B2(D3226_Y),     .Y(D1417_Y), .A(D3288_Y));
KC_AOI31_X1 D968 ( .B0(D11024_Y), .B1(D8364_Y), .B2(D8371_Y),     .Y(D968_Y), .A(D970_Y));
KC_AOI31_X1 D632 ( .B0(D12695_Y), .B1(D12718_Y), .B2(D13225_Y),     .Y(D632_Y), .A(D13364_Y));
KC_AOI31_X1 D627 ( .B0(D12768_Y), .B1(D13359_Y), .B2(D13385_Y),     .Y(D627_Y), .A(D13364_Y));
KC_AOI31_X1 D568 ( .B0(D16089_Y), .B1(D15262_Y), .B2(D16086_Y),     .Y(D568_Y), .A(D15337_Y));
KC_AOI31_X1 D281 ( .B0(D6028_Y), .B1(D5992_Y), .B2(D7441_Y),     .Y(D281_Y), .A(D7177_Y));
KC_AOI31_X1 D276 ( .B0(D5951_Y), .B1(D7504_Y), .B2(D6040_Y),     .Y(D276_Y), .A(D6028_Y));
KC_AOI31_X1 D215 ( .B0(D9482_Y), .B1(D7251_Y), .B2(D5657_Y),     .Y(D215_Y), .A(D5650_Y));
KC_AOI31_X1 D181 ( .B0(D7113_Y), .B1(D7114_Y), .B2(D8706_Y),     .Y(D181_Y), .A(D8708_Y));
KC_AOI31_X1 D71 ( .B0(D7501_Y), .B1(D7469_Y), .B2(D1904_Y), .Y(D71_Y),     .A(D6075_Y));
KC_NAND2_X1 D16694 ( .Y(D16694_Y), .B(D16671_Y), .A(D1395_Q));
KC_NAND2_X1 D16692 ( .Y(D16692_Y), .B(D16691_Y), .A(D16681_Q));
KC_NAND2_X1 D16690 ( .Y(D16690_Y), .B(D16689_Y), .A(D16682_Q));
KC_NAND2_X1 D16688 ( .Y(D16688_Y), .B(D16695_Y), .A(D16684_Q));
KC_NAND2_X1 D16670 ( .Y(D16670_Y), .B(D16643_Y), .A(D16650_Q));
KC_NAND2_X1 D16668 ( .Y(D16668_Y), .B(D16646_Y), .A(D1373_Q));
KC_NAND2_X1 D16666 ( .Y(D16666_Y), .B(D16669_Y), .A(D16660_Q));
KC_NAND2_X1 D16653 ( .Y(D16653_Y), .B(D1395_Q), .A(D16650_Q));
KC_NAND2_X1 D16642 ( .Y(D16642_Y), .B(D16640_Y), .A(D1396_Q));
KC_NAND2_X1 D16574 ( .Y(D16574_Y), .B(D16570_Y), .A(D16586_Y));
KC_NAND2_X1 D16573 ( .Y(D16573_Y), .B(D16382_Y), .A(D16285_Y));
KC_NAND2_X1 D16544 ( .Y(D16544_Y), .B(D16771_Y), .A(D1385_Q));
KC_NAND2_X1 D16542 ( .Y(D16542_Y), .B(D16557_Q), .A(D16543_Y));
KC_NAND2_X1 D16535 ( .Y(D16535_Y), .B(D16537_Y), .A(D16771_Y));
KC_NAND2_X1 D16531 ( .Y(D16531_Y), .B(D16550_Y), .A(D16551_Y));
KC_NAND2_X1 D16487 ( .Y(D16487_Y), .B(D16488_Y), .A(D16528_Y));
KC_NAND2_X1 D16485 ( .Y(D16485_Y), .B(D13988_Y), .A(D14651_Y));
KC_NAND2_X1 D16417 ( .Y(D16417_Y), .B(D16459_Q), .A(D1324_Q));
KC_NAND2_X1 D16408 ( .Y(D16408_Y), .B(D13966_Y), .A(D16430_Y));
KC_NAND2_X1 D16375 ( .Y(D16375_Y), .B(D16438_Y), .A(D16425_Y));
KC_NAND2_X1 D16374 ( .Y(D16374_Y), .B(D16299_Y), .A(D16399_Q));
KC_NAND2_X1 D16264 ( .Y(D16264_Y), .B(D16259_Y), .A(D16272_Y));
KC_NAND2_X1 D16253 ( .Y(D16253_Y), .B(D16268_Y), .A(D16299_Y));
KC_NAND2_X1 D16251 ( .Y(D16251_Y), .B(D16268_Y), .A(D14057_Y));
KC_NAND2_X1 D16250 ( .Y(D16250_Y), .B(D15630_Y), .A(D16274_Y));
KC_NAND2_X1 D16247 ( .Y(D16247_Y), .B(D16273_Y), .A(D16293_Q));
KC_NAND2_X1 D16191 ( .Y(D16191_Y), .B(D16458_Y), .A(D16192_Y));
KC_NAND2_X1 D16187 ( .Y(D16187_Y), .B(D16095_Y), .A(D16148_Y));
KC_NAND2_X1 D16113 ( .Y(D16113_Y), .B(D16137_Y), .A(D14654_Y));
KC_NAND2_X1 D16112 ( .Y(D16112_Y), .B(D16170_Y), .A(D16131_Y));
KC_NAND2_X1 D16109 ( .Y(D16109_Y), .B(D16168_Y), .A(D16186_Y));
KC_NAND2_X1 D16100 ( .Y(D16100_Y), .B(D16120_Y), .A(D16051_Y));
KC_NAND2_X1 D16065 ( .Y(D16065_Y), .B(D16094_Y), .A(D16059_Y));
KC_NAND2_X1 D16058 ( .Y(D16058_Y), .B(D16043_Y), .A(D16094_Y));
KC_NAND2_X1 D16056 ( .Y(D16056_Y), .B(D16054_Y), .A(D16057_Y));
KC_NAND2_X1 D15917 ( .Y(D15917_Y), .B(D15936_S), .A(D15916_Y));
KC_NAND2_X1 D15916 ( .Y(D15916_Y), .B(D15961_Y), .A(D15994_Q));
KC_NAND2_X1 D15912 ( .Y(D15912_Y), .B(D15859_S), .A(D15904_Y));
KC_NAND2_X1 D15908 ( .Y(D15908_Y), .B(D15897_Y), .A(D15948_Q));
KC_NAND2_X1 D15904 ( .Y(D15904_Y), .B(D15882_Y), .A(D16010_Q));
KC_NAND2_X1 D15901 ( .Y(D15901_Y), .B(D15856_S), .A(D15894_Y));
KC_NAND2_X1 D15898 ( .Y(D15898_Y), .B(D15888_Y), .A(D15947_Q));
KC_NAND2_X1 D15894 ( .Y(D15894_Y), .B(D15883_Y), .A(D16388_Q));
KC_NAND2_X1 D15893 ( .Y(D15893_Y), .B(D15858_S), .A(D15898_Y));
KC_NAND2_X1 D15638 ( .Y(D15638_Y), .B(D15637_Y), .A(D15628_Y));
KC_NAND2_X1 D15637 ( .Y(D15637_Y), .B(D14827_Y), .A(D15496_Y));
KC_NAND2_X1 D15636 ( .Y(D15636_Y), .B(D749_Y), .A(D15633_Y));
KC_NAND2_X1 D15627 ( .Y(D15627_Y), .B(D15618_Y), .A(D15467_Y));
KC_NAND2_X1 D15626 ( .Y(D15626_Y), .B(D15495_Y), .A(D14826_Y));
KC_NAND2_X1 D15625 ( .Y(D15625_Y), .B(D15620_Y), .A(D15628_Y));
KC_NAND2_X1 D15619 ( .Y(D15619_Y), .B(D15003_Y), .A(D16461_Y));
KC_NAND2_X1 D15618 ( .Y(D15618_Y), .B(D15076_Y), .A(D16461_Y));
KC_NAND2_X1 D15609 ( .Y(D15609_Y), .B(D15580_Y), .A(D15577_Y));
KC_NAND2_X1 D15534 ( .Y(D15534_Y), .B(D15362_Y), .A(D15530_Y));
KC_NAND2_X1 D15530 ( .Y(D15530_Y), .B(D15345_Y), .A(D16461_Y));
KC_NAND2_X1 D15525 ( .Y(D15525_Y), .B(D15494_Y), .A(D15388_Y));
KC_NAND2_X1 D15524 ( .Y(D15524_Y), .B(D15803_Y), .A(D15563_Y));
KC_NAND2_X1 D15523 ( .Y(D15523_Y), .B(D15386_Y), .A(D15493_Y));
KC_NAND2_X1 D15517 ( .Y(D15517_Y), .B(D15507_Y), .A(D15387_Y));
KC_NAND2_X1 D15507 ( .Y(D15507_Y), .B(D14390_Y), .A(D16461_Y));
KC_NAND2_X1 D15502 ( .Y(D15502_Y), .B(D16242_Q), .A(D15476_Y));
KC_NAND2_X1 D15496 ( .Y(D15496_Y), .B(D15449_Y), .A(D14813_Y));
KC_NAND2_X1 D15495 ( .Y(D15495_Y), .B(D8885_Y), .A(D14813_Y));
KC_NAND2_X1 D15494 ( .Y(D15494_Y), .B(D15955_Y), .A(D16461_Y));
KC_NAND2_X1 D15493 ( .Y(D15493_Y), .B(D2647_Y), .A(D16461_Y));
KC_NAND2_X1 D15492 ( .Y(D15492_Y), .B(D651_Y), .A(D14813_Y));
KC_NAND2_X1 D15487 ( .Y(D15487_Y), .B(D16270_Y), .A(D1273_Y));
KC_NAND2_X1 D15483 ( .Y(D15483_Y), .B(D15482_Y), .A(D2607_Y));
KC_NAND2_X1 D15482 ( .Y(D15482_Y), .B(D14514_Y), .A(D15463_Y));
KC_NAND2_X1 D15475 ( .Y(D15475_Y), .B(D816_Q), .A(D16242_Q));
KC_NAND2_X1 D15470 ( .Y(D15470_Y), .B(D749_Y), .A(D15465_Y));
KC_NAND2_X1 D15469 ( .Y(D15469_Y), .B(D12140_Y), .A(D14720_Y));
KC_NAND2_X1 D15468 ( .Y(D15468_Y), .B(D15482_Y), .A(D14719_Y));
KC_NAND2_X1 D15467 ( .Y(D15467_Y), .B(D16198_Y), .A(D14813_Y));
KC_NAND2_X1 D15466 ( .Y(D15466_Y), .B(D15473_Y), .A(D15465_Y));
KC_NAND2_X1 D15465 ( .Y(D15465_Y), .B(D15463_Y), .A(D14720_Y));
KC_NAND2_X1 D15461 ( .Y(D15461_Y), .B(D636_Y), .A(D15513_Y));
KC_NAND2_X1 D15403 ( .Y(D15403_Y), .B(D15517_Y), .A(D15353_Y));
KC_NAND2_X1 D15394 ( .Y(D15394_Y), .B(D16125_Y), .A(D14654_Y));
KC_NAND2_X1 D15392 ( .Y(D15392_Y), .B(D2590_Y), .A(D15405_Y));
KC_NAND2_X1 D15391 ( .Y(D15391_Y), .B(D2590_Y), .A(D15406_Y));
KC_NAND2_X1 D15389 ( .Y(D15389_Y), .B(D2589_Y), .A(D15409_Y));
KC_NAND2_X1 D15388 ( .Y(D15388_Y), .B(D15433_Y), .A(D15522_Y));
KC_NAND2_X1 D15387 ( .Y(D15387_Y), .B(D6975_Y), .A(D15522_Y));
KC_NAND2_X1 D15386 ( .Y(D15386_Y), .B(D6977_Y), .A(D15522_Y));
KC_NAND2_X1 D15385 ( .Y(D15385_Y), .B(D16139_Y), .A(D15522_Y));
KC_NAND2_X1 D15384 ( .Y(D15384_Y), .B(D6524_Y), .A(D15522_Y));
KC_NAND2_X1 D15383 ( .Y(D15383_Y), .B(D2589_Y), .A(D15327_Y));
KC_NAND2_X1 D15382 ( .Y(D15382_Y), .B(D2589_Y), .A(D15397_Y));
KC_NAND2_X1 D15379 ( .Y(D15379_Y), .B(D15441_Y), .A(D16107_Y));
KC_NAND2_X1 D15376 ( .Y(D15376_Y), .B(D15373_Y), .A(D15363_Y));
KC_NAND2_X1 D15375 ( .Y(D15375_Y), .B(D12214_Y), .A(D15377_Y));
KC_NAND2_X1 D15374 ( .Y(D15374_Y), .B(D15371_Y), .A(D15377_Y));
KC_NAND2_X1 D15373 ( .Y(D15373_Y), .B(D14513_Y), .A(D15371_Y));
KC_NAND2_X1 D15364 ( .Y(D15364_Y), .B(D15366_Y), .A(D636_Y));
KC_NAND2_X1 D15363 ( .Y(D15363_Y), .B(D14624_Y), .A(D15377_Y));
KC_NAND2_X1 D15362 ( .Y(D15362_Y), .B(D636_Y), .A(D15374_Y));
KC_NAND2_X1 D15361 ( .Y(D15361_Y), .B(D15344_Y), .A(D15374_Y));
KC_NAND2_X1 D15351 ( .Y(D15351_Y), .B(D15514_Y), .A(D15353_Y));
KC_NAND2_X1 D15350 ( .Y(D15350_Y), .B(D15373_Y), .A(D15530_Y));
KC_NAND2_X1 D15310 ( .Y(D15310_Y), .B(D15283_Y), .A(D15326_Y));
KC_NAND2_X1 D15306 ( .Y(D15306_Y), .B(D567_Y), .A(D15282_Y));
KC_NAND2_X1 D15299 ( .Y(D15299_Y), .B(D15305_Y), .A(D15284_Y));
KC_NAND2_X1 D15298 ( .Y(D15298_Y), .B(D15304_Y), .A(D15284_Y));
KC_NAND2_X1 D15294 ( .Y(D15294_Y), .B(D2590_Y), .A(D15303_Y));
KC_NAND2_X1 D15293 ( .Y(D15293_Y), .B(D2590_Y), .A(D15301_Y));
KC_NAND2_X1 D15289 ( .Y(D15289_Y), .B(D2590_Y), .A(D16052_Y));
KC_NAND2_X1 D15279 ( .Y(D15279_Y), .B(D16053_Y), .A(D15320_Y));
KC_NAND2_X1 D15278 ( .Y(D15278_Y), .B(D15273_Y), .A(D15326_Y));
KC_NAND2_X1 D15277 ( .Y(D15277_Y), .B(D15283_Y), .A(D15309_Y));
KC_NAND2_X1 D15276 ( .Y(D15276_Y), .B(D15273_Y), .A(D15309_Y));
KC_NAND2_X1 D15271 ( .Y(D15271_Y), .B(D567_Y), .A(D15326_Y));
KC_NAND2_X1 D15270 ( .Y(D15270_Y), .B(D567_Y), .A(D15309_Y));
KC_NAND2_X1 D15267 ( .Y(D15267_Y), .B(D15273_Y), .A(D15282_Y));
KC_NAND2_X1 D15240 ( .Y(D15240_Y), .B(D15183_Y), .A(D15228_Y));
KC_NAND2_X1 D15096 ( .Y(D15096_Y), .B(D15070_S), .A(D15092_Y));
KC_NAND2_X1 D15092 ( .Y(D15092_Y), .B(D15094_Y), .A(D15133_Q));
KC_NAND2_X1 D15047 ( .Y(D15047_Y), .B(D15068_S), .A(D15046_Y));
KC_NAND2_X1 D15046 ( .Y(D15046_Y), .B(D2529_Y), .A(D2572_Q));
KC_NAND2_X1 D15014 ( .Y(D15014_Y), .B(D15072_S), .A(D15012_Y));
KC_NAND2_X1 D15012 ( .Y(D15012_Y), .B(D15099_Y), .A(D1158_Q));
KC_NAND2_X1 D14827 ( .Y(D14827_Y), .B(D14381_Y), .A(D15562_Y));
KC_NAND2_X1 D14826 ( .Y(D14826_Y), .B(D2579_Y), .A(D15562_Y));
KC_NAND2_X1 D14747 ( .Y(D14747_Y), .B(D14044_Y), .A(D14785_Y));
KC_NAND2_X1 D14744 ( .Y(D14744_Y), .B(D14664_Y), .A(D14044_Y));
KC_NAND2_X1 D14728 ( .Y(D14728_Y), .B(D14514_Y), .A(D12140_Y));
KC_NAND2_X1 D14719 ( .Y(D14719_Y), .B(D15490_Y), .A(D14720_Y));
KC_NAND2_X1 D14649 ( .Y(D14649_Y), .B(D13958_Y), .A(D13988_Y));
KC_NAND2_X1 D14646 ( .Y(D14646_Y), .B(D14587_Y), .A(D14655_Y));
KC_NAND2_X1 D14642 ( .Y(D14642_Y), .B(D15433_Y), .A(D2509_Y));
KC_NAND2_X1 D14641 ( .Y(D14641_Y), .B(D13952_Y), .A(D13997_Q));
KC_NAND2_X1 D14640 ( .Y(D14640_Y), .B(D13947_Y), .A(D14635_Y));
KC_NAND2_X1 D14639 ( .Y(D14639_Y), .B(D14644_Y), .A(D14742_Y));
KC_NAND2_X1 D14638 ( .Y(D14638_Y), .B(D2871_Y), .A(D2509_Y));
KC_NAND2_X1 D14637 ( .Y(D14637_Y), .B(D14673_Y), .A(D15499_Y));
KC_NAND2_X1 D14629 ( .Y(D14629_Y), .B(D14622_Y), .A(D14634_Y));
KC_NAND2_X1 D14628 ( .Y(D14628_Y), .B(D8889_Y), .A(D2509_Y));
KC_NAND2_X1 D14625 ( .Y(D14625_Y), .B(D14513_Y), .A(D12214_Y));
KC_NAND2_X1 D14621 ( .Y(D14621_Y), .B(D637_Y), .A(D14686_Q));
KC_NAND2_X1 D14620 ( .Y(D14620_Y), .B(D637_Y), .A(D722_Q));
KC_NAND2_X1 D14614 ( .Y(D14614_Y), .B(D14707_Y), .A(D14650_Y));
KC_NAND2_X1 D16770 ( .Y(D16770_Y), .B(D14609_Y), .A(D14519_Q));
KC_NAND2_X1 D14608 ( .Y(D14608_Y), .B(D14607_Y), .A(D14518_Q));
KC_NAND2_X1 D14606 ( .Y(D14606_Y), .B(D14605_Y), .A(D2512_Y));
KC_NAND2_X1 D14604 ( .Y(D14604_Y), .B(D14687_Q), .A(D14688_Q));
KC_NAND2_X1 D14602 ( .Y(D14602_Y), .B(D16769_Y), .A(D14601_Q));
KC_NAND2_X1 D14556 ( .Y(D14556_Y), .B(D14687_Q), .A(D14688_Q));
KC_NAND2_X1 D14541 ( .Y(D14541_Y), .B(D14539_Y), .A(D608_Q));
KC_NAND2_X1 D14534 ( .Y(D14534_Y), .B(D14576_Y), .A(D14519_Q));
KC_NAND2_X1 D14446 ( .Y(D14446_Y), .B(D15214_Q), .A(D14408_Y));
KC_NAND2_X1 D14141 ( .Y(D14141_Y), .B(D14023_Y), .A(D14026_Y));
KC_NAND2_X1 D14137 ( .Y(D14137_Y), .B(D14020_Y), .A(D14882_Y));
KC_NAND2_X1 D14134 ( .Y(D14134_Y), .B(D14020_Y), .A(D14879_Y));
KC_NAND2_X1 D14133 ( .Y(D14133_Y), .B(D14020_Y), .A(D14880_Y));
KC_NAND2_X1 D14132 ( .Y(D14132_Y), .B(D14020_Y), .A(D14881_Y));
KC_NAND2_X1 D14043 ( .Y(D14043_Y), .B(D14123_Y), .A(D14046_Y));
KC_NAND2_X1 D14024 ( .Y(D14024_Y), .B(D14025_Y), .A(D16275_Y));
KC_NAND2_X1 D14023 ( .Y(D14023_Y), .B(D12856_Q), .A(D13328_Y));
KC_NAND2_X1 D13962 ( .Y(D13962_Y), .B(D13996_Q), .A(D2461_Y));
KC_NAND2_X1 D13958 ( .Y(D13958_Y), .B(D2518_Q), .A(D13275_Q));
KC_NAND2_X1 D13953 ( .Y(D13953_Y), .B(D696_Q), .A(D13275_Q));
KC_NAND2_X1 D13952 ( .Y(D13952_Y), .B(D695_Q), .A(D13275_Q));
KC_NAND2_X1 D13948 ( .Y(D13948_Y), .B(D8902_Y), .A(D2509_Y));
KC_NAND2_X1 D13947 ( .Y(D13947_Y), .B(D13946_Y), .A(D13945_Y));
KC_NAND2_X1 D13940 ( .Y(D13940_Y), .B(D13941_Y), .A(D13930_Y));
KC_NAND2_X1 D13939 ( .Y(D13939_Y), .B(D14683_Y), .A(D14616_Y));
KC_NAND2_X1 D13935 ( .Y(D13935_Y), .B(D14665_Y), .A(D13275_Q));
KC_NAND2_X1 D13933 ( .Y(D13933_Y), .B(D13953_Y), .A(D13941_Y));
KC_NAND2_X1 D13924 ( .Y(D13924_Y), .B(D14603_Y), .A(D608_Q));
KC_NAND2_X1 D13922 ( .Y(D13922_Y), .B(D13925_Y), .A(D14520_Q));
KC_NAND2_X1 D13903 ( .Y(D13903_Y), .B(D13209_Q), .A(D13254_Y));
KC_NAND2_X1 D13900 ( .Y(D13900_Y), .B(D6977_Y), .A(D2509_Y));
KC_NAND2_X1 D13899 ( .Y(D13899_Y), .B(D12680_Q), .A(D13254_Y));
KC_NAND2_X1 D13898 ( .Y(D13898_Y), .B(D6524_Y), .A(D2509_Y));
KC_NAND2_X1 D13897 ( .Y(D13897_Y), .B(D16800_Y), .A(D2509_Y));
KC_NAND2_X1 D13889 ( .Y(D13889_Y), .B(D14000_Y), .A(D13928_Y));
KC_NAND2_X1 D13880 ( .Y(D13880_Y), .B(D12689_Q), .A(D13254_Y));
KC_NAND2_X1 D13875 ( .Y(D13875_Y), .B(D13211_Q), .A(D13254_Y));
KC_NAND2_X1 D13873 ( .Y(D13873_Y), .B(D13872_Q), .A(D13865_Q));
KC_NAND2_X1 D13871 ( .Y(D13871_Y), .B(D13874_Y), .A(D13864_Q));
KC_NAND2_X1 D13868 ( .Y(D13868_Y), .B(D13870_Y), .A(D543_Q));
KC_NAND2_X1 D13555 ( .Y(D13555_Y), .B(D2436_Y), .A(D13506_Y));
KC_NAND2_X1 D13554 ( .Y(D13554_Y), .B(D13543_Y), .A(D13506_Y));
KC_NAND2_X1 D13547 ( .Y(D13547_Y), .B(D13548_Y), .A(D13506_Y));
KC_NAND2_X1 D13546 ( .Y(D13546_Y), .B(D13567_Y), .A(D13506_Y));
KC_NAND2_X1 D13545 ( .Y(D13545_Y), .B(D2436_Y), .A(D13338_Y));
KC_NAND2_X1 D13542 ( .Y(D13542_Y), .B(D13553_Y), .A(D13578_Y));
KC_NAND2_X1 D13541 ( .Y(D13541_Y), .B(D13417_Y), .A(D13578_Y));
KC_NAND2_X1 D13536 ( .Y(D13536_Y), .B(D13393_Y), .A(D12754_Q));
KC_NAND2_X1 D13470 ( .Y(D13470_Y), .B(D13323_Y), .A(D7669_Y));
KC_NAND2_X1 D13456 ( .Y(D13456_Y), .B(D13468_Y), .A(D928_Q));
KC_NAND2_X1 D13455 ( .Y(D13455_Y), .B(D10216_Y), .A(D13460_Y));
KC_NAND2_X1 D13448 ( .Y(D13448_Y), .B(D13578_Y), .A(D2436_Y));
KC_NAND2_X1 D13447 ( .Y(D13447_Y), .B(D2438_Y), .A(D13553_Y));
KC_NAND2_X1 D13446 ( .Y(D13446_Y), .B(D13441_Y), .A(D13578_Y));
KC_NAND2_X1 D13445 ( .Y(D13445_Y), .B(D13458_Y), .A(D13464_Y));
KC_NAND2_X1 D13429 ( .Y(D13429_Y), .B(D2435_Y), .A(D13464_Y));
KC_NAND2_X1 D13428 ( .Y(D13428_Y), .B(D2438_Y), .A(D13464_Y));
KC_NAND2_X1 D13420 ( .Y(D13420_Y), .B(D2435_Y), .A(D13553_Y));
KC_NAND2_X1 D13419 ( .Y(D13419_Y), .B(D13409_Y), .A(D2432_Y));
KC_NAND2_X1 D13365 ( .Y(D13365_Y), .B(D13358_Y), .A(D13267_Q));
KC_NAND2_X1 D13356 ( .Y(D13356_Y), .B(D13347_Y), .A(D13353_Y));
KC_NAND2_X1 D13339 ( .Y(D13339_Y), .B(D13357_Y), .A(D13336_Y));
KC_NAND2_X1 D13334 ( .Y(D13334_Y), .B(D13475_Y), .A(D13328_Y));
KC_NAND2_X1 D13331 ( .Y(D13331_Y), .B(D13329_Y), .A(D12241_Y));
KC_NAND2_X1 D13330 ( .Y(D13330_Y), .B(D13327_Y), .A(D13335_Y));
KC_NAND2_X1 D13322 ( .Y(D13322_Y), .B(D2312_Y), .A(D2353_Y));
KC_NAND2_X1 D13321 ( .Y(D13321_Y), .B(D7670_Y), .A(D2353_Y));
KC_NAND2_X1 D13320 ( .Y(D13320_Y), .B(D13376_Y), .A(D16471_Q));
KC_NAND2_X1 D13319 ( .Y(D13319_Y), .B(D13256_Y), .A(D13315_Y));
KC_NAND2_X1 D13313 ( .Y(D13313_Y), .B(D13315_Y), .A(D161_Y));
KC_NAND2_X1 D13308 ( .Y(D13308_Y), .B(D2343_Y), .A(D13316_Y));
KC_NAND2_X1 D13301 ( .Y(D13301_Y), .B(D13317_Y), .A(D13316_Y));
KC_NAND2_X1 D13241 ( .Y(D13241_Y), .B(D13245_Y), .A(D13257_Y));
KC_NAND2_X1 D13240 ( .Y(D13240_Y), .B(D2390_Q), .A(D13254_Y));
KC_NAND2_X1 D13235 ( .Y(D13235_Y), .B(D13257_Y), .A(D10216_Y));
KC_NAND2_X1 D13224 ( .Y(D13224_Y), .B(D13257_Y), .A(D11276_Y));
KC_NAND2_X1 D13177 ( .Y(D13177_Y), .B(D13210_Q), .A(D13254_Y));
KC_NAND2_X1 D13176 ( .Y(D13176_Y), .B(D13203_Q), .A(D13254_Y));
KC_NAND2_X1 D16763 ( .Y(D16763_Y), .B(D13869_Y), .A(D13175_Q));
KC_NAND2_X1 D13019 ( .Y(D13019_Y), .B(D13539_Y), .A(D13578_Y));
KC_NAND2_X1 D13011 ( .Y(D13011_Y), .B(D13538_Y), .A(D13578_Y));
KC_NAND2_X1 D12950 ( .Y(D12950_Y), .B(D12991_Q), .A(D12952_Y));
KC_NAND2_X1 D12946 ( .Y(D12946_Y), .B(D12947_Y), .A(D13590_Y));
KC_NAND2_X1 D12894 ( .Y(D12894_Y), .B(D13469_Y), .A(D13696_Y));
KC_NAND2_X1 D12888 ( .Y(D12888_Y), .B(D14057_Y), .A(D14859_Y));
KC_NAND2_X1 D12887 ( .Y(D12887_Y), .B(D961_Y), .A(D843_Q));
KC_NAND2_X1 D12875 ( .Y(D12875_Y), .B(D961_Y), .A(D12854_Q));
KC_NAND2_X1 D12874 ( .Y(D12874_Y), .B(D961_Y), .A(D12749_Q));
KC_NAND2_X1 D12873 ( .Y(D12873_Y), .B(D961_Y), .A(D12857_Q));
KC_NAND2_X1 D12869 ( .Y(D12869_Y), .B(D14057_Y), .A(D15694_Y));
KC_NAND2_X1 D12825 ( .Y(D12825_Y), .B(D13402_Y), .A(D15474_Y));
KC_NAND2_X1 D12808 ( .Y(D12808_Y), .B(D12697_Y), .A(D14003_Y));
KC_NAND2_X1 D12807 ( .Y(D12807_Y), .B(D12792_Y), .A(D12697_Y));
KC_NAND2_X1 D12797 ( .Y(D12797_Y), .B(D12815_Y), .A(D12804_Y));
KC_NAND2_X1 D12793 ( .Y(D12793_Y), .B(D12773_Y), .A(D12856_Q));
KC_NAND2_X1 D12792 ( .Y(D12792_Y), .B(D13402_Y), .A(D15491_Y));
KC_NAND2_X1 D12791 ( .Y(D12791_Y), .B(D13402_Y), .A(D12788_Y));
KC_NAND2_X1 D12785 ( .Y(D12785_Y), .B(D12725_Y), .A(D12754_Q));
KC_NAND2_X1 D12784 ( .Y(D12784_Y), .B(D13402_Y), .A(D12787_Y));
KC_NAND2_X1 D12777 ( .Y(D12777_Y), .B(D12773_Y), .A(D12804_Y));
KC_NAND2_X1 D12771 ( .Y(D12771_Y), .B(D14057_Y), .A(D15583_Y));
KC_NAND2_X1 D12770 ( .Y(D12770_Y), .B(D14057_Y), .A(D14786_Y));
KC_NAND2_X1 D12760 ( .Y(D12760_Y), .B(D12751_Y), .A(D13234_Y));
KC_NAND2_X1 D12720 ( .Y(D12720_Y), .B(D12188_Y), .A(D7669_Y));
KC_NAND2_X1 D12717 ( .Y(D12717_Y), .B(D13226_Y), .A(D12731_Y));
KC_NAND2_X1 D12713 ( .Y(D12713_Y), .B(D7305_Y), .A(D12260_Y));
KC_NAND2_X1 D12711 ( .Y(D12711_Y), .B(D12791_Y), .A(D12697_Y));
KC_NAND2_X1 D12708 ( .Y(D12708_Y), .B(D13225_Y), .A(D12713_Y));
KC_NAND2_X1 D12702 ( .Y(D12702_Y), .B(D12825_Y), .A(D12697_Y));
KC_NAND2_X1 D12701 ( .Y(D12701_Y), .B(D12729_Y), .A(D699_Q));
KC_NAND2_X1 D12700 ( .Y(D12700_Y), .B(D12279_Q), .A(D12729_Y));
KC_NAND2_X1 D12699 ( .Y(D12699_Y), .B(D12697_Y), .A(D13950_Y));
KC_NAND2_X1 D12696 ( .Y(D12696_Y), .B(D12784_Y), .A(D12697_Y));
KC_NAND2_X1 D12661 ( .Y(D12661_Y), .B(D13216_Q), .A(D13275_Q));
KC_NAND2_X1 D12313 ( .Y(D12313_Y), .B(D12315_Y), .A(D14057_Y));
KC_NAND2_X1 D12199 ( .Y(D12199_Y), .B(D12200_Y), .A(D13257_Y));
KC_NAND2_X1 D12196 ( .Y(D12196_Y), .B(D13257_Y), .A(D10134_Y));
KC_NAND2_X1 D12195 ( .Y(D12195_Y), .B(D7782_Y), .A(D10134_Y));
KC_NAND2_X1 D12194 ( .Y(D12194_Y), .B(D4747_Y), .A(D6281_Y));
KC_NAND2_X1 D12190 ( .Y(D12190_Y), .B(D12212_Y), .A(D12198_Y));
KC_NAND2_X1 D12189 ( .Y(D12189_Y), .B(D13257_Y), .A(D12210_Y));
KC_NAND2_X1 D12027 ( .Y(D12027_Y), .B(D12028_Y), .A(D8222_Y));
KC_NAND2_X1 D12018 ( .Y(D12018_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D11957 ( .Y(D11957_Y), .B(D11421_Y), .A(D760_Y));
KC_NAND2_X1 D11956 ( .Y(D11956_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D11945 ( .Y(D11945_Y), .B(D11954_Y), .A(D8222_Y));
KC_NAND2_X1 D11942 ( .Y(D11942_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D11941 ( .Y(D11941_Y), .B(D11421_Y), .A(D760_Y));
KC_NAND2_X1 D11940 ( .Y(D11940_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D11645 ( .Y(D11645_Y), .B(D11651_Y), .A(D10181_Y));
KC_NAND2_X1 D11591 ( .Y(D11591_Y), .B(D2243_Y), .A(D1823_Y));
KC_NAND2_X1 D11554 ( .Y(D11554_Y), .B(D8472_Y), .A(D11546_Y));
KC_NAND2_X1 D11553 ( .Y(D11553_Y), .B(D2243_Y), .A(D1823_Y));
KC_NAND2_X1 D11552 ( .Y(D11552_Y), .B(D11551_Y), .A(D8473_Y));
KC_NAND2_X1 D11550 ( .Y(D11550_Y), .B(D11476_Y), .A(D2243_Y));
KC_NAND2_X1 D11549 ( .Y(D11549_Y), .B(D11546_Y), .A(D8472_Y));
KC_NAND2_X1 D11548 ( .Y(D11548_Y), .B(D11505_Y), .A(D2243_Y));
KC_NAND2_X1 D11547 ( .Y(D11547_Y), .B(D8473_Y), .A(D11551_Y));
KC_NAND2_X1 D11365 ( .Y(D11365_Y), .B(D11363_Y), .A(D8302_Y));
KC_NAND2_X1 D11358 ( .Y(D11358_Y), .B(D8302_Y), .A(D11363_Y));
KC_NAND2_X1 D11191 ( .Y(D11191_Y), .B(D11762_Y), .A(D10787_Y));
KC_NAND2_X1 D11152 ( .Y(D11152_Y), .B(D11322_Y), .A(D10861_Y));
KC_NAND2_X1 D11148 ( .Y(D11148_Y), .B(D11476_Y), .A(D11322_Y));
KC_NAND2_X1 D11144 ( .Y(D11144_Y), .B(D8258_Y), .A(D11145_Y));
KC_NAND2_X1 D11143 ( .Y(D11143_Y), .B(D11145_Y), .A(D8258_Y));
KC_NAND2_X1 D11090 ( .Y(D11090_Y), .B(D11098_Y), .A(D11112_Y));
KC_NAND2_X1 D10975 ( .Y(D10975_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D10972 ( .Y(D10972_Y), .B(D11421_Y), .A(D760_Y));
KC_NAND2_X1 D10971 ( .Y(D10971_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D10967 ( .Y(D10967_Y), .B(D8540_Y), .A(D8222_Y));
KC_NAND2_X1 D10966 ( .Y(D10966_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D10965 ( .Y(D10965_Y), .B(D8540_Y), .A(D8222_Y));
KC_NAND2_X1 D10963 ( .Y(D10963_Y), .B(D11421_Y), .A(D760_Y));
KC_NAND2_X1 D10855 ( .Y(D10855_Y), .B(D10854_Y), .A(D1961_Y));
KC_NAND2_X1 D10852 ( .Y(D10852_Y), .B(D11308_Y), .A(D10861_Y));
KC_NAND2_X1 D10847 ( .Y(D10847_Y), .B(D1961_Y), .A(D10854_Y));
KC_NAND2_X1 D10846 ( .Y(D10846_Y), .B(D11476_Y), .A(D11308_Y));
KC_NAND2_X1 D10734 ( .Y(D10734_Y), .B(D5403_Y), .A(D8222_Y));
KC_NAND2_X1 D10730 ( .Y(D10730_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D10729 ( .Y(D10729_Y), .B(D2206_Y), .A(D760_Y));
KC_NAND2_X1 D10728 ( .Y(D10728_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D10467 ( .Y(D10467_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D10465 ( .Y(D10465_Y), .B(D10994_Q), .A(D10505_Y));
KC_NAND2_X1 D10318 ( .Y(D10318_Y), .B(D10359_Q), .A(D10360_Q));
KC_NAND2_X1 D10258 ( .Y(D10258_Y), .B(D774_Y), .A(D848_Y));
KC_NAND2_X1 D10242 ( .Y(D10242_Y), .B(D2176_Y), .A(D9538_Y));
KC_NAND2_X1 D10136 ( .Y(D10136_Y), .B(D10137_Y), .A(D10629_Y));
KC_NAND2_X1 D10080 ( .Y(D10080_Y), .B(D9985_Y), .A(D9943_Y));
KC_NAND2_X1 D10075 ( .Y(D10075_Y), .B(D10076_Y), .A(D9218_Q));
KC_NAND2_X1 D10069 ( .Y(D10069_Y), .B(D10072_Y), .A(D10073_Y));
KC_NAND2_X1 D10068 ( .Y(D10068_Y), .B(D10071_Y), .A(D419_Q));
KC_NAND2_X1 D10037 ( .Y(D10037_Y), .B(D2166_Q), .A(D8900_Y));
KC_NAND2_X1 D10021 ( .Y(D10021_Y), .B(D10006_Q), .A(D2070_Y));
KC_NAND2_X1 D10017 ( .Y(D10017_Y), .B(D10031_Q), .A(D8900_Y));
KC_NAND2_X1 D10011 ( .Y(D10011_Y), .B(D10031_Q), .A(D7313_Y));
KC_NAND2_X1 D10002 ( .Y(D10002_Y), .B(D9983_Q), .A(D8900_Y));
KC_NAND2_X1 D9999 ( .Y(D9999_Y), .B(D10007_Q), .A(D2070_Y));
KC_NAND2_X1 D9995 ( .Y(D9995_Y), .B(D10008_Q), .A(D2070_Y));
KC_NAND2_X1 D9992 ( .Y(D9992_Y), .B(D10009_Q), .A(D8900_Y));
KC_NAND2_X1 D9527 ( .Y(D9527_Y), .B(D9528_Y), .A(D9575_Q));
KC_NAND2_X1 D9510 ( .Y(D9510_Y), .B(D9575_Q), .A(D9576_Q));
KC_NAND2_X1 D9509 ( .Y(D9509_Y), .B(D2039_Y), .A(D9575_Q));
KC_NAND2_X1 D9508 ( .Y(D9508_Y), .B(D2039_Y), .A(D9521_Y));
KC_NAND2_X1 D9502 ( .Y(D9502_Y), .B(D2039_Y), .A(D9528_Y));
KC_NAND2_X1 D9501 ( .Y(D9501_Y), .B(D9575_Q), .A(D9578_Q));
KC_NAND2_X1 D9498 ( .Y(D9498_Y), .B(D9502_Y), .A(D9539_Y));
KC_NAND2_X1 D9418 ( .Y(D9418_Y), .B(D625_Y), .A(D643_Y));
KC_NAND2_X1 D9417 ( .Y(D9417_Y), .B(D9439_Y), .A(D625_Y));
KC_NAND2_X1 D9412 ( .Y(D9412_Y), .B(D8083_Y), .A(D2063_Y));
KC_NAND2_X1 D9405 ( .Y(D9405_Y), .B(D8221_Y), .A(D9404_Y));
KC_NAND2_X1 D9398 ( .Y(D9398_Y), .B(D9441_Y), .A(D8221_Y));
KC_NAND2_X1 D9393 ( .Y(D9393_Y), .B(D8156_Y), .A(D9405_Y));
KC_NAND2_X1 D9392 ( .Y(D9392_Y), .B(D9421_Y), .A(D8079_Y));
KC_NAND2_X1 D9391 ( .Y(D9391_Y), .B(D9513_Y), .A(D1987_Y));
KC_NAND2_X1 D9369 ( .Y(D9369_Y), .B(D6288_Y), .A(D2312_Y));
KC_NAND2_X1 D9344 ( .Y(D9344_Y), .B(D9172_Y), .A(D4540_Y));
KC_NAND2_X1 D9299 ( .Y(D9299_Y), .B(D9247_Y), .A(D9246_Y));
KC_NAND2_X1 D9242 ( .Y(D9242_Y), .B(D7626_Y), .A(D9249_Y));
KC_NAND2_X1 D9240 ( .Y(D9240_Y), .B(D9147_Y), .A(D41_Y));
KC_NAND2_X1 D9192 ( .Y(D9192_Y), .B(D9213_Y), .A(D7683_Y));
KC_NAND2_X1 D9180 ( .Y(D9180_Y), .B(D9147_Y), .A(D8951_Q));
KC_NAND2_X1 D9175 ( .Y(D9175_Y), .B(D9147_Y), .A(D7481_Q));
KC_NAND2_X1 D9167 ( .Y(D9167_Y), .B(D9147_Y), .A(D57_Y));
KC_NAND2_X1 D9101 ( .Y(D9101_Y), .B(D9147_Y), .A(D8953_Q));
KC_NAND2_X1 D9164 ( .Y(D9164_Y), .B(D5966_Y), .A(D7470_Y));
KC_NAND2_X1 D9125 ( .Y(D9125_Y), .B(D9119_Y), .A(D9119_Y));
KC_NAND2_X1 D9121 ( .Y(D9121_Y), .B(D7635_Y), .A(D383_Y));
KC_NAND2_X1 D9113 ( .Y(D9113_Y), .B(D9147_Y), .A(D7501_Y));
KC_NAND2_X1 D9107 ( .Y(D9107_Y), .B(D9101_Y), .A(D9162_Y));
KC_NAND2_X1 D9027 ( .Y(D9027_Y), .B(D9029_Y), .A(D9028_Y));
KC_NAND2_X1 D8984 ( .Y(D8984_Y), .B(D8986_Y), .A(D2095_Y));
KC_NAND2_X1 D8970 ( .Y(D8970_Y), .B(D266_Y), .A(D5684_Y));
KC_NAND2_X1 D8964 ( .Y(D8964_Y), .B(D8986_Y), .A(D9481_Y));
KC_NAND2_X1 D8963 ( .Y(D8963_Y), .B(D8986_Y), .A(D9477_Y));
KC_NAND2_X1 D8919 ( .Y(D8919_Y), .B(D8937_Y), .A(D8904_Y));
KC_NAND2_X1 D8918 ( .Y(D8918_Y), .B(D283_Y), .A(D8950_Y));
KC_NAND2_X1 D8916 ( .Y(D8916_Y), .B(D7456_Y), .A(D9021_Q));
KC_NAND2_X1 D8913 ( .Y(D8913_Y), .B(D7456_Y), .A(D8951_Q));
KC_NAND2_X1 D8912 ( .Y(D8912_Y), .B(D7393_Y), .A(D2095_Y));
KC_NAND2_X1 D8910 ( .Y(D8910_Y), .B(D7393_Y), .A(D9477_Y));
KC_NAND2_X1 D8907 ( .Y(D8907_Y), .B(D7393_Y), .A(D9480_Y));
KC_NAND2_X1 D8871 ( .Y(D8871_Y), .B(D7393_Y), .A(D9475_Y));
KC_NAND2_X1 D8870 ( .Y(D8870_Y), .B(D7393_Y), .A(D9481_Y));
KC_NAND2_X1 D8864 ( .Y(D8864_Y), .B(D8859_Y), .A(D9012_Y));
KC_NAND2_X1 D8860 ( .Y(D8860_Y), .B(D8874_Y), .A(D9015_Y));
KC_NAND2_X1 D8853 ( .Y(D8853_Y), .B(D7393_Y), .A(D9476_Y));
KC_NAND2_X1 D8849 ( .Y(D8849_Y), .B(D7393_Y), .A(D9479_Y));
KC_NAND2_X1 D8848 ( .Y(D8848_Y), .B(D7393_Y), .A(D9482_Y));
KC_NAND2_X1 D8768 ( .Y(D8768_Y), .B(D8770_Y), .A(D8664_Y));
KC_NAND2_X1 D8766 ( .Y(D8766_Y), .B(D8767_Y), .A(D205_Y));
KC_NAND2_X1 D8764 ( .Y(D8764_Y), .B(D8762_Y), .A(D7110_Y));
KC_NAND2_X1 D8763 ( .Y(D8763_Y), .B(D8740_Y), .A(D8746_Y));
KC_NAND2_X1 D8758 ( .Y(D8758_Y), .B(D8772_Y), .A(D9480_Y));
KC_NAND2_X1 D8742 ( .Y(D8742_Y), .B(D2026_Y), .A(D9479_Y));
KC_NAND2_X1 D8740 ( .Y(D8740_Y), .B(D9981_Q), .A(D9980_Q));
KC_NAND2_X1 D8737 ( .Y(D8737_Y), .B(D8738_Y), .A(D8735_Y));
KC_NAND2_X1 D8736 ( .Y(D8736_Y), .B(D8737_Y), .A(D8738_Y));
KC_NAND2_X1 D8668 ( .Y(D8668_Y), .B(D9941_Q), .A(D8712_Q));
KC_NAND2_X1 D8500 ( .Y(D8500_Y), .B(D8534_Y), .A(D8466_Y));
KC_NAND2_X1 D8496 ( .Y(D8496_Y), .B(D5508_Y), .A(D8466_Y));
KC_NAND2_X1 D8419 ( .Y(D8419_Y), .B(D8463_Q), .A(D545_Y));
KC_NAND2_X1 D8413 ( .Y(D8413_Y), .B(D8368_Y), .A(D8382_Y));
KC_NAND2_X1 D8412 ( .Y(D8412_Y), .B(D8397_Y), .A(D8457_Y));
KC_NAND2_X1 D8403 ( .Y(D8403_Y), .B(D8414_Y), .A(D8405_Y));
KC_NAND2_X1 D8393 ( .Y(D8393_Y), .B(D8376_Y), .A(D7928_Y));
KC_NAND2_X1 D8392 ( .Y(D8392_Y), .B(D8460_Q), .A(D545_Y));
KC_NAND2_X1 D8386 ( .Y(D8386_Y), .B(D8405_Y), .A(D8387_Y));
KC_NAND2_X1 D8385 ( .Y(D8385_Y), .B(D8376_Y), .A(D8435_Y));
KC_NAND2_X1 D8378 ( .Y(D8378_Y), .B(D8410_Y), .A(D8279_Y));
KC_NAND2_X1 D8377 ( .Y(D8377_Y), .B(D6787_Y), .A(D8460_Q));
KC_NAND2_X1 D8370 ( .Y(D8370_Y), .B(D8418_Y), .A(D8279_Y));
KC_NAND2_X1 D8369 ( .Y(D8369_Y), .B(D11390_Q), .A(D545_Y));
KC_NAND2_X1 D8368 ( .Y(D8368_Y), .B(D11475_Q), .A(D545_Y));
KC_NAND2_X1 D8361 ( .Y(D8361_Y), .B(D8377_Y), .A(D8360_Y));
KC_NAND2_X1 D8360 ( .Y(D8360_Y), .B(D5496_Y), .A(D8466_Y));
KC_NAND2_X1 D8357 ( .Y(D8357_Y), .B(D8294_Y), .A(D6773_Y));
KC_NAND2_X1 D8293 ( .Y(D8293_Y), .B(D8245_Q), .A(D8244_Q));
KC_NAND2_X1 D8291 ( .Y(D8291_Y), .B(D8290_Y), .A(D8292_Y));
KC_NAND2_X1 D8289 ( .Y(D8289_Y), .B(D8292_Y), .A(D8048_Y));
KC_NAND2_X1 D8288 ( .Y(D8288_Y), .B(D16755_Y), .A(D8047_Y));
KC_NAND2_X1 D8281 ( .Y(D8281_Y), .B(D942_Y), .A(D957_Y));
KC_NAND2_X1 D8280 ( .Y(D8280_Y), .B(D8415_Y), .A(D8286_Y));
KC_NAND2_X1 D8262 ( .Y(D8262_Y), .B(D8219_Y), .A(D8239_Y));
KC_NAND2_X1 D8204 ( .Y(D8204_Y), .B(D8248_Q), .A(D8202_Y));
KC_NAND2_X1 D8199 ( .Y(D8199_Y), .B(D8459_Q), .A(D7916_Y));
KC_NAND2_X1 D8198 ( .Y(D8198_Y), .B(D8210_Y), .A(D5288_Y));
KC_NAND2_X1 D8190 ( .Y(D8190_Y), .B(D8220_Y), .A(D9559_Y));
KC_NAND2_X1 D8185 ( .Y(D8185_Y), .B(D7669_Y), .A(D7668_Y));
KC_NAND2_X1 D8182 ( .Y(D8182_Y), .B(D8240_Y), .A(D6709_Y));
KC_NAND2_X1 D8181 ( .Y(D8181_Y), .B(D8240_Y), .A(D3776_Y));
KC_NAND2_X1 D8115 ( .Y(D8115_Y), .B(D7782_Y), .A(D6014_Y));
KC_NAND2_X1 D8109 ( .Y(D8109_Y), .B(D8106_Y), .A(D8120_Y));
KC_NAND2_X1 D8094 ( .Y(D8094_Y), .B(D8220_Y), .A(D1984_Y));
KC_NAND2_X1 D8093 ( .Y(D8093_Y), .B(D9444_Y), .A(D8125_Y));
KC_NAND2_X1 D8092 ( .Y(D8092_Y), .B(D7475_Q), .A(D8098_Y));
KC_NAND2_X1 D8091 ( .Y(D8091_Y), .B(D8128_Y), .A(D8090_Y));
KC_NAND2_X1 D8081 ( .Y(D8081_Y), .B(D5213_Y), .A(D8240_Y));
KC_NAND2_X1 D8018 ( .Y(D8018_Y), .B(D1849_Y), .A(D8015_Y));
KC_NAND2_X1 D8017 ( .Y(D8017_Y), .B(D7670_Y), .A(D8001_Y));
KC_NAND2_X1 D7985 ( .Y(D7985_Y), .B(D7963_Y), .A(D7947_Y));
KC_NAND2_X1 D7946 ( .Y(D7946_Y), .B(D7948_Y), .A(D531_Q));
KC_NAND2_X1 D7938 ( .Y(D7938_Y), .B(D7942_Y), .A(D531_Q));
KC_NAND2_X1 D7937 ( .Y(D7937_Y), .B(D7941_Y), .A(D7942_Y));
KC_NAND2_X1 D7925 ( .Y(D7925_Y), .B(D532_Q), .A(D533_Q));
KC_NAND2_X1 D7924 ( .Y(D7924_Y), .B(D7917_Y), .A(D533_Q));
KC_NAND2_X1 D7923 ( .Y(D7923_Y), .B(D7917_Y), .A(D7926_Y));
KC_NAND2_X1 D7922 ( .Y(D7922_Y), .B(D7926_Y), .A(D532_Q));
KC_NAND2_X1 D7918 ( .Y(D7918_Y), .B(D7913_Y), .A(D9375_Y));
KC_NAND2_X1 D7853 ( .Y(D7853_Y), .B(D7874_Y), .A(D7902_Y));
KC_NAND2_X1 D7852 ( .Y(D7852_Y), .B(D6441_Y), .A(D7858_Y));
KC_NAND2_X1 D7848 ( .Y(D7848_Y), .B(D7842_Y), .A(D7866_Y));
KC_NAND2_X1 D7847 ( .Y(D7847_Y), .B(D7867_Y), .A(D7875_Y));
KC_NAND2_X1 D7842 ( .Y(D7842_Y), .B(D6787_Y), .A(D7953_Y));
KC_NAND2_X1 D7838 ( .Y(D7838_Y), .B(D7827_Y), .A(D7888_Q));
KC_NAND2_X1 D7837 ( .Y(D7837_Y), .B(D7834_Y), .A(D1860_Y));
KC_NAND2_X1 D7832 ( .Y(D7832_Y), .B(D7839_Y), .A(D7833_Y));
KC_NAND2_X1 D7831 ( .Y(D7831_Y), .B(D7835_Y), .A(D7927_Y));
KC_NAND2_X1 D7830 ( .Y(D7830_Y), .B(D7862_Y), .A(D7831_Y));
KC_NAND2_X1 D7829 ( .Y(D7829_Y), .B(D7835_Y), .A(D533_Q));
KC_NAND2_X1 D7762 ( .Y(D7762_Y), .B(D7775_Y), .A(D9254_Y));
KC_NAND2_X1 D7753 ( .Y(D7753_Y), .B(D9210_Y), .A(D7706_Y));
KC_NAND2_X1 D7683 ( .Y(D7683_Y), .B(D9147_Y), .A(D9021_Q));
KC_NAND2_X1 D7620 ( .Y(D7620_Y), .B(D6075_Y), .A(D7671_Y));
KC_NAND2_X1 D7565 ( .Y(D7565_Y), .B(D7587_Q), .A(D7586_Q));
KC_NAND2_X1 D7564 ( .Y(D7564_Y), .B(D102_Y), .A(D4150_Y));
KC_NAND2_X1 D7563 ( .Y(D7563_Y), .B(D1787_Y), .A(D102_Y));
KC_NAND2_X1 D7510 ( .Y(D7510_Y), .B(D7418_Y), .A(D5684_Y));
KC_NAND2_X1 D7508 ( .Y(D7508_Y), .B(D9147_Y), .A(D7479_Q));
KC_NAND2_X1 D7504 ( .Y(D7504_Y), .B(D1871_Y), .A(D11642_Y));
KC_NAND2_X1 D7503 ( .Y(D7503_Y), .B(D7501_Y), .A(D7499_Y));
KC_NAND2_X1 D7500 ( .Y(D7500_Y), .B(D7501_Y), .A(D5969_Y));
KC_NAND2_X1 D7491 ( .Y(D7491_Y), .B(D36_Y), .A(D9041_Y));
KC_NAND2_X1 D7445 ( .Y(D7445_Y), .B(D7456_Y), .A(D7481_Q));
KC_NAND2_X1 D7444 ( .Y(D7444_Y), .B(D7315_Y), .A(D273_Y));
KC_NAND2_X1 D7427 ( .Y(D7427_Y), .B(D7426_Y), .A(D9473_Y));
KC_NAND2_X1 D7414 ( .Y(D7414_Y), .B(D24_Y), .A(D7413_Y));
KC_NAND2_X1 D7413 ( .Y(D7413_Y), .B(D9147_Y), .A(D36_Y));
KC_NAND2_X1 D7359 ( .Y(D7359_Y), .B(D257_Y), .A(D7153_Y));
KC_NAND2_X1 D7358 ( .Y(D7358_Y), .B(D2892_Y), .A(D257_Y));
KC_NAND2_X1 D7352 ( .Y(D7352_Y), .B(D7143_Y), .A(D5804_Y));
KC_NAND2_X1 D7343 ( .Y(D7343_Y), .B(D7323_Y), .A(D5656_Y));
KC_NAND2_X1 D7316 ( .Y(D7316_Y), .B(D5677_Y), .A(D12176_Y));
KC_NAND2_X1 D7303 ( .Y(D7303_Y), .B(D7110_Y), .A(D7109_Y));
KC_NAND2_X1 D7259 ( .Y(D7259_Y), .B(D5804_Y), .A(D7195_Y));
KC_NAND2_X1 D7258 ( .Y(D7258_Y), .B(D6333_Y), .A(D7141_Y));
KC_NAND2_X1 D7246 ( .Y(D7246_Y), .B(D6470_Y), .A(D7140_Y));
KC_NAND2_X1 D7245 ( .Y(D7245_Y), .B(D7236_Y), .A(D7248_Y));
KC_NAND2_X1 D7238 ( .Y(D7238_Y), .B(D7188_Y), .A(D8760_Y));
KC_NAND2_X1 D7237 ( .Y(D7237_Y), .B(D8778_Y), .A(D7239_Y));
KC_NAND2_X1 D7236 ( .Y(D7236_Y), .B(D8778_Y), .A(D8741_Y));
KC_NAND2_X1 D7229 ( .Y(D7229_Y), .B(D1887_Y), .A(D7217_Y));
KC_NAND2_X1 D7224 ( .Y(D7224_Y), .B(D8754_Y), .A(D7228_Y));
KC_NAND2_X1 D7216 ( .Y(D7216_Y), .B(D8778_Y), .A(D2026_Y));
KC_NAND2_X1 D7211 ( .Y(D7211_Y), .B(D7219_Y), .A(D5768_Y));
KC_NAND2_X1 D7206 ( .Y(D7206_Y), .B(D8749_Y), .A(D8876_Y));
KC_NAND2_X1 D7198 ( .Y(D7198_Y), .B(D1970_Y), .A(D7182_Y));
KC_NAND2_X1 D7197 ( .Y(D7197_Y), .B(D4444_Y), .A(D247_Y));
KC_NAND2_X1 D7187 ( .Y(D7187_Y), .B(D8752_Y), .A(D7238_Y));
KC_NAND2_X1 D7181 ( .Y(D7181_Y), .B(D202_Y), .A(D7175_Y));
KC_NAND2_X1 D7180 ( .Y(D7180_Y), .B(D209_Y), .A(D7186_Y));
KC_NAND2_X1 D7179 ( .Y(D7179_Y), .B(D7175_Y), .A(D7171_Y));
KC_NAND2_X1 D7178 ( .Y(D7178_Y), .B(D8756_Y), .A(D7209_Y));
KC_NAND2_X1 D7176 ( .Y(D7176_Y), .B(D7239_Y), .A(D8812_Y));
KC_NAND2_X1 D7175 ( .Y(D7175_Y), .B(D7188_Y), .A(D7239_Y));
KC_NAND2_X1 D7169 ( .Y(D7169_Y), .B(D7214_Y), .A(D8754_Y));
KC_NAND2_X1 D7115 ( .Y(D7115_Y), .B(D7144_Q), .A(D7146_Q));
KC_NAND2_X1 D7111 ( .Y(D7111_Y), .B(D7124_Y), .A(D5880_Y));
KC_NAND2_X1 D7105 ( .Y(D7105_Y), .B(D5804_Y), .A(D7108_Y));
KC_NAND2_X1 D7104 ( .Y(D7104_Y), .B(D189_Y), .A(D7137_Y));
KC_NAND2_X1 D7097 ( .Y(D7097_Y), .B(D7106_Y), .A(D7099_Y));
KC_NAND2_X1 D7096 ( .Y(D7096_Y), .B(D5864_Y), .A(D7098_Y));
KC_NAND2_X1 D7095 ( .Y(D7095_Y), .B(D7098_Y), .A(D6334_Y));
KC_NAND2_X1 D6938 ( .Y(D6938_Y), .B(D7830_Y), .A(D6877_Y));
KC_NAND2_X1 D6935 ( .Y(D6935_Y), .B(D8540_Y), .A(D8222_Y));
KC_NAND2_X1 D6934 ( .Y(D6934_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D6928 ( .Y(D6928_Y), .B(D8466_Y), .A(D5501_Y));
KC_NAND2_X1 D6854 ( .Y(D6854_Y), .B(D8540_Y), .A(D8222_Y));
KC_NAND2_X1 D6842 ( .Y(D6842_Y), .B(D8371_Y), .A(D968_Y));
KC_NAND2_X1 D6782 ( .Y(D6782_Y), .B(D5403_Y), .A(D8222_Y));
KC_NAND2_X1 D6780 ( .Y(D6780_Y), .B(D6800_Y), .A(D5214_Y));
KC_NAND2_X1 D6719 ( .Y(D6719_Y), .B(D6618_Y), .A(D8240_Y));
KC_NAND2_X1 D6516 ( .Y(D6516_Y), .B(D6566_Y), .A(D6517_Y));
KC_NAND2_X1 D6447 ( .Y(D6447_Y), .B(D1793_Q), .A(D6259_Y));
KC_NAND2_X1 D6443 ( .Y(D6443_Y), .B(D3408_Y), .A(D6449_Y));
KC_NAND2_X1 D6437 ( .Y(D6437_Y), .B(D6463_Y), .A(D6426_Y));
KC_NAND2_X1 D6433 ( .Y(D6433_Y), .B(D6432_Y), .A(D6486_Q));
KC_NAND2_X1 D6430 ( .Y(D6430_Y), .B(D5031_Y), .A(D4866_Y));
KC_NAND2_X1 D6363 ( .Y(D6363_Y), .B(D6375_Q), .A(D6376_Q));
KC_NAND2_X1 D6362 ( .Y(D6362_Y), .B(D1698_Y), .A(D444_Q));
KC_NAND2_X1 D14139 ( .Y(D14139_Y), .B(D6238_Y), .A(D6254_Y));
KC_NAND2_X1 D12130 ( .Y(D12130_Y), .B(D6240_Y), .A(D6212_Y));
KC_NAND2_X1 D6234 ( .Y(D6234_Y), .B(D6245_Y), .A(D6252_Y));
KC_NAND2_X1 D6227 ( .Y(D6227_Y), .B(D6228_Y), .A(D6244_Y));
KC_NAND2_X1 D9105 ( .Y(D9105_Y), .B(D6183_Y), .A(D6157_Y));
KC_NAND2_X1 D6145 ( .Y(D6145_Y), .B(D6253_Y), .A(D6144_Y));
KC_NAND2_X1 D6368 ( .Y(D6368_Y), .B(D6105_Y), .A(D16143_Y));
KC_NAND2_X1 D6097 ( .Y(D6097_Y), .B(D1787_Y), .A(D20_Y));
KC_NAND2_X1 D6096 ( .Y(D6096_Y), .B(D1713_Y), .A(D20_Y));
KC_NAND2_X1 D6036 ( .Y(D6036_Y), .B(D4493_Y), .A(D1719_Y));
KC_NAND2_X1 D6035 ( .Y(D6035_Y), .B(D6013_Y), .A(D5698_Y));
KC_NAND2_X1 D6034 ( .Y(D6034_Y), .B(D6054_Y), .A(D5871_Y));
KC_NAND2_X1 D6021 ( .Y(D6021_Y), .B(D4402_Y), .A(D7242_Y));
KC_NAND2_X1 D6011 ( .Y(D6011_Y), .B(D6000_Y), .A(D5755_Y));
KC_NAND2_X1 D6010 ( .Y(D6010_Y), .B(D5984_Y), .A(D5755_Y));
KC_NAND2_X1 D6009 ( .Y(D6009_Y), .B(D6013_Y), .A(D5646_Y));
KC_NAND2_X1 D5985 ( .Y(D5985_Y), .B(D6046_Y), .A(D6033_Y));
KC_NAND2_X1 D5978 ( .Y(D5978_Y), .B(D6024_Y), .A(D5641_Y));
KC_NAND2_X1 D5975 ( .Y(D5975_Y), .B(D4416_Y), .A(D277_Y));
KC_NAND2_X1 D5974 ( .Y(D5974_Y), .B(D277_Y), .A(D239_Q));
KC_NAND2_X1 D5973 ( .Y(D5973_Y), .B(D4150_Y), .A(D235_Y));
KC_NAND2_X1 D5972 ( .Y(D5972_Y), .B(D6024_Y), .A(D6001_Y));
KC_NAND2_X1 D5963 ( .Y(D5963_Y), .B(D6075_Y), .A(D5970_Y));
KC_NAND2_X1 D5957 ( .Y(D5957_Y), .B(D1712_Y), .A(D6033_Y));
KC_NAND2_X1 D5956 ( .Y(D5956_Y), .B(D165_Y), .A(D4149_Q));
KC_NAND2_X1 D5955 ( .Y(D5955_Y), .B(D4149_Q), .A(D8313_Q));
KC_NAND2_X1 D5888 ( .Y(D5888_Y), .B(D7984_Y), .A(D5698_Y));
KC_NAND2_X1 D5887 ( .Y(D5887_Y), .B(D6024_Y), .A(D6034_Y));
KC_NAND2_X1 D5886 ( .Y(D5886_Y), .B(D5852_Y), .A(D5968_Y));
KC_NAND2_X1 D5885 ( .Y(D5885_Y), .B(D4350_Y), .A(D5684_Y));
KC_NAND2_X1 D5884 ( .Y(D5884_Y), .B(D266_Y), .A(D6039_Y));
KC_NAND2_X1 D5876 ( .Y(D5876_Y), .B(D7242_Y), .A(D5889_Y));
KC_NAND2_X1 D5875 ( .Y(D5875_Y), .B(D7372_Y), .A(D5945_Y));
KC_NAND2_X1 D5874 ( .Y(D5874_Y), .B(D7984_Y), .A(D5871_Y));
KC_NAND2_X1 D5865 ( .Y(D5865_Y), .B(D7371_Y), .A(D5945_Y));
KC_NAND2_X1 D5864 ( .Y(D5864_Y), .B(D5890_Y), .A(D7242_Y));
KC_NAND2_X1 D5857 ( .Y(D5857_Y), .B(D4340_Y), .A(D7242_Y));
KC_NAND2_X1 D5849 ( .Y(D5849_Y), .B(D4282_Y), .A(D7100_Y));
KC_NAND2_X1 D5848 ( .Y(D5848_Y), .B(D5997_Y), .A(D4425_Y));
KC_NAND2_X1 D5847 ( .Y(D5847_Y), .B(D4233_Y), .A(D5851_Y));
KC_NAND2_X1 D5846 ( .Y(D5846_Y), .B(D5877_Y), .A(D262_Y));
KC_NAND2_X1 D5840 ( .Y(D5840_Y), .B(D6001_Y), .A(D5866_Y));
KC_NAND2_X1 D5834 ( .Y(D5834_Y), .B(D4233_Y), .A(D5646_Y));
KC_NAND2_X1 D5829 ( .Y(D5829_Y), .B(D5763_Y), .A(D6032_Y));
KC_NAND2_X1 D5828 ( .Y(D5828_Y), .B(D7329_Y), .A(D5763_Y));
KC_NAND2_X1 D5771 ( .Y(D5771_Y), .B(D7092_Y), .A(D186_Y));
KC_NAND2_X1 D5769 ( .Y(D5769_Y), .B(D5804_Y), .A(D7234_Y));
KC_NAND2_X1 D5762 ( .Y(D5762_Y), .B(D1734_Y), .A(D5715_Y));
KC_NAND2_X1 D5761 ( .Y(D5761_Y), .B(D1617_Y), .A(D5737_Y));
KC_NAND2_X1 D5753 ( .Y(D5753_Y), .B(D1739_Y), .A(D5742_Y));
KC_NAND2_X1 D5747 ( .Y(D5747_Y), .B(D6039_Y), .A(D5755_Y));
KC_NAND2_X1 D5746 ( .Y(D5746_Y), .B(D5980_Y), .A(D5841_Y));
KC_NAND2_X1 D5745 ( .Y(D5745_Y), .B(D5722_Y), .A(D4305_Y));
KC_NAND2_X1 D5744 ( .Y(D5744_Y), .B(D7500_Y), .A(D5644_Y));
KC_NAND2_X1 D5743 ( .Y(D5743_Y), .B(D6056_Y), .A(D5671_Y));
KC_NAND2_X1 D5728 ( .Y(D5728_Y), .B(D5744_Y), .A(D1726_Y));
KC_NAND2_X1 D5727 ( .Y(D5727_Y), .B(D7193_Y), .A(D9477_Y));
KC_NAND2_X1 D5721 ( .Y(D5721_Y), .B(D5768_Y), .A(D203_Y));
KC_NAND2_X1 D5713 ( .Y(D5713_Y), .B(D7292_Y), .A(D203_Y));
KC_NAND2_X1 D5712 ( .Y(D5712_Y), .B(D4226_Y), .A(D4119_Q));
KC_NAND2_X1 D5668 ( .Y(D5668_Y), .B(D5669_Y), .A(D5689_Q));
KC_NAND2_X1 D5663 ( .Y(D5663_Y), .B(D5664_Y), .A(D5660_Y));
KC_NAND2_X1 D5662 ( .Y(D5662_Y), .B(D5660_Y), .A(D5691_Q));
KC_NAND2_X1 D5661 ( .Y(D5661_Y), .B(D5664_Y), .A(D5690_Q));
KC_NAND2_X1 D5658 ( .Y(D5658_Y), .B(D5670_Y), .A(D5804_Y));
KC_NAND2_X1 D5654 ( .Y(D5654_Y), .B(D5667_Y), .A(D5688_Q));
KC_NAND2_X1 D5651 ( .Y(D5651_Y), .B(D186_Y), .A(D7093_Y));
KC_NAND2_X1 D5647 ( .Y(D5647_Y), .B(D5652_Y), .A(D5653_Y));
KC_NAND2_X1 D5520 ( .Y(D5520_Y), .B(D5432_Y), .A(D760_Y));
KC_NAND2_X1 D5518 ( .Y(D5518_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D5442 ( .Y(D5442_Y), .B(D5432_Y), .A(D760_Y));
KC_NAND2_X1 D5431 ( .Y(D5431_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D5368 ( .Y(D5368_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D5359 ( .Y(D5359_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D5358 ( .Y(D5358_Y), .B(D5403_Y), .A(D8222_Y));
KC_NAND2_X1 D5357 ( .Y(D5357_Y), .B(D5432_Y), .A(D760_Y));
KC_NAND2_X1 D5350 ( .Y(D5350_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D5267 ( .Y(D5267_Y), .B(D5432_Y), .A(D760_Y));
KC_NAND2_X1 D5097 ( .Y(D5097_Y), .B(D3633_Y), .A(D5064_Y));
KC_NAND2_X1 D5042 ( .Y(D5042_Y), .B(D3371_Y), .A(D1565_Y));
KC_NAND2_X1 D5041 ( .Y(D5041_Y), .B(D3498_Y), .A(D1537_Y));
KC_NAND2_X1 D5040 ( .Y(D5040_Y), .B(D5011_Y), .A(D4880_Y));
KC_NAND2_X1 D5031 ( .Y(D5031_Y), .B(D5012_Y), .A(D4900_Y));
KC_NAND2_X1 D5030 ( .Y(D5030_Y), .B(D5033_Y), .A(D4985_Y));
KC_NAND2_X1 D5021 ( .Y(D5021_Y), .B(D3371_Y), .A(D4886_Y));
KC_NAND2_X1 D5020 ( .Y(D5020_Y), .B(D3371_Y), .A(D3499_Y));
KC_NAND2_X1 D5019 ( .Y(D5019_Y), .B(D4886_Y), .A(D3498_Y));
KC_NAND2_X1 D5018 ( .Y(D5018_Y), .B(D4868_Y), .A(D3484_Q));
KC_NAND2_X1 D5005 ( .Y(D5005_Y), .B(D5012_Y), .A(D3599_Y));
KC_NAND2_X1 D5001 ( .Y(D5001_Y), .B(D3594_Y), .A(D3509_Y));
KC_NAND2_X1 D5000 ( .Y(D5000_Y), .B(D4996_Y), .A(D4883_Y));
KC_NAND2_X1 D4999 ( .Y(D4999_Y), .B(D5009_Y), .A(D3599_Y));
KC_NAND2_X1 D4998 ( .Y(D4998_Y), .B(D1565_Y), .A(D4985_Y));
KC_NAND2_X1 D4992 ( .Y(D4992_Y), .B(D3509_Y), .A(D3446_Y));
KC_NAND2_X1 D4991 ( .Y(D4991_Y), .B(D5038_Y), .A(D4877_Y));
KC_NAND2_X1 D4983 ( .Y(D4983_Y), .B(D5033_Y), .A(D4877_Y));
KC_NAND2_X1 D4982 ( .Y(D4982_Y), .B(D5079_Y), .A(D5082_Y));
KC_NAND2_X1 D4923 ( .Y(D4923_Y), .B(D3371_Y), .A(D3400_Y));
KC_NAND2_X1 D4922 ( .Y(D4922_Y), .B(D4926_Y), .A(D3388_Q));
KC_NAND2_X1 D4921 ( .Y(D4921_Y), .B(D448_Y), .A(D4962_Y));
KC_NAND2_X1 D4916 ( .Y(D4916_Y), .B(D1570_Y), .A(D1537_Y));
KC_NAND2_X1 D4915 ( .Y(D4915_Y), .B(D3416_Y), .A(D1537_Y));
KC_NAND2_X1 D4914 ( .Y(D4914_Y), .B(D4926_Y), .A(D3400_Y));
KC_NAND2_X1 D4909 ( .Y(D4909_Y), .B(D4920_Y), .A(D4900_Y));
KC_NAND2_X1 D4902 ( .Y(D4902_Y), .B(D3416_Y), .A(D4897_Y));
KC_NAND2_X1 D4901 ( .Y(D4901_Y), .B(D3501_Y), .A(D4903_Y));
KC_NAND2_X1 D4896 ( .Y(D4896_Y), .B(D3421_Y), .A(D3499_Y));
KC_NAND2_X1 D4895 ( .Y(D4895_Y), .B(D4920_Y), .A(D3499_Y));
KC_NAND2_X1 D4894 ( .Y(D4894_Y), .B(D4906_Y), .A(D1537_Y));
KC_NAND2_X1 D4893 ( .Y(D4893_Y), .B(D4900_Y), .A(D3499_Y));
KC_NAND2_X1 D4888 ( .Y(D4888_Y), .B(D4868_Y), .A(D3499_Y));
KC_NAND2_X1 D4881 ( .Y(D4881_Y), .B(D4874_Y), .A(D1537_Y));
KC_NAND2_X1 D4880 ( .Y(D4880_Y), .B(D3509_Y), .A(D4874_Y));
KC_NAND2_X1 D4879 ( .Y(D4879_Y), .B(D3371_Y), .A(D4891_Y));
KC_NAND2_X1 D4865 ( .Y(D4865_Y), .B(D4883_Y), .A(D3365_Y));
KC_NAND2_X1 D4858 ( .Y(D4858_Y), .B(D4856_Y), .A(D4824_Q));
KC_NAND2_X1 D4855 ( .Y(D4855_Y), .B(D4852_Y), .A(D4823_Q));
KC_NAND2_X1 D4854 ( .Y(D4854_Y), .B(D4848_Y), .A(D4825_Q));
KC_NAND2_X1 D4851 ( .Y(D4851_Y), .B(D4849_Y), .A(D1655_Q));
KC_NAND2_X1 D4850 ( .Y(D4850_Y), .B(D4853_Y), .A(D4817_Q));
KC_NAND2_X1 D4847 ( .Y(D4847_Y), .B(D3993_Y), .A(D4826_Q));
KC_NAND2_X1 D4843 ( .Y(D4843_Y), .B(D4779_Y), .A(D4700_Y));
KC_NAND2_X1 D4772 ( .Y(D4772_Y), .B(D4771_Y), .A(D1456_Y));
KC_NAND2_X1 D4770 ( .Y(D4770_Y), .B(D9345_Y), .A(D4576_Y));
KC_NAND2_X1 D4758 ( .Y(D4758_Y), .B(D4812_Y), .A(D4812_Y));
KC_NAND2_X1 D4748 ( .Y(D4748_Y), .B(D402_Y), .A(D4920_Y));
KC_NAND2_X1 D4696 ( .Y(D4696_Y), .B(D1573_Y), .A(D4709_Y));
KC_NAND2_X1 D4695 ( .Y(D4695_Y), .B(D4659_Y), .A(D3126_Y));
KC_NAND2_X1 D4693 ( .Y(D4693_Y), .B(D4575_Y), .A(D4688_Y));
KC_NAND2_X1 D4692 ( .Y(D4692_Y), .B(D372_Y), .A(D3255_Y));
KC_NAND2_X1 D4690 ( .Y(D4690_Y), .B(D1606_Y), .A(D4737_Y));
KC_NAND2_X1 D4684 ( .Y(D4684_Y), .B(D372_Y), .A(D4666_Y));
KC_NAND2_X1 D4673 ( .Y(D4673_Y), .B(D4675_Y), .A(D4524_Y));
KC_NAND2_X1 D4672 ( .Y(D4672_Y), .B(D4668_Y), .A(D4727_Q));
KC_NAND2_X1 D4671 ( .Y(D4671_Y), .B(D4666_Y), .A(D4668_Y));
KC_NAND2_X1 D4663 ( .Y(D4663_Y), .B(D4660_Y), .A(D3214_Y));
KC_NAND2_X1 D4658 ( .Y(D4658_Y), .B(D12653_Y), .A(D3258_Y));
KC_NAND2_X1 D4605 ( .Y(D4605_Y), .B(D4601_Y), .A(D4503_Y));
KC_NAND2_X1 D4601 ( .Y(D4601_Y), .B(D4640_Q), .A(D4591_Y));
KC_NAND2_X1 D4586 ( .Y(D4586_Y), .B(D4636_Q), .A(D4640_Q));
KC_NAND2_X1 D4585 ( .Y(D4585_Y), .B(D4581_Y), .A(D4595_Y));
KC_NAND2_X1 D4580 ( .Y(D4580_Y), .B(D4595_Y), .A(D4638_Q));
KC_NAND2_X1 D4579 ( .Y(D4579_Y), .B(D4589_Y), .A(D4636_Q));
KC_NAND2_X1 D4509 ( .Y(D4509_Y), .B(D3016_Y), .A(D3041_Y));
KC_NAND2_X1 D4504 ( .Y(D4504_Y), .B(D4501_Y), .A(D312_Y));
KC_NAND2_X1 D4499 ( .Y(D4499_Y), .B(D3012_Y), .A(D3018_Y));
KC_NAND2_X1 D4498 ( .Y(D4498_Y), .B(D4505_Y), .A(D1578_Y));
KC_NAND2_X1 D4448 ( .Y(D4448_Y), .B(D4434_Y), .A(D4116_Y));
KC_NAND2_X1 D4447 ( .Y(D4447_Y), .B(D2878_Y), .A(D4116_Y));
KC_NAND2_X1 D4446 ( .Y(D4446_Y), .B(D6033_Y), .A(D5988_Y));
KC_NAND2_X1 D4426 ( .Y(D4426_Y), .B(D4489_Q), .A(D5772_Y));
KC_NAND2_X1 D4425 ( .Y(D4425_Y), .B(D4427_Y), .A(D1787_Y));
KC_NAND2_X1 D4420 ( .Y(D4420_Y), .B(D4418_Y), .A(D4149_Q));
KC_NAND2_X1 D4419 ( .Y(D4419_Y), .B(D4438_Y), .A(D239_Q));
KC_NAND2_X1 D4415 ( .Y(D4415_Y), .B(D4294_Y), .A(D228_Q));
KC_NAND2_X1 D4413 ( .Y(D4413_Y), .B(D4235_Q), .A(D228_Q));
KC_NAND2_X1 D4410 ( .Y(D4410_Y), .B(D4412_Y), .A(D4235_Q));
KC_NAND2_X1 D4409 ( .Y(D4409_Y), .B(D4294_Y), .A(D4412_Y));
KC_NAND2_X1 D4360 ( .Y(D4360_Y), .B(D4306_Y), .A(D4345_Y));
KC_NAND2_X1 D4359 ( .Y(D4359_Y), .B(D7503_Y), .A(D4292_Y));
KC_NAND2_X1 D4358 ( .Y(D4358_Y), .B(D4348_Y), .A(D4345_Y));
KC_NAND2_X1 D4349 ( .Y(D4349_Y), .B(D4301_Y), .A(D5889_Y));
KC_NAND2_X1 D4348 ( .Y(D4348_Y), .B(D4306_Y), .A(D4291_Y));
KC_NAND2_X1 D4347 ( .Y(D4347_Y), .B(D4430_Y), .A(D5872_Y));
KC_NAND2_X1 D4337 ( .Y(D4337_Y), .B(D7394_Y), .A(D7295_Y));
KC_NAND2_X1 D4326 ( .Y(D4326_Y), .B(D4322_Y), .A(D4277_Y));
KC_NAND2_X1 D4325 ( .Y(D4325_Y), .B(D7737_Q), .A(D4368_Y));
KC_NAND2_X1 D4324 ( .Y(D4324_Y), .B(D7730_Y), .A(D4390_Y));
KC_NAND2_X1 D4323 ( .Y(D4323_Y), .B(D5890_Y), .A(D4320_Y));
KC_NAND2_X1 D4317 ( .Y(D4317_Y), .B(D4315_Y), .A(D4277_Y));
KC_NAND2_X1 D4316 ( .Y(D4316_Y), .B(D4319_Y), .A(D4318_Y));
KC_NAND2_X1 D4315 ( .Y(D4315_Y), .B(D4318_Y), .A(D262_Y));
KC_NAND2_X1 D4309 ( .Y(D4309_Y), .B(D5855_Y), .A(D4233_Y));
KC_NAND2_X1 D4303 ( .Y(D4303_Y), .B(D4327_Y), .A(D5863_Y));
KC_NAND2_X1 D4302 ( .Y(D4302_Y), .B(D4283_Y), .A(D4296_Y));
KC_NAND2_X1 D4292 ( .Y(D4292_Y), .B(D4456_Y), .A(D165_Y));
KC_NAND2_X1 D4283 ( .Y(D4283_Y), .B(D4441_Y), .A(D4276_Y));
KC_NAND2_X1 D4282 ( .Y(D4282_Y), .B(D3038_Y), .A(D4276_Y));
KC_NAND2_X1 D4281 ( .Y(D4281_Y), .B(D4303_Y), .A(D4293_Y));
KC_NAND2_X1 D4280 ( .Y(D4280_Y), .B(D5833_Y), .A(D1629_Y));
KC_NAND2_X1 D4279 ( .Y(D4279_Y), .B(D4282_Y), .A(D4287_Y));
KC_NAND2_X1 D4268 ( .Y(D4268_Y), .B(D4266_Y), .A(D8838_Y));
KC_NAND2_X1 D4265 ( .Y(D4265_Y), .B(D235_Y), .A(D4150_Y));
KC_NAND2_X1 D4260 ( .Y(D4260_Y), .B(D2810_Y), .A(D228_Q));
KC_NAND2_X1 D4259 ( .Y(D4259_Y), .B(D4253_Y), .A(D229_Q));
KC_NAND2_X1 D4255 ( .Y(D4255_Y), .B(D4261_Y), .A(D165_Y));
KC_NAND2_X1 D4254 ( .Y(D4254_Y), .B(D5693_Q), .A(D4136_Q));
KC_NAND2_X1 D4251 ( .Y(D4251_Y), .B(D4258_Y), .A(D232_Q));
KC_NAND2_X1 D4202 ( .Y(D4202_Y), .B(D4370_Y), .A(D5863_Y));
KC_NAND2_X1 D4201 ( .Y(D4201_Y), .B(D4166_Y), .A(D4191_Y));
KC_NAND2_X1 D4197 ( .Y(D4197_Y), .B(D4168_Y), .A(D4187_Y));
KC_NAND2_X1 D4166 ( .Y(D4166_Y), .B(D4356_Y), .A(D5863_Y));
KC_NAND2_X1 D4165 ( .Y(D4165_Y), .B(D241_Y), .A(D4164_Y));
KC_NAND2_X1 D4152 ( .Y(D4152_Y), .B(D4256_Y), .A(D4149_Q));
KC_NAND2_X1 D4147 ( .Y(D4147_Y), .B(D4252_Y), .A(D4121_Q));
KC_NAND2_X1 D4143 ( .Y(D4143_Y), .B(D4141_Y), .A(D4120_Q));
KC_NAND2_X1 D4142 ( .Y(D4142_Y), .B(D4139_Y), .A(D4122_Q));
KC_NAND2_X1 D4140 ( .Y(D4140_Y), .B(D4148_Y), .A(D4119_Q));
KC_NAND2_X1 D3992 ( .Y(D3992_Y), .B(D1407_Y), .A(D8471_Y));
KC_NAND2_X1 D3991 ( .Y(D3991_Y), .B(D8471_Y), .A(D1407_Y));
KC_NAND2_X1 D3987 ( .Y(D3987_Y), .B(D3881_Y), .A(D169_Y));
KC_NAND2_X1 D3986 ( .Y(D3986_Y), .B(D169_Y), .A(D6794_Y));
KC_NAND2_X1 D3839 ( .Y(D3839_Y), .B(D5387_Y), .A(D6794_Y));
KC_NAND2_X1 D3838 ( .Y(D3838_Y), .B(D8309_Y), .A(D3841_Y));
KC_NAND2_X1 D3837 ( .Y(D3837_Y), .B(D3841_Y), .A(D8309_Y));
KC_NAND2_X1 D3836 ( .Y(D3836_Y), .B(D3881_Y), .A(D5387_Y));
KC_NAND2_X1 D3714 ( .Y(D3714_Y), .B(D3713_Y), .A(D561_Y));
KC_NAND2_X1 D3594 ( .Y(D3594_Y), .B(D5020_Y), .A(D4882_Y));
KC_NAND2_X1 D3538 ( .Y(D3538_Y), .B(D4911_Y), .A(D3400_Y));
KC_NAND2_X1 D3537 ( .Y(D3537_Y), .B(D3533_Y), .A(D3540_Y));
KC_NAND2_X1 D3533 ( .Y(D3533_Y), .B(D1570_Y), .A(D3576_Q));
KC_NAND2_X1 D3520 ( .Y(D3520_Y), .B(D4911_Y), .A(D4874_Y));
KC_NAND2_X1 D3519 ( .Y(D3519_Y), .B(D3533_Y), .A(D4874_Y));
KC_NAND2_X1 D3516 ( .Y(D3516_Y), .B(D4911_Y), .A(D3599_Y));
KC_NAND2_X1 D3515 ( .Y(D3515_Y), .B(D3516_Y), .A(D3446_Y));
KC_NAND2_X1 D3508 ( .Y(D3508_Y), .B(D3413_Y), .A(D4985_Y));
KC_NAND2_X1 D3447 ( .Y(D3447_Y), .B(D4960_Y), .A(D1537_Y));
KC_NAND2_X1 D3439 ( .Y(D3439_Y), .B(D3447_Y), .A(D4915_Y));
KC_NAND2_X1 D3438 ( .Y(D3438_Y), .B(D3304_Y), .A(D1570_Y));
KC_NAND2_X1 D3429 ( .Y(D3429_Y), .B(D3428_Y), .A(D3388_Q));
KC_NAND2_X1 D3428 ( .Y(D3428_Y), .B(D3599_Y), .A(D3479_Y));
KC_NAND2_X1 D3427 ( .Y(D3427_Y), .B(D4903_Y), .A(D3432_Y));
KC_NAND2_X1 D3422 ( .Y(D3422_Y), .B(D3408_Y), .A(D446_Q));
KC_NAND2_X1 D3421 ( .Y(D3421_Y), .B(D3516_Y), .A(D4916_Y));
KC_NAND2_X1 D3420 ( .Y(D3420_Y), .B(D3432_Y), .A(D3430_Y));
KC_NAND2_X1 D3415 ( .Y(D3415_Y), .B(D3477_Y), .A(D1537_Y));
KC_NAND2_X1 D3414 ( .Y(D3414_Y), .B(D4960_Y), .A(D3416_Y));
KC_NAND2_X1 D3405 ( .Y(D3405_Y), .B(D3446_Y), .A(D3365_Y));
KC_NAND2_X1 D3331 ( .Y(D3331_Y), .B(D3209_Y), .A(D3346_Y));
KC_NAND2_X1 D3325 ( .Y(D3325_Y), .B(D3137_Y), .A(D3349_Y));
KC_NAND2_X1 D3304 ( .Y(D3304_Y), .B(D3374_Q), .A(D3375_Q));
KC_NAND2_X1 D3239 ( .Y(D3239_Y), .B(D1423_Y), .A(D3225_Y));
KC_NAND2_X1 D3237 ( .Y(D3237_Y), .B(D3282_Q), .A(D3281_Q));
KC_NAND2_X1 D3229 ( .Y(D3229_Y), .B(D1456_Y), .A(D3283_Q));
KC_NAND2_X1 D3221 ( .Y(D3221_Y), .B(D3368_Y), .A(D3270_Y));
KC_NAND2_X1 D3218 ( .Y(D3218_Y), .B(D3360_Y), .A(D3247_Y));
KC_NAND2_X1 D3214 ( .Y(D3214_Y), .B(D3329_Y), .A(D3360_Y));
KC_NAND2_X1 D3213 ( .Y(D3213_Y), .B(D4658_Y), .A(D3380_Y));
KC_NAND2_X1 D3206 ( .Y(D3206_Y), .B(D3215_Y), .A(D3368_Y));
KC_NAND2_X1 D3152 ( .Y(D3152_Y), .B(D3146_Y), .A(D3138_Y));
KC_NAND2_X1 D3151 ( .Y(D3151_Y), .B(D3185_Q), .A(D3188_Q));
KC_NAND2_X1 D3142 ( .Y(D3142_Y), .B(D3141_Y), .A(D3143_Y));
KC_NAND2_X1 D3141 ( .Y(D3141_Y), .B(D3040_Y), .A(D9345_Y));
KC_NAND2_X1 D3132 ( .Y(D3132_Y), .B(D3186_Q), .A(D3189_Q));
KC_NAND2_X1 D3119 ( .Y(D3119_Y), .B(D3137_Y), .A(D3124_Y));
KC_NAND2_X1 D3118 ( .Y(D3118_Y), .B(D3140_Y), .A(D3130_Y));
KC_NAND2_X1 D3107 ( .Y(D3107_Y), .B(D336_Y), .A(D3112_Y));
KC_NAND2_X1 D3030 ( .Y(D3030_Y), .B(D3024_Y), .A(D3025_Y));
KC_NAND2_X1 D3026 ( .Y(D3026_Y), .B(D3079_Q), .A(D3078_Q));
KC_NAND2_X1 D3019 ( .Y(D3019_Y), .B(D39_Y), .A(D3087_Y));
KC_NAND2_X1 D3014 ( .Y(D3014_Y), .B(D3015_Y), .A(D3079_Q));
KC_NAND2_X1 D3013 ( .Y(D3013_Y), .B(D3015_Y), .A(D44_Y));
KC_NAND2_X1 D2945 ( .Y(D2945_Y), .B(D1439_Y), .A(D2854_Y));
KC_NAND2_X1 D2944 ( .Y(D2944_Y), .B(D2825_Y), .A(D2857_Y));
KC_NAND2_X1 D2943 ( .Y(D2943_Y), .B(D1459_Y), .A(D2857_Y));
KC_NAND2_X1 D2942 ( .Y(D2942_Y), .B(D1439_Y), .A(D2857_Y));
KC_NAND2_X1 D2941 ( .Y(D2941_Y), .B(D2825_Y), .A(D2854_Y));
KC_NAND2_X1 D2940 ( .Y(D2940_Y), .B(D1459_Y), .A(D2854_Y));
KC_NAND2_X1 D2939 ( .Y(D2939_Y), .B(D2941_Y), .A(D2859_Y));
KC_NAND2_X1 D2935 ( .Y(D2935_Y), .B(D2944_Y), .A(D2824_Y));
KC_NAND2_X1 D2934 ( .Y(D2934_Y), .B(D2894_Y), .A(D2937_Y));
KC_NAND2_X1 D2932 ( .Y(D2932_Y), .B(D1435_Y), .A(D1488_Y));
KC_NAND2_X1 D2930 ( .Y(D2930_Y), .B(D2937_Y), .A(D2859_Y));
KC_NAND2_X1 D2929 ( .Y(D2929_Y), .B(D2985_Y), .A(D1438_Y));
KC_NAND2_X1 D2928 ( .Y(D2928_Y), .B(D2860_Y), .A(D2944_Y));
KC_NAND2_X1 D2927 ( .Y(D2927_Y), .B(D2945_Y), .A(D2859_Y));
KC_NAND2_X1 D2926 ( .Y(D2926_Y), .B(D1488_Y), .A(D1438_Y));
KC_NAND2_X1 D2925 ( .Y(D2925_Y), .B(D1435_Y), .A(D2985_Y));
KC_NAND2_X1 D2922 ( .Y(D2922_Y), .B(D2942_Y), .A(D2824_Y));
KC_NAND2_X1 D2921 ( .Y(D2921_Y), .B(D1438_Y), .A(D2987_Y));
KC_NAND2_X1 D2920 ( .Y(D2920_Y), .B(D2943_Y), .A(D2824_Y));
KC_NAND2_X1 D2919 ( .Y(D2919_Y), .B(D2986_Y), .A(D1438_Y));
KC_NAND2_X1 D2918 ( .Y(D2918_Y), .B(D2943_Y), .A(D2860_Y));
KC_NAND2_X1 D2917 ( .Y(D2917_Y), .B(D2942_Y), .A(D2860_Y));
KC_NAND2_X1 D2915 ( .Y(D2915_Y), .B(D2940_Y), .A(D2859_Y));
KC_NAND2_X1 D2914 ( .Y(D2914_Y), .B(D1490_Y), .A(D1438_Y));
KC_NAND2_X1 D2907 ( .Y(D2907_Y), .B(D1435_Y), .A(D1491_Y));
KC_NAND2_X1 D2906 ( .Y(D2906_Y), .B(D1491_Y), .A(D1438_Y));
KC_NAND2_X1 D2900 ( .Y(D2900_Y), .B(D2788_Y), .A(D2885_Q));
KC_NAND2_X1 D2850 ( .Y(D2850_Y), .B(D2858_Y), .A(D2852_Y));
KC_NAND2_X1 D2846 ( .Y(D2846_Y), .B(D1440_Y), .A(D2850_Y));
KC_NAND2_X1 D2838 ( .Y(D2838_Y), .B(D2822_Y), .A(D2836_Y));
KC_NAND2_X1 D2831 ( .Y(D2831_Y), .B(D4366_Y), .A(D2956_Y));
KC_NAND2_X1 D2825 ( .Y(D2825_Y), .B(D2885_Q), .A(D2884_Q));
KC_NAND2_X1 D2766 ( .Y(D2766_Y), .B(D2780_Y), .A(D2782_Y));
KC_NAND2_X1 D2753 ( .Y(D2753_Y), .B(D2850_Y), .A(D2744_Y));
KC_NAND2_X1 D2746 ( .Y(D2746_Y), .B(D2769_Y), .A(D2773_Y));
KC_NAND2_X1 D2745 ( .Y(D2745_Y), .B(D2747_Y), .A(D2741_Y));
KC_NAND2_X1 D2744 ( .Y(D2744_Y), .B(D2746_Y), .A(D1956_Y));
KC_NAND2_X1 D2715 ( .Y(D2715_Y), .B(D2750_Y), .A(D2725_Y));
KC_NAND2_X1 D2714 ( .Y(D2714_Y), .B(D2750_Y), .A(D2726_Y));
KC_NAND2_X1 D2713 ( .Y(D2713_Y), .B(D2750_Y), .A(D2730_Y));
KC_NAND2_X1 D2712 ( .Y(D2712_Y), .B(D2750_Y), .A(D2729_Y));
KC_NAND2_X1 D2711 ( .Y(D2711_Y), .B(D2750_Y), .A(D2724_Y));
KC_NAND2_X1 D2710 ( .Y(D2710_Y), .B(D2750_Y), .A(D2723_Y));
KC_NAND2_X1 D2709 ( .Y(D2709_Y), .B(D2750_Y), .A(D2731_Y));
KC_NAND2_X1 D2708 ( .Y(D2708_Y), .B(D2750_Y), .A(D2722_Y));
KC_NAND2_X1 D2707 ( .Y(D2707_Y), .B(D2750_Y), .A(D2732_Y));
KC_NAND2_X1 D2706 ( .Y(D2706_Y), .B(D2750_Y), .A(D2721_Y));
KC_NAND2_X1 D2705 ( .Y(D2705_Y), .B(D2750_Y), .A(D2733_Y));
KC_NAND2_X1 D2704 ( .Y(D2704_Y), .B(D2750_Y), .A(D2720_Y));
KC_NAND2_X1 D2703 ( .Y(D2703_Y), .B(D2750_Y), .A(D2734_Y));
KC_NAND2_X1 D2702 ( .Y(D2702_Y), .B(D2750_Y), .A(D2719_Y));
KC_NAND2_X1 D2701 ( .Y(D2701_Y), .B(D2750_Y), .A(D2735_Y));
KC_NAND2_X1 D2700 ( .Y(D2700_Y), .B(D2750_Y), .A(D2718_Y));
KC_NAND2_X1 D2691 ( .Y(D2691_Y), .B(D16665_Y), .A(D16599_Q));
KC_NAND2_X1 D2651 ( .Y(D2651_Y), .B(D16087_Y), .A(D16064_Y));
KC_NAND2_X1 D2650 ( .Y(D2650_Y), .B(D2651_Y), .A(D14654_Y));
KC_NAND2_X1 D2607 ( .Y(D2607_Y), .B(D2609_Y), .A(D15562_Y));
KC_NAND2_X1 D2606 ( .Y(D2606_Y), .B(D15471_Y), .A(D749_Y));
KC_NAND2_X1 D2595 ( .Y(D2595_Y), .B(D15861_S), .A(D15908_Y));
KC_NAND2_X1 D2593 ( .Y(D2593_Y), .B(D15271_Y), .A(D15270_Y));
KC_NAND2_X1 D2547 ( .Y(D2547_Y), .B(D14497_Y), .A(D2512_Y));
KC_NAND2_X1 D2546 ( .Y(D2546_Y), .B(D14497_Y), .A(D14501_Y));
KC_NAND2_X1 D2487 ( .Y(D2487_Y), .B(D13419_Y), .A(D13297_Y));
KC_NAND2_X1 D2478 ( .Y(D2478_Y), .B(D14518_Q), .A(D14711_Y));
KC_NAND2_X1 D2438 ( .Y(D2438_Y), .B(D13478_Y), .A(D13294_Y));
KC_NAND2_X1 D2436 ( .Y(D2436_Y), .B(D13294_Y), .A(D13318_Y));
KC_NAND2_X1 D2435 ( .Y(D2435_Y), .B(D14019_Y), .A(D13294_Y));
KC_NAND2_X1 D2426 ( .Y(D2426_Y), .B(D13466_Y), .A(D13464_Y));
KC_NAND2_X1 D2421 ( .Y(D2421_Y), .B(D13419_Y), .A(D13295_Y));
KC_NAND2_X1 D2420 ( .Y(D2420_Y), .B(D13419_Y), .A(D13297_Y));
KC_NAND2_X1 D2409 ( .Y(D2409_Y), .B(D2405_Y), .A(D2343_Y));
KC_NAND2_X1 D2408 ( .Y(D2408_Y), .B(D2312_Y), .A(D12659_Y));
KC_NAND2_X1 D2407 ( .Y(D2407_Y), .B(D7668_Y), .A(D2405_Y));
KC_NAND2_X1 D2401 ( .Y(D2401_Y), .B(D12919_Q), .A(D12870_Y));
KC_NAND2_X1 D2376 ( .Y(D2376_Y), .B(D12819_Y), .A(D12815_Y));
KC_NAND2_X1 D2372 ( .Y(D2372_Y), .B(D12997_Q), .A(D2375_Y));
KC_NAND2_X1 D2371 ( .Y(D2371_Y), .B(D2391_Q), .A(D2374_Y));
KC_NAND2_X1 D2370 ( .Y(D2370_Y), .B(D13552_Y), .A(D13578_Y));
KC_NAND2_X1 D2361 ( .Y(D2361_Y), .B(D12188_Y), .A(D2353_Y));
KC_NAND2_X1 D2329 ( .Y(D2329_Y), .B(D12137_Y), .A(D12131_Y));
KC_NAND2_X1 D2229 ( .Y(D2229_Y), .B(D8473_Y), .A(D6792_Y));
KC_NAND2_X1 D2136 ( .Y(D2136_Y), .B(D2862_Y), .A(D10232_Y));
KC_NAND2_X1 D2127 ( .Y(D2127_Y), .B(D245_Y), .A(D8948_Y));
KC_NAND2_X1 D2117 ( .Y(D2117_Y), .B(D1983_Y), .A(D10299_Q));
KC_NAND2_X1 D2109 ( .Y(D2109_Y), .B(D2061_Y), .A(D9672_Y));
KC_NAND2_X1 D2024 ( .Y(D2024_Y), .B(D8883_Y), .A(D272_Y));
KC_NAND2_X1 D2013 ( .Y(D2013_Y), .B(D8986_Y), .A(D9475_Y));
KC_NAND2_X1 D2002 ( .Y(D2002_Y), .B(D9147_Y), .A(D51_Y));
KC_NAND2_X1 D2001 ( .Y(D2001_Y), .B(D7631_Y), .A(D5981_Y));
KC_NAND2_X1 D1993 ( .Y(D1993_Y), .B(D7670_Y), .A(D6288_Y));
KC_NAND2_X1 D1992 ( .Y(D1992_Y), .B(D1985_Y), .A(D9398_Y));
KC_NAND2_X1 D1986 ( .Y(D1986_Y), .B(D1990_Y), .A(D8156_Y));
KC_NAND2_X1 D1985 ( .Y(D1985_Y), .B(D8105_Y), .A(D643_Y));
KC_NAND2_X1 D1887 ( .Y(D1887_Y), .B(D8877_Y), .A(D8748_Y));
KC_NAND2_X1 D1885 ( .Y(D1885_Y), .B(D7214_Y), .A(D1970_Y));
KC_NAND2_X1 D1880 ( .Y(D1880_Y), .B(D177_Y), .A(D7409_Q));
KC_NAND2_X1 D1879 ( .Y(D1879_Y), .B(D7329_Y), .A(D7442_Y));
KC_NAND2_X1 D1873 ( .Y(D1873_Y), .B(D8952_Q), .A(D7361_Y));
KC_NAND2_X1 D1865 ( .Y(D1865_Y), .B(D382_Y), .A(D7469_Y));
KC_NAND2_X1 D1858 ( .Y(D1858_Y), .B(D1856_Y), .A(D7944_Y));
KC_NAND2_X1 D1857 ( .Y(D1857_Y), .B(D7965_Y), .A(D1901_Y));
KC_NAND2_X1 D1856 ( .Y(D1856_Y), .B(D7927_Y), .A(D7948_Y));
KC_NAND2_X1 D1855 ( .Y(D1855_Y), .B(D7835_Y), .A(D7947_Y));
KC_NAND2_X1 D1849 ( .Y(D1849_Y), .B(D1922_Y), .A(D6483_Y));
KC_NAND2_X1 D1846 ( .Y(D1846_Y), .B(D9368_Y), .A(D1845_Y));
KC_NAND2_X1 D1844 ( .Y(D1844_Y), .B(D6580_Y), .A(D8240_Y));
KC_NAND2_X1 D1839 ( .Y(D1839_Y), .B(D1915_Y), .A(D8202_Y));
KC_NAND2_X1 D1837 ( .Y(D1837_Y), .B(D11325_Q), .A(D545_Y));
KC_NAND2_X1 D1836 ( .Y(D1836_Y), .B(D8279_Y), .A(D8401_Y));
KC_NAND2_X1 D1835 ( .Y(D1835_Y), .B(D6702_Y), .A(D2353_Y));
KC_NAND2_X1 D1822 ( .Y(D1822_Y), .B(D1645_Q), .A(D8212_Y));
KC_NAND2_X1 D1735 ( .Y(D1735_Y), .B(D5736_Y), .A(D5886_Y));
KC_NAND2_X1 D1734 ( .Y(D1734_Y), .B(D5881_Y), .A(D5736_Y));
KC_NAND2_X1 D1733 ( .Y(D1733_Y), .B(D5877_Y), .A(D5646_Y));
KC_NAND2_X1 D1732 ( .Y(D1732_Y), .B(D5738_Y), .A(D5877_Y));
KC_NAND2_X1 D1731 ( .Y(D1731_Y), .B(D5877_Y), .A(D6039_Y));
KC_NAND2_X1 D1724 ( .Y(D1724_Y), .B(D214_Y), .A(D7326_Y));
KC_NAND2_X1 D1722 ( .Y(D1722_Y), .B(D6113_Y), .A(D5852_Y));
KC_NAND2_X1 D1721 ( .Y(D1721_Y), .B(D7295_Y), .A(D5969_Y));
KC_NAND2_X1 D1720 ( .Y(D1720_Y), .B(D4454_Y), .A(D7305_Y));
KC_NAND2_X1 D1711 ( .Y(D1711_Y), .B(D6065_Y), .A(D4416_Y));
KC_NAND2_X1 D1710 ( .Y(D1710_Y), .B(D6062_Y), .A(D5872_Y));
KC_NAND2_X1 D1702 ( .Y(D1702_Y), .B(D1701_Y), .A(D4746_Y));
KC_NAND2_X1 D1698 ( .Y(D1698_Y), .B(D1700_Y), .A(D1699_Y));
KC_NAND2_X1 D1685 ( .Y(D1685_Y), .B(D10514_Y), .A(D1143_Y));
KC_NAND2_X1 D1684 ( .Y(D1684_Y), .B(D8466_Y), .A(D5599_Y));
KC_NAND2_X1 D1683 ( .Y(D1683_Y), .B(D8466_Y), .A(D7068_Y));
KC_NAND2_X1 D1674 ( .Y(D1674_Y), .B(D5141_Q), .A(D8212_Y));
KC_NAND2_X1 D1583 ( .Y(D1583_Y), .B(D8980_Y), .A(D4272_Y));
KC_NAND2_X1 D1582 ( .Y(D1582_Y), .B(D5985_Y), .A(D1591_Y));
KC_NAND2_X1 D1573 ( .Y(D1573_Y), .B(D4577_Y), .A(D4572_Y));
KC_NAND2_X1 D1569 ( .Y(D1569_Y), .B(D3446_Y), .A(D4985_Y));
KC_NAND2_X1 D1564 ( .Y(D1564_Y), .B(D4926_Y), .A(D4913_Y));
KC_NAND2_X1 D1556 ( .Y(D1556_Y), .B(D5479_Y), .A(D5480_Y));
KC_NAND2_X1 D1529 ( .Y(D1529_Y), .B(D2898_Y), .A(D1524_Q));
KC_NAND2_X1 D1528 ( .Y(D1528_Y), .B(D2766_Y), .A(D1529_Y));
KC_NAND2_X1 D1440 ( .Y(D1440_Y), .B(D1525_Y), .A(D1442_Y));
KC_NAND2_X1 D1439 ( .Y(D1439_Y), .B(D2821_Y), .A(D2885_Q));
KC_NAND2_X1 D1423 ( .Y(D1423_Y), .B(D3225_Y), .A(D1421_Y));
KC_NAND2_X1 D1413 ( .Y(D1413_Y), .B(D3881_Y), .A(D11308_Y));
KC_NAND2_X1 D1412 ( .Y(D1412_Y), .B(D561_Y), .A(D3713_Y));
KC_NAND2_X1 D1411 ( .Y(D1411_Y), .B(D11308_Y), .A(D6794_Y));
KC_NAND2_X1 D1406 ( .Y(D1406_Y), .B(D1320_Q), .A(D1400_Q));
KC_NAND2_X1 D1341 ( .Y(D1341_Y), .B(D16488_Y), .A(D16539_Y));
KC_NAND2_X1 D1340 ( .Y(D1340_Y), .B(D16613_Q), .A(D1374_Q));
KC_NAND2_X1 D981 ( .Y(D981_Y), .B(D11476_Y), .A(D11322_Y));
KC_NAND2_X1 D980 ( .Y(D980_Y), .B(D11322_Y), .A(D10861_Y));
KC_NAND2_X1 D961 ( .Y(D961_Y), .B(D13393_Y), .A(D12813_Y));
KC_NAND2_X1 D874 ( .Y(D874_Y), .B(D14025_Y), .A(D13312_Y));
KC_NAND2_X1 D863 ( .Y(D863_Y), .B(D6698_Y), .A(D8240_Y));
KC_NAND2_X1 D752 ( .Y(D752_Y), .B(D8887_Y), .A(D14813_Y));
KC_NAND2_X1 D749 ( .Y(D749_Y), .B(D14514_Y), .A(D15490_Y));
KC_NAND2_X1 D733 ( .Y(D733_Y), .B(D8240_Y), .A(D6693_Y));
KC_NAND2_X1 D639 ( .Y(D639_Y), .B(D13992_Q), .A(D13254_Y));
KC_NAND2_X1 D636 ( .Y(D636_Y), .B(D14513_Y), .A(D14624_Y));
KC_NAND2_X1 D635 ( .Y(D635_Y), .B(D14619_Y), .A(D14631_Y));
KC_NAND2_X1 D622 ( .Y(D622_Y), .B(D9421_Y), .A(D1984_Y));
KC_NAND2_X1 D570 ( .Y(D570_Y), .B(D16057_Y), .A(D15335_Y));
KC_NAND2_X1 D564 ( .Y(D564_Y), .B(D16062_Y), .A(D15335_Y));
KC_NAND2_X1 D560 ( .Y(D560_Y), .B(D12661_Y), .A(D161_Y));
KC_NAND2_X1 D471 ( .Y(D471_Y), .B(D1563_Y), .A(D5038_Y));
KC_NAND2_X1 D469 ( .Y(D469_Y), .B(D7839_Y), .A(D7920_Y));
KC_NAND2_X1 D434 ( .Y(D434_Y), .B(D9147_Y), .A(D7613_Y));
KC_NAND2_X1 D3391 ( .Y(D3391_Y), .B(D4846_Y), .A(D3385_Q));
KC_NAND2_X1 D405 ( .Y(D405_Y), .B(D4797_Y), .A(D3361_Y));
KC_NAND2_X1 D372 ( .Y(D372_Y), .B(D3234_Y), .A(D4687_Y));
KC_NAND2_X1 D371 ( .Y(D371_Y), .B(D4656_Y), .A(D4774_Y));
KC_NAND2_X1 D369 ( .Y(D369_Y), .B(D3214_Y), .A(D3218_Y));
KC_NAND2_X1 D339 ( .Y(D339_Y), .B(D4587_Y), .A(D6291_Y));
KC_NAND2_X1 D238 ( .Y(D238_Y), .B(D4267_Y), .A(D239_Q));
KC_NAND2_X1 D237 ( .Y(D237_Y), .B(D2815_Y), .A(D4235_Q));
KC_NAND2_X1 D216 ( .Y(D216_Y), .B(D8768_Y), .A(D8759_Y));
KC_NAND2_X1 D213 ( .Y(D213_Y), .B(D174_Y), .A(D7092_Y));
KC_NAND2_X1 D211 ( .Y(D211_Y), .B(D209_Y), .A(D8772_Y));
KC_NAND2_X1 D210 ( .Y(D210_Y), .B(D7276_Y), .A(D7234_Y));
KC_NAND2_X1 D204 ( .Y(D204_Y), .B(D7183_Y), .A(D9481_Y));
KC_NAND2_X1 D176 ( .Y(D176_Y), .B(D5649_Y), .A(D4092_Y));
KC_NAND2_X1 D89 ( .Y(D89_Y), .B(D13374_Y), .A(D16271_Y));
KC_NAND2_X1 D86 ( .Y(D86_Y), .B(D13419_Y), .A(D13295_Y));
KC_NAND2_X1 D73 ( .Y(D73_Y), .B(D6062_Y), .A(D275_Y));
KC_NAND2_X1 D69 ( .Y(D69_Y), .B(D4920_Y), .A(D3373_Q));
KC_NAND4_X1 D16654 ( .Y(D16654_Y), .D(D16658_Y), .C(D16609_Y),     .B(D1395_Q), .A(D16650_Q));
KC_NAND4_X1 D16624 ( .Y(D16624_Y), .D(D16655_Y), .C(D16657_Y),     .B(D1400_Q), .A(D16667_Y));
KC_NAND4_X1 D16623 ( .Y(D16623_Y), .D(D16652_Y), .C(D16667_Y),     .B(D16647_Y), .A(D14698_Y));
KC_NAND4_X1 D16600 ( .Y(D16600_Y), .D(D16590_Q), .C(D16564_Q),     .B(D16613_Q), .A(D1374_Q));
KC_NAND4_X1 D16571 ( .Y(D16571_Y), .D(D16564_Q), .C(D16611_Q),     .B(D16572_Y), .A(D16285_Y));
KC_NAND4_X1 D16570 ( .Y(D16570_Y), .D(D16533_Y), .C(D16489_Y),     .B(D16555_Q), .A(D16586_Y));
KC_NAND4_X1 D16523 ( .Y(D16523_Y), .D(D16499_Y), .C(D16528_Y),     .B(D16771_Y), .A(D1385_Q));
KC_NAND4_X1 D16519 ( .Y(D16519_Y), .D(D16001_Y), .C(D16504_Y),     .B(D16523_Y), .A(D16612_Y));
KC_NAND4_X1 D16500 ( .Y(D16500_Y), .D(D16488_Y), .C(D16536_Y),     .B(D16538_Y), .A(D1385_Q));
KC_NAND4_X1 D16495 ( .Y(D16495_Y), .D(D16505_Y), .C(D16549_Y),     .B(D16524_Y), .A(D16548_Y));
KC_NAND4_X1 D16490 ( .Y(D16490_Y), .D(D16488_Y), .C(D16379_Y),     .B(D16538_Y), .A(D16539_Y));
KC_NAND4_X1 D16489 ( .Y(D16489_Y), .D(D16549_Y), .C(D15958_Y),     .B(D14744_Y), .A(D16548_Y));
KC_NAND4_X1 D16442 ( .Y(D16442_Y), .D(D16454_Y), .C(D16422_Y),     .B(D16451_Y), .A(D16413_Y));
KC_NAND4_X1 D16437 ( .Y(D16437_Y), .D(D16452_Y), .C(D16451_Y),     .B(D1276_Y), .A(D16458_Y));
KC_NAND4_X1 D16432 ( .Y(D16432_Y), .D(D16425_Y), .C(D16426_Y),     .B(D16471_Q), .A(D16436_Y));
KC_NAND4_X1 D16431 ( .Y(D16431_Y), .D(D16433_Y), .C(D16425_Y),     .B(D16426_Y), .A(D1378_Q));
KC_NAND4_X1 D16428 ( .Y(D16428_Y), .D(D16408_Y), .C(D16398_Y),     .B(D16413_Y), .A(D16440_Y));
KC_NAND4_X1 D16427 ( .Y(D16427_Y), .D(D16454_Y), .C(D16460_Y),     .B(D15985_Y), .A(D16410_Y));
KC_NAND4_X1 D16424 ( .Y(D16424_Y), .D(D16425_Y), .C(D16433_Y),     .B(D1378_Q), .A(D1322_Q));
KC_NAND4_X1 D16423 ( .Y(D16423_Y), .D(D16425_Y), .C(D16426_Y),     .B(D1378_Q), .A(D16471_Q));
KC_NAND4_X1 D16421 ( .Y(D16421_Y), .D(D16460_Y), .C(D16422_Y),     .B(D16398_Y), .A(D16410_Y));
KC_NAND4_X1 D16416 ( .Y(D16416_Y), .D(D16438_Y), .C(D16426_Y),     .B(D16435_Y), .A(D16459_Q));
KC_NAND4_X1 D16263 ( .Y(D16263_Y), .D(D16256_Y), .C(D16274_Y),     .B(D16293_Q), .A(D2681_Q));
KC_NAND4_X1 D16259 ( .Y(D16259_Y), .D(D16265_Y), .C(D16274_Y),     .B(D16293_Q), .A(D16292_Q));
KC_NAND4_X1 D16190 ( .Y(D16190_Y), .D(D16458_Y), .C(D16192_Y),     .B(D15508_Y), .A(D16382_Y));
KC_NAND4_X1 D16064 ( .Y(D16064_Y), .D(D15327_Y), .C(D16094_Y),     .B(D16059_Y), .A(D15335_Y));
KC_NAND4_X1 D16063 ( .Y(D16063_Y), .D(D15282_Y), .C(D16094_Y),     .B(D16059_Y), .A(D15335_Y));
KC_NAND4_X1 D16055 ( .Y(D16055_Y), .D(D16072_Y), .C(D16094_Y),     .B(D15335_Y), .A(D16059_Y));
KC_NAND4_X1 D16048 ( .Y(D16048_Y), .D(D16054_Y), .C(D2590_Y),     .B(D16060_Y), .A(D16062_Y));
KC_NAND4_X1 D15966 ( .Y(D15966_Y), .D(D15915_Y), .C(D15179_Y),     .B(D15109_Y), .A(D1279_Y));
KC_NAND4_X1 D15887 ( .Y(D15887_Y), .D(D15880_Y), .C(D15879_Y),     .B(D15885_Y), .A(D15088_Y));
KC_NAND4_X1 D15881 ( .Y(D15881_Y), .D(D1228_Q), .C(D15998_Q),     .B(D15995_Q), .A(D15996_Q));
KC_NAND4_X1 D15835 ( .Y(D15835_Y), .D(D16389_Q), .C(D16364_Q),     .B(D16391_Q), .A(D16365_Q));
KC_NAND4_X1 D15822 ( .Y(D15822_Y), .D(D16369_Q), .C(D15872_Q),     .B(D16354_Q), .A(D15871_Q));
KC_NAND4_X1 D15819 ( .Y(D15819_Y), .D(D15946_Y), .C(D15989_Y),     .B(D15866_Y), .A(D1117_Y));
KC_NAND4_X1 D15714 ( .Y(D15714_Y), .D(D2600_Y), .C(D15712_Y),     .B(D2599_Y), .A(D15036_Y));
KC_NAND4_X1 D15288 ( .Y(D15288_Y), .D(D15278_Y), .C(D15310_Y),     .B(D15277_Y), .A(D15276_Y));
KC_NAND4_X1 D15269 ( .Y(D15269_Y), .D(D15436_Y), .C(D15333_Y),     .B(D2592_Y), .A(D16069_Y));
KC_NAND4_X1 D15171 ( .Y(D15171_Y), .D(D15233_Q), .C(D1386_Q),     .B(D15231_Q), .A(D15238_Q));
KC_NAND4_X1 D15170 ( .Y(D15170_Y), .D(D1278_Y), .C(D15168_Y),     .B(D15175_Y), .A(D15178_Y));
KC_NAND4_X1 D15091 ( .Y(D15091_Y), .D(D15085_Y), .C(D15087_Y),     .B(D15886_Y), .A(D15093_Y));
KC_NAND4_X1 D15089 ( .Y(D15089_Y), .D(D15086_Y), .C(D15104_Y),     .B(D14318_Y), .A(D14331_Y));
KC_NAND4_X1 D15042 ( .Y(D15042_Y), .D(D15832_Y), .C(D15816_Y),     .B(D15817_Y), .A(D15040_Y));
KC_NAND4_X1 D15037 ( .Y(D15037_Y), .D(D15034_Y), .C(D15030_Y),     .B(D15026_Y), .A(D14824_Y));
KC_NAND4_X1 D15031 ( .Y(D15031_Y), .D(D15033_Y), .C(D15015_Y),     .B(D15028_Y), .A(D14838_Y));
KC_NAND4_X1 D15022 ( .Y(D15022_Y), .D(D15035_Y), .C(D15017_Y),     .B(D15029_Y), .A(D14825_Y));
KC_NAND4_X1 D14959 ( .Y(D14959_Y), .D(D15797_Q), .C(D15711_Q),     .B(D1074_Q), .A(D14997_Q));
KC_NAND4_X1 D14952 ( .Y(D14952_Y), .D(D15726_Y), .C(D2535_Y),     .B(D14942_Y), .A(D15742_Y));
KC_NAND4_X1 D14940 ( .Y(D14940_Y), .D(D15737_Y), .C(D15736_Y),     .B(D15733_Y), .A(D14943_Y));
KC_NAND4_X1 D14929 ( .Y(D14929_Y), .D(D15719_Y), .C(D15718_Y),     .B(D15725_Y), .A(D14931_Y));
KC_NAND4_X1 D14926 ( .Y(D14926_Y), .D(D14936_Y), .C(D16318_Q),     .B(D16314_Q), .A(D15794_Q));
KC_NAND4_X1 D14923 ( .Y(D14923_Y), .D(D14960_Y), .C(D985_Y),     .B(D15095_Y), .A(D15038_Y));
KC_NAND4_X1 D14921 ( .Y(D14921_Y), .D(D14913_Y), .C(D14919_Y),     .B(D14917_Y), .A(D871_Y));
KC_NAND4_X1 D14843 ( .Y(D14843_Y), .D(D14844_Y), .C(D14865_Y),     .B(D14861_Y), .A(D14849_Y));
KC_NAND4_X1 D14842 ( .Y(D14842_Y), .D(D948_Y), .C(D14868_Y),     .B(D14910_Y), .A(D14159_Y));
KC_NAND4_X1 D14836 ( .Y(D14836_Y), .D(D14831_Y), .C(D14955_Y),     .B(D14834_Y), .A(D14822_Y));
KC_NAND4_X1 D14835 ( .Y(D14835_Y), .D(D14832_Y), .C(D14956_Y),     .B(D14818_Y), .A(D14823_Y));
KC_NAND4_X1 D14820 ( .Y(D14820_Y), .D(D14833_Y), .C(D2533_Y),     .B(D14819_Y), .A(D14125_Y));
KC_NAND4_X1 D14817 ( .Y(D14817_Y), .D(D925_Q), .C(D14874_Q),     .B(D15670_Q), .A(D1054_Q));
KC_NAND4_X1 D14753 ( .Y(D14753_Y), .D(D14704_Y), .C(D13968_Y),     .B(D14057_Y), .A(D14748_Y));
KC_NAND4_X1 D14636 ( .Y(D14636_Y), .D(D14632_Y), .C(D15418_Y),     .B(D14646_Y), .A(D14706_Y));
KC_NAND4_X1 D14618 ( .Y(D14618_Y), .D(D14652_Y), .C(D645_Y),     .B(D14668_Y), .A(D13931_Y));
KC_NAND4_X1 D14540 ( .Y(D14540_Y), .D(D14562_Y), .C(D14601_Q),     .B(D14520_Q), .A(D6976_Y));
KC_NAND4_X1 D14444 ( .Y(D14444_Y), .D(D14496_Q), .C(D15235_Q),     .B(D1379_Q), .A(D1380_Q));
KC_NAND4_X1 D14437 ( .Y(D14437_Y), .D(D14422_Y), .C(D14421_Y),     .B(D14434_Y), .A(D14420_Y));
KC_NAND4_X1 D14436 ( .Y(D14436_Y), .D(D14472_Y), .C(D14473_Y),     .B(D13797_Y), .A(D13755_Y));
KC_NAND4_X1 D14435 ( .Y(D14435_Y), .D(D13808_Q), .C(D14492_Q),     .B(D13759_Q), .A(D14495_Q));
KC_NAND4_X1 D14340 ( .Y(D14340_Y), .D(D14342_Y), .C(D13669_Y),     .B(D14341_Y), .A(D1184_Y));
KC_NAND4_X1 D14338 ( .Y(D14338_Y), .D(D15103_Y), .C(D15156_Y),     .B(D1181_Y), .A(D14397_Y));
KC_NAND4_X1 D14328 ( .Y(D14328_Y), .D(D14320_Y), .C(D14323_Y),     .B(D14319_Y), .A(D14423_Y));
KC_NAND4_X1 D14327 ( .Y(D14327_Y), .D(D1180_Y), .C(D14357_Y),     .B(D14325_Y), .A(D14333_Y));
KC_NAND4_X1 D14324 ( .Y(D14324_Y), .D(D1178_Y), .C(D2479_Y),     .B(D14326_Y), .A(D14339_Y));
KC_NAND4_X1 D14285 ( .Y(D14285_Y), .D(D1094_Y), .C(D2481_Y),     .B(D14272_Y), .A(D11100_Y));
KC_NAND4_X1 D14281 ( .Y(D14281_Y), .D(D14278_Y), .C(D2484_Y),     .B(D14280_Y), .A(D2483_Y));
KC_NAND4_X1 D14274 ( .Y(D14274_Y), .D(D14271_Y), .C(D2482_Y),     .B(D14283_Y), .A(D14273_Y));
KC_NAND4_X1 D14221 ( .Y(D14221_Y), .D(D14219_Y), .C(D14218_Y),     .B(D2490_Y), .A(D14213_Y));
KC_NAND4_X1 D14216 ( .Y(D14216_Y), .D(D989_Y), .C(D14214_Y),     .B(D14211_Y), .A(D14215_Y));
KC_NAND4_X1 D14208 ( .Y(D14208_Y), .D(D14230_Y), .C(D14269_Y),     .B(D14925_Y), .A(D14122_Y));
KC_NAND4_X1 D14207 ( .Y(D14207_Y), .D(D14265_Q), .C(D14242_Q),     .B(D14245_Q), .A(D14244_Q));
KC_NAND4_X1 D14203 ( .Y(D14203_Y), .D(D14205_Y), .C(D14270_Y),     .B(D14286_Y), .A(D14355_Y));
KC_NAND4_X1 D14202 ( .Y(D14202_Y), .D(D14234_Y), .C(D14235_Y),     .B(D14985_Y), .A(D14232_Y));
KC_NAND4_X1 D14201 ( .Y(D14201_Y), .D(D14267_Y), .C(D14268_Y),     .B(D15007_Y), .A(D15005_Y));
KC_NAND4_X1 D14131 ( .Y(D14131_Y), .D(D13495_Y), .C(D13519_Y),     .B(D1067_Y), .A(D14142_Y));
KC_NAND4_X1 D14120 ( .Y(D14120_Y), .D(D926_Q), .C(D14164_Q),     .B(D14167_Q), .A(D14241_Q));
KC_NAND4_X1 D13957 ( .Y(D13957_Y), .D(D14638_Y), .C(D13960_Y),     .B(D15393_Y), .A(D83_Y));
KC_NAND4_X1 D13956 ( .Y(D13956_Y), .D(D13980_Y), .C(D13962_Y),     .B(D13961_Y), .A(D638_Y));
KC_NAND4_X1 D13951 ( .Y(D13951_Y), .D(D13948_Y), .C(D13999_Y),     .B(D15381_Y), .A(D13981_Y));
KC_NAND4_X1 D13943 ( .Y(D13943_Y), .D(D14642_Y), .C(D13949_Y),     .B(D14623_Y), .A(D13944_Y));
KC_NAND4_X1 D13938 ( .Y(D13938_Y), .D(D14631_Y), .C(D13275_Q),     .B(D13946_Y), .A(D722_Q));
KC_NAND4_X1 D13896 ( .Y(D13896_Y), .D(D13177_Y), .C(D13959_Y),     .B(D571_Y), .A(D13881_Y));
KC_NAND4_X1 D13895 ( .Y(D13895_Y), .D(D13898_Y), .C(D13180_Y),     .B(D14737_Y), .A(D562_Y));
KC_NAND4_X1 D13894 ( .Y(D13894_Y), .D(D13897_Y), .C(D13891_Y),     .B(D14633_Y), .A(D13892_Y));
KC_NAND4_X1 D13893 ( .Y(D13893_Y), .D(D13899_Y), .C(D14041_Y),     .B(D13882_Y), .A(D13884_Y));
KC_NAND4_X1 D13888 ( .Y(D13888_Y), .D(D13903_Y), .C(D14752_Y),     .B(D13886_Y), .A(D13887_Y));
KC_NAND4_X1 D13885 ( .Y(D13885_Y), .D(D13176_Y), .C(D13927_Y),     .B(D13901_Y), .A(D565_Y));
KC_NAND4_X1 D13879 ( .Y(D13879_Y), .D(D13875_Y), .C(D14039_Y),     .B(D563_Y), .A(D13182_Y));
KC_NAND4_X1 D13878 ( .Y(D13878_Y), .D(D13880_Y), .C(D14741_Y),     .B(D13876_Y), .A(D13883_Y));
KC_NAND4_X1 D13845 ( .Y(D13845_Y), .D(D109_Y), .C(D349_Y),     .B(D13855_Y), .A(D13854_Y));
KC_NAND4_X1 D13715 ( .Y(D13715_Y), .D(D13806_Q), .C(D13827_Q),     .B(D13813_Q), .A(D1401_Q));
KC_NAND4_X1 D13644 ( .Y(D13644_Y), .D(D2474_Q), .C(D14316_Q),     .B(D14297_Q), .A(D14308_Q));
KC_NAND4_X1 D13465 ( .Y(D13465_Y), .D(D13533_Y), .C(D13522_Y),     .B(D1069_Y), .A(D13490_Y));
KC_NAND4_X1 D13427 ( .Y(D13427_Y), .D(D13537_Y), .C(D13518_Y),     .B(D1068_Y), .A(D13482_Y));
KC_NAND4_X1 D13418 ( .Y(D13418_Y), .D(D876_Y), .C(D2473_Y),     .B(D13626_Y), .A(D2444_Y));
KC_NAND4_X1 D13363 ( .Y(D13363_Y), .D(D13347_Y), .C(D13269_Q),     .B(D13267_Q), .A(D13333_Y));
KC_NAND4_X1 D13362 ( .Y(D13362_Y), .D(D13222_Y), .C(D13355_Y),     .B(D13363_Y), .A(D13354_Y));
KC_NAND4_X1 D13361 ( .Y(D13361_Y), .D(D13358_Y), .C(D13267_Q),     .B(D13333_Y), .A(D13398_Q));
KC_NAND4_X1 D13360 ( .Y(D13360_Y), .D(D13385_Y), .C(D12823_Y),     .B(D12797_Y), .A(D13363_Y));
KC_NAND4_X1 D13355 ( .Y(D13355_Y), .D(D13347_Y), .C(D13357_Y),     .B(D13352_Y), .A(D13335_Y));
KC_NAND4_X1 D13345 ( .Y(D13345_Y), .D(D13357_Y), .C(D13383_Y),     .B(D13353_Y), .A(D13398_Q));
KC_NAND4_X1 D13344 ( .Y(D13344_Y), .D(D2376_Y), .C(D13222_Y),     .B(D13345_Y), .A(D840_Y));
KC_NAND4_X1 D13343 ( .Y(D13343_Y), .D(D13353_Y), .C(D13398_Q),     .B(D13336_Y), .A(D13397_Q));
KC_NAND4_X1 D13342 ( .Y(D13342_Y), .D(D13370_Y), .C(D13345_Y),     .B(D13343_Y), .A(D13338_Y));
KC_NAND4_X1 D13338 ( .Y(D13338_Y), .D(D13357_Y), .C(D13335_Y),     .B(D13353_Y), .A(D13398_Q));
KC_NAND4_X1 D13239 ( .Y(D13239_Y), .D(D14628_Y), .C(D13237_Y),     .B(D14626_Y), .A(D13238_Y));
KC_NAND4_X1 D13230 ( .Y(D13230_Y), .D(D13240_Y), .C(D13965_Y),     .B(D13284_Y), .A(D14684_Y));
KC_NAND4_X1 D13183 ( .Y(D13183_Y), .D(D13900_Y), .C(D13181_Y),     .B(D14657_Y), .A(D13217_Y));
KC_NAND4_X1 D13152 ( .Y(D13152_Y), .D(D13169_Y), .C(D13167_Y),     .B(D12645_Y), .A(D12646_Y));
KC_NAND4_X1 D13113 ( .Y(D13113_Y), .D(D13128_Y), .C(D13132_Y),     .B(D12557_Y), .A(D13106_Y));
KC_NAND4_X1 D13111 ( .Y(D13111_Y), .D(D13125_Y), .C(D13112_Y),     .B(D1262_Y), .A(D13104_Y));
KC_NAND4_X1 D13103 ( .Y(D13103_Y), .D(D13123_Y), .C(D13101_Y),     .B(D12563_Y), .A(D13107_Y));
KC_NAND4_X1 D13074 ( .Y(D13074_Y), .D(D13131_Y), .C(D13092_Y),     .B(D13055_Y), .A(D13110_Y));
KC_NAND4_X1 D13073 ( .Y(D13073_Y), .D(D13126_Y), .C(D13076_Y),     .B(D13054_Y), .A(D13105_Y));
KC_NAND4_X1 D13072 ( .Y(D13072_Y), .D(D13127_Y), .C(D13069_Y),     .B(D13078_Y), .A(D13109_Y));
KC_NAND4_X1 D13067 ( .Y(D13067_Y), .D(D13130_Y), .C(D13063_Y),     .B(D13061_Y), .A(D13071_Y));
KC_NAND4_X1 D13066 ( .Y(D13066_Y), .D(D13121_Y), .C(D13068_Y),     .B(D13062_Y), .A(D2366_Y));
KC_NAND4_X1 D13058 ( .Y(D13058_Y), .D(D13124_Y), .C(D13065_Y),     .B(D13075_Y), .A(D13070_Y));
KC_NAND4_X1 D13057 ( .Y(D13057_Y), .D(D13122_Y), .C(D13064_Y),     .B(D13059_Y), .A(D2367_Y));
KC_NAND4_X1 D13056 ( .Y(D13056_Y), .D(D13133_Y), .C(D13077_Y),     .B(D13060_Y), .A(D13108_Y));
KC_NAND4_X1 D12959 ( .Y(D12959_Y), .D(D12966_Y), .C(D13005_Y),     .B(D13627_Y), .A(D13596_Y));
KC_NAND4_X1 D12954 ( .Y(D12954_Y), .D(D12962_Y), .C(D12999_Y),     .B(D13577_Y), .A(D13637_Y));
KC_NAND4_X1 D12948 ( .Y(D12948_Y), .D(D12961_Y), .C(D13002_Y),     .B(D13625_Y), .A(D13587_Y));
KC_NAND4_X1 D12943 ( .Y(D12943_Y), .D(D12941_Y), .C(D2397_Y),     .B(D2398_Y), .A(D13452_Y));
KC_NAND4_X1 D12880 ( .Y(D12880_Y), .D(D13469_Y), .C(D12876_Y),     .B(D12881_Y), .A(D12877_Y));
KC_NAND4_X1 D12871 ( .Y(D12871_Y), .D(D12971_Y), .C(D13516_Y),     .B(D12927_Y), .A(D12937_Y));
KC_NAND4_X1 D12801 ( .Y(D12801_Y), .D(D12799_Y), .C(D12809_Y),     .B(D12798_Y), .A(D12800_Y));
KC_NAND4_X1 D12710 ( .Y(D12710_Y), .D(D12813_Y), .C(D13268_Q),     .B(D12714_Y), .A(D12698_Y));
KC_NAND4_X1 D12657 ( .Y(D12657_Y), .D(D12325_Y), .C(D12716_Y),     .B(D12715_Y), .A(D12248_Y));
KC_NAND4_X1 D12624 ( .Y(D12624_Y), .D(D12652_Y), .C(D12635_Y),     .B(D12638_Y), .A(D12647_Y));
KC_NAND4_X1 D12622 ( .Y(D12622_Y), .D(D12641_Y), .C(D12644_Y),     .B(D12648_Y), .A(D12633_Y));
KC_NAND4_X1 D12621 ( .Y(D12621_Y), .D(D12639_Y), .C(D12640_Y),     .B(D12651_Y), .A(D16762_Y));
KC_NAND4_X1 D12570 ( .Y(D12570_Y), .D(D12587_Y), .C(D12556_Y),     .B(D12552_Y), .A(D12562_Y));
KC_NAND4_X1 D12569 ( .Y(D12569_Y), .D(D12591_Y), .C(D12565_Y),     .B(D12553_Y), .A(D12561_Y));
KC_NAND4_X1 D12568 ( .Y(D12568_Y), .D(D1372_Y), .C(D12554_Y),     .B(D12566_Y), .A(D12559_Y));
KC_NAND4_X1 D12567 ( .Y(D12567_Y), .D(D12590_Y), .C(D12564_Y),     .B(D12555_Y), .A(D12560_Y));
KC_NAND4_X1 D12538 ( .Y(D12538_Y), .D(D12616_Y), .C(D12523_Y),     .B(D12524_Y), .A(D12519_Y));
KC_NAND4_X1 D12537 ( .Y(D12537_Y), .D(D12589_Y), .C(D12516_Y),     .B(D12535_Y), .A(D12009_Y));
KC_NAND4_X1 D12530 ( .Y(D12530_Y), .D(D12592_Y), .C(D12532_Y),     .B(D12527_Y), .A(D1174_Y));
KC_NAND4_X1 D12529 ( .Y(D12529_Y), .D(D12595_Y), .C(D12522_Y),     .B(D12528_Y), .A(D12526_Y));
KC_NAND4_X1 D12525 ( .Y(D12525_Y), .D(D12593_Y), .C(D12515_Y),     .B(D12521_Y), .A(D12014_Y));
KC_NAND4_X1 D12520 ( .Y(D12520_Y), .D(D12586_Y), .C(D12514_Y),     .B(D12518_Y), .A(D12008_Y));
KC_NAND4_X1 D12517 ( .Y(D12517_Y), .D(D12594_Y), .C(D12533_Y),     .B(D12536_Y), .A(D12007_Y));
KC_NAND4_X1 D12493 ( .Y(D12493_Y), .D(D13048_Y), .C(D2368_Y),     .B(D12512_Y), .A(D12479_Y));
KC_NAND4_X1 D12492 ( .Y(D12492_Y), .D(D13047_Y), .C(D81_Y),     .B(D12475_Y), .A(D12480_Y));
KC_NAND4_X1 D12491 ( .Y(D12491_Y), .D(D12510_Y), .C(D13020_Y),     .B(D12478_Y), .A(D12485_Y));
KC_NAND4_X1 D12490 ( .Y(D12490_Y), .D(D1145_Y), .C(D13021_Y),     .B(D12481_Y), .A(D12486_Y));
KC_NAND4_X1 D12489 ( .Y(D12489_Y), .D(D13046_Y), .C(D978_Y),     .B(D12488_Y), .A(D2320_Y));
KC_NAND4_X1 D12484 ( .Y(D12484_Y), .D(D12509_Y), .C(D2315_Y),     .B(D12476_Y), .A(D12427_Y));
KC_NAND4_X1 D12483 ( .Y(D12483_Y), .D(D12508_Y), .C(D12487_Y),     .B(D12474_Y), .A(D12426_Y));
KC_NAND4_X1 D12446 ( .Y(D12446_Y), .D(D1047_Y), .C(D12444_Y),     .B(D2322_Y), .A(D12385_Y));
KC_NAND4_X1 D12440 ( .Y(D12440_Y), .D(D12470_Y), .C(D12445_Y),     .B(D12434_Y), .A(D12438_Y));
KC_NAND4_X1 D12439 ( .Y(D12439_Y), .D(D12469_Y), .C(D12441_Y),     .B(D12433_Y), .A(D12437_Y));
KC_NAND4_X1 D12436 ( .Y(D12436_Y), .D(D12990_Y), .C(D12428_Y),     .B(D2317_Y), .A(D12432_Y));
KC_NAND4_X1 D12431 ( .Y(D12431_Y), .D(D12989_Y), .C(D12940_Y),     .B(D2316_Y), .A(D12430_Y));
KC_NAND4_X1 D12423 ( .Y(D12423_Y), .D(D12411_Y), .C(D12388_Y),     .B(D2323_Y), .A(D12386_Y));
KC_NAND4_X1 D12391 ( .Y(D12391_Y), .D(D12412_Y), .C(D12392_Y),     .B(D12390_Y), .A(D12387_Y));
KC_NAND4_X1 D12381 ( .Y(D12381_Y), .D(D2354_Y), .C(D12389_Y),     .B(D12377_Y), .A(D12383_Y));
KC_NAND4_X1 D12380 ( .Y(D12380_Y), .D(D12413_Y), .C(D12376_Y),     .B(D12384_Y), .A(D12382_Y));
KC_NAND4_X1 D12375 ( .Y(D12375_Y), .D(D12471_Y), .C(D12443_Y),     .B(D12378_Y), .A(D12374_Y));
KC_NAND4_X1 D12324 ( .Y(D12324_Y), .D(D12359_Q), .C(D12368_Q),     .B(D12358_Q), .A(D12274_Q));
KC_NAND4_X1 D12311 ( .Y(D12311_Y), .D(D12342_Q), .C(D2355_Q),     .B(D12416_Q), .A(D12351_Q));
KC_NAND4_X1 D12310 ( .Y(D12310_Y), .D(D12343_Q), .C(D12348_Q),     .B(D12346_Q), .A(D12367_Q));
KC_NAND4_X1 D12255 ( .Y(D12255_Y), .D(D2311_Y), .C(D12207_Y),     .B(D11660_Y), .A(D2310_Y));
KC_NAND4_X1 D12246 ( .Y(D12246_Y), .D(D12266_Y), .C(D12737_Y),     .B(D12265_Y), .A(D12264_Y));
KC_NAND4_X1 D12244 ( .Y(D12244_Y), .D(D12335_Y), .C(D653_Y),     .B(D12334_Y), .A(D12307_Y));
KC_NAND4_X1 D12205 ( .Y(D12205_Y), .D(D10179_Y), .C(D11660_Y),     .B(D12193_Y), .A(D10177_Y));
KC_NAND4_X1 D12204 ( .Y(D12204_Y), .D(D16130_Y), .C(D12744_Y),     .B(D12232_Y), .A(D12221_Y));
KC_NAND4_X1 D12186 ( .Y(D12186_Y), .D(D12187_Y), .C(D2363_Y),     .B(D9371_Y), .A(D12213_Y));
KC_NAND4_X1 D12133 ( .Y(D12133_Y), .D(D511_Y), .C(D2342_Y),     .B(D12642_Y), .A(D12230_Y));
KC_NAND4_X1 D12077 ( .Y(D12077_Y), .D(D12101_Y), .C(D12075_Y),     .B(D12062_Y), .A(D12078_Y));
KC_NAND4_X1 D12072 ( .Y(D12072_Y), .D(D12099_Y), .C(D12081_Y),     .B(D12064_Y), .A(D12083_Y));
KC_NAND4_X1 D12071 ( .Y(D12071_Y), .D(D12098_Y), .C(D12068_Y),     .B(D12066_Y), .A(D12079_Y));
KC_NAND4_X1 D12070 ( .Y(D12070_Y), .D(D12097_Y), .C(D12080_Y),     .B(D12063_Y), .A(D12076_Y));
KC_NAND4_X1 D12067 ( .Y(D12067_Y), .D(D12100_Y), .C(D12082_Y),     .B(D12065_Y), .A(D12073_Y));
KC_NAND4_X1 D12061 ( .Y(D12061_Y), .D(D12124_Y), .C(D12069_Y),     .B(D1261_Y), .A(D12074_Y));
KC_NAND4_X1 D12022 ( .Y(D12022_Y), .D(D12588_Y), .C(D12531_Y),     .B(D12534_Y), .A(D12021_Y));
KC_NAND4_X1 D12004 ( .Y(D12004_Y), .D(D12103_Y), .C(D12002_Y),     .B(D12019_Y), .A(D11998_Y));
KC_NAND4_X1 D12003 ( .Y(D12003_Y), .D(D12102_Y), .C(D12001_Y),     .B(D11997_Y), .A(D12020_Y));
KC_NAND4_X1 D11947 ( .Y(D11947_Y), .D(D11985_Y), .C(D11883_Y),     .B(D2268_Y), .A(D11892_Y));
KC_NAND4_X1 D11900 ( .Y(D11900_Y), .D(D11927_Y), .C(D11899_Y),     .B(D11894_Y), .A(D11897_Y));
KC_NAND4_X1 D11888 ( .Y(D11888_Y), .D(D11986_Y), .C(D11880_Y),     .B(D11885_Y), .A(D11890_Y));
KC_NAND4_X1 D11887 ( .Y(D11887_Y), .D(D11987_Y), .C(D11884_Y),     .B(D11879_Y), .A(D11891_Y));
KC_NAND4_X1 D11878 ( .Y(D11878_Y), .D(D11873_Y), .C(D11830_Y),     .B(D11828_Y), .A(D11839_Y));
KC_NAND4_X1 D11837 ( .Y(D11837_Y), .D(D11872_Y), .C(D11833_Y),     .B(D11831_Y), .A(D11841_Y));
KC_NAND4_X1 D11834 ( .Y(D11834_Y), .D(D11874_Y), .C(D11829_Y),     .B(D11824_Y), .A(D11840_Y));
KC_NAND4_X1 D11827 ( .Y(D11827_Y), .D(D11877_Y), .C(D11821_Y),     .B(D11819_Y), .A(D11838_Y));
KC_NAND4_X1 D11826 ( .Y(D11826_Y), .D(D11876_Y), .C(D11820_Y),     .B(D11822_Y), .A(D11835_Y));
KC_NAND4_X1 D11815 ( .Y(D11815_Y), .D(D11875_Y), .C(D11823_Y),     .B(D11825_Y), .A(D11836_Y));
KC_NAND4_X1 D11771 ( .Y(D11771_Y), .D(D11808_Y), .C(D11763_Y),     .B(D11773_Y), .A(D11769_Y));
KC_NAND4_X1 D11770 ( .Y(D11770_Y), .D(D11810_Y), .C(D11765_Y),     .B(D11686_Y), .A(D11768_Y));
KC_NAND4_X1 D11767 ( .Y(D11767_Y), .D(D12353_Q), .C(D12352_Q),     .B(D12349_Q), .A(D12350_Q));
KC_NAND4_X1 D11762 ( .Y(D11762_Y), .D(D11807_Y), .C(D11750_Y),     .B(D11757_Y), .A(D11747_Y));
KC_NAND4_X1 D11761 ( .Y(D11761_Y), .D(D2299_Y), .C(D11748_Y),     .B(D11759_Y), .A(D11751_Y));
KC_NAND4_X1 D11760 ( .Y(D11760_Y), .D(D11809_Y), .C(D11758_Y),     .B(D11756_Y), .A(D11745_Y));
KC_NAND4_X1 D11754 ( .Y(D11754_Y), .D(D2298_Y), .C(D11740_Y),     .B(D11755_Y), .A(D11746_Y));
KC_NAND4_X1 D11753 ( .Y(D11753_Y), .D(D11805_Y), .C(D11741_Y),     .B(D11749_Y), .A(D11752_Y));
KC_NAND4_X1 D11744 ( .Y(D11744_Y), .D(D11806_Y), .C(D11739_Y),     .B(D11743_Y), .A(D11742_Y));
KC_NAND4_X1 D11709 ( .Y(D11709_Y), .D(D11664_Y), .C(D11708_Y),     .B(D11707_Y), .A(D11692_Y));
KC_NAND4_X1 D11704 ( .Y(D11704_Y), .D(D2305_Y), .C(D11702_Y),     .B(D11701_Y), .A(D11689_Y));
KC_NAND4_X1 D11699 ( .Y(D11699_Y), .D(D11730_Y), .C(D11698_Y),     .B(D11705_Y), .A(D11696_Y));
KC_NAND4_X1 D11697 ( .Y(D11697_Y), .D(D11729_Y), .C(D11703_Y),     .B(D11695_Y), .A(D11691_Y));
KC_NAND4_X1 D11683 ( .Y(D11683_Y), .D(D11728_Y), .C(D11685_Y),     .B(D11688_Y), .A(D11680_Y));
KC_NAND4_X1 D11682 ( .Y(D11682_Y), .D(D11727_Y), .C(D11684_Y),     .B(D11687_Y), .A(D11681_Y));
KC_NAND4_X1 D11428 ( .Y(D11428_Y), .D(D11403_Y), .C(D1086_Y),     .B(D11427_Y), .A(D10968_Y));
KC_NAND4_X1 D11350 ( .Y(D11350_Y), .D(D11404_Y), .C(D79_Y),     .B(D1085_Y), .A(D10977_Y));
KC_NAND4_X1 D11222 ( .Y(D11222_Y), .D(D11132_Y), .C(D11215_Y),     .B(D11136_Y), .A(D11226_Y));
KC_NAND4_X1 D11218 ( .Y(D11218_Y), .D(D11278_Y), .C(D11211_Y),     .B(D628_Y), .A(D748_Y));
KC_NAND4_X1 D11217 ( .Y(D11217_Y), .D(D11277_Y), .C(D11216_Y),     .B(D11225_Y), .A(D11220_Y));
KC_NAND4_X1 D11214 ( .Y(D11214_Y), .D(D11130_Y), .C(D11213_Y),     .B(D626_Y), .A(D11224_Y));
KC_NAND4_X1 D11140 ( .Y(D11140_Y), .D(D11131_Y), .C(D11221_Y),     .B(D11137_Y), .A(D11138_Y));
KC_NAND4_X1 D11139 ( .Y(D11139_Y), .D(D604_Y), .C(D11219_Y),     .B(D10668_Y), .A(D11223_Y));
KC_NAND4_X1 D11058 ( .Y(D11058_Y), .D(D11111_Y), .C(D11059_Y),     .B(D11096_Y), .A(D10587_Y));
KC_NAND4_X1 D10978 ( .Y(D10978_Y), .D(D10957_Y), .C(D2185_Y),     .B(D10970_Y), .A(D10969_Y));
KC_NAND4_X1 D10962 ( .Y(D10962_Y), .D(D140_Y), .C(D10934_Y),     .B(D10932_Y), .A(D10933_Y));
KC_NAND4_X1 D10935 ( .Y(D10935_Y), .D(D11344_Y), .C(D10931_Y),     .B(D2198_Y), .A(D2192_Y));
KC_NAND4_X1 D10929 ( .Y(D10929_Y), .D(D1045_Y), .C(D10918_Y),     .B(D10920_Y), .A(D10925_Y));
KC_NAND4_X1 D10926 ( .Y(D10926_Y), .D(D10961_Y), .C(D10922_Y),     .B(D10921_Y), .A(D10927_Y));
KC_NAND4_X1 D10916 ( .Y(D10916_Y), .D(D11406_Y), .C(D10914_Y),     .B(D10906_Y), .A(D10974_Y));
KC_NAND4_X1 D10911 ( .Y(D10911_Y), .D(D10959_Y), .C(D10909_Y),     .B(D10900_Y), .A(D2182_Y));
KC_NAND4_X1 D10908 ( .Y(D10908_Y), .D(D10958_Y), .C(D10915_Y),     .B(D10907_Y), .A(D10973_Y));
KC_NAND4_X1 D10901 ( .Y(D10901_Y), .D(D10960_Y), .C(D10910_Y),     .B(D10899_Y), .A(D2181_Y));
KC_NAND4_X1 D10845 ( .Y(D10845_Y), .D(D923_Y), .C(D2194_Y),     .B(D10837_Y), .A(D10832_Y));
KC_NAND4_X1 D10841 ( .Y(D10841_Y), .D(D11343_Y), .C(D10835_Y),     .B(D10834_Y), .A(D10840_Y));
KC_NAND4_X1 D10839 ( .Y(D10839_Y), .D(D922_Y), .C(D2196_Y),     .B(D10836_Y), .A(D10833_Y));
KC_NAND4_X1 D10760 ( .Y(D10760_Y), .D(D10657_Y), .C(D10752_Y),     .B(D10670_Y), .A(D10755_Y));
KC_NAND4_X1 D10756 ( .Y(D10756_Y), .D(D10659_Y), .C(D10661_Y),     .B(D10669_Y), .A(D10662_Y));
KC_NAND4_X1 D10754 ( .Y(D10754_Y), .D(D602_Y), .C(D747_Y),     .B(D10665_Y), .A(D10759_Y));
KC_NAND4_X1 D10699 ( .Y(D10699_Y), .D(D2225_Y), .C(D10703_Y),     .B(D10689_Y), .A(D10683_Y));
KC_NAND4_X1 D10698 ( .Y(D10698_Y), .D(D2224_Y), .C(D10702_Y),     .B(D10690_Y), .A(D10684_Y));
KC_NAND4_X1 D10697 ( .Y(D10697_Y), .D(D601_Y), .C(D10695_Y),     .B(D10682_Y), .A(D10696_Y));
KC_NAND4_X1 D10692 ( .Y(D10692_Y), .D(D10654_Y), .C(D10694_Y),     .B(D10700_Y), .A(D10686_Y));
KC_NAND4_X1 D10691 ( .Y(D10691_Y), .D(D10658_Y), .C(D10671_Y),     .B(D10685_Y), .A(D10678_Y));
KC_NAND4_X1 D10680 ( .Y(D10680_Y), .D(D10655_Y), .C(D10673_Y),     .B(D10677_Y), .A(D10679_Y));
KC_NAND4_X1 D10676 ( .Y(D10676_Y), .D(D10656_Y), .C(D10758_Y),     .B(D10666_Y), .A(D10667_Y));
KC_NAND4_X1 D10675 ( .Y(D10675_Y), .D(D11129_Y), .C(D630_Y),     .B(D10674_Y), .A(D10687_Y));
KC_NAND4_X1 D10591 ( .Y(D10591_Y), .D(D10626_Y), .C(D1266_Y),     .B(D10574_Y), .A(D10586_Y));
KC_NAND4_X1 D10590 ( .Y(D10590_Y), .D(D10628_Y), .C(D11061_Y),     .B(D10589_Y), .A(D10575_Y));
KC_NAND4_X1 D10585 ( .Y(D10585_Y), .D(D11087_Y), .C(D10582_Y),     .B(D10581_Y), .A(D2112_Y));
KC_NAND4_X1 D10584 ( .Y(D10584_Y), .D(D10623_Y), .C(D10588_Y),     .B(D10566_Y), .A(D10567_Y));
KC_NAND4_X1 D10583 ( .Y(D10583_Y), .D(D11086_Y), .C(D10580_Y),     .B(D1263_Y), .A(D10573_Y));
KC_NAND4_X1 D10579 ( .Y(D10579_Y), .D(D1371_Y), .C(D10576_Y),     .B(D1260_Y), .A(D10577_Y));
KC_NAND4_X1 D10569 ( .Y(D10569_Y), .D(D10619_Y), .C(D1258_Y),     .B(D10564_Y), .A(D9872_Y));
KC_NAND4_X1 D10568 ( .Y(D10568_Y), .D(D10620_Y), .C(D9863_Y),     .B(D9858_Y), .A(D10572_Y));
KC_NAND4_X1 D10565 ( .Y(D10565_Y), .D(D10625_Y), .C(D10578_Y),     .B(D10571_Y), .A(D10570_Y));
KC_NAND4_X1 D10531 ( .Y(D10531_Y), .D(D10556_Y), .C(D10537_Y),     .B(D10529_Y), .A(D10561_Y));
KC_NAND4_X1 D10530 ( .Y(D10530_Y), .D(D10557_Y), .C(D10538_Y),     .B(D10528_Y), .A(D10526_Y));
KC_NAND4_X1 D10522 ( .Y(D10522_Y), .D(D2164_Y), .C(D1168_Y),     .B(D10525_Y), .A(D10523_Y));
KC_NAND4_X1 D10521 ( .Y(D10521_Y), .D(D2165_Y), .C(D9802_Y),     .B(D1169_Y), .A(D10524_Y));
KC_NAND4_X1 D10471 ( .Y(D10471_Y), .D(D1146_Y), .C(D10533_Y),     .B(D10469_Y), .A(D2129_Y));
KC_NAND4_X1 D10470 ( .Y(D10470_Y), .D(D11008_Y), .C(D10540_Y),     .B(D10468_Y), .A(D10461_Y));
KC_NAND4_X1 D10402 ( .Y(D10402_Y), .D(D10437_Y), .C(D10401_Y),     .B(D10395_Y), .A(D10380_Y));
KC_NAND4_X1 D10400 ( .Y(D10400_Y), .D(D10436_Y), .C(D10403_Y),     .B(D10445_Y), .A(D10381_Y));
KC_NAND4_X1 D10399 ( .Y(D10399_Y), .D(D1046_Y), .C(D10396_Y),     .B(D10441_Y), .A(D10377_Y));
KC_NAND4_X1 D10391 ( .Y(D10391_Y), .D(D10435_Y), .C(D10919_Y),     .B(D10390_Y), .A(D2113_Y));
KC_NAND4_X1 D10385 ( .Y(D10385_Y), .D(D10439_Y), .C(D10443_Y),     .B(D10442_Y), .A(D974_Y));
KC_NAND4_X1 D10384 ( .Y(D10384_Y), .D(D10438_Y), .C(D10386_Y),     .B(D10379_Y), .A(D10378_Y));
KC_NAND4_X1 D10383 ( .Y(D10383_Y), .D(D10440_Y), .C(D10398_Y),     .B(D10392_Y), .A(D10382_Y));
KC_NAND4_X1 D10376 ( .Y(D10376_Y), .D(D10432_Y), .C(D10397_Y),     .B(D10393_Y), .A(D10375_Y));
KC_NAND4_X1 D10200 ( .Y(D10200_Y), .D(D603_Y), .C(D10693_Y),     .B(D629_Y), .A(D10688_Y));
KC_NAND4_X1 D10194 ( .Y(D10194_Y), .D(D10213_Y), .C(D2151_Y),     .B(D10286_Y), .A(D10211_Y));
KC_NAND4_X1 D10193 ( .Y(D10193_Y), .D(D15457_Y), .C(D15460_Y),     .B(D9453_Y), .A(D10212_Y));
KC_NAND4_X1 D10153 ( .Y(D10153_Y), .D(D10157_Y), .C(D10160_Y),     .B(D10158_Y), .A(D481_Y));
KC_NAND4_X1 D10084 ( .Y(D10084_Y), .D(D9012_Y), .C(D9118_Y),     .B(D8904_Y), .A(D8972_Y));
KC_NAND4_X1 D10038 ( .Y(D10038_Y), .D(D10011_Y), .C(D10037_Y),     .B(D8907_Y), .A(D2125_Y));
KC_NAND4_X1 D10035 ( .Y(D10035_Y), .D(D9013_Y), .C(D8950_Y),     .B(D8949_Y), .A(D10045_Y));
KC_NAND4_X1 D10034 ( .Y(D10034_Y), .D(D9015_Y), .C(D10044_Y),     .B(D10043_Y), .A(D8973_Y));
KC_NAND4_X1 D10020 ( .Y(D10020_Y), .D(D10021_Y), .C(D10017_Y),     .B(D8853_Y), .A(D10019_Y));
KC_NAND4_X1 D9998 ( .Y(D9998_Y), .D(D9995_Y), .C(D10002_Y),     .B(D8870_Y), .A(D9989_Y));
KC_NAND4_X1 D9994 ( .Y(D9994_Y), .D(D9999_Y), .C(D9992_Y), .B(D8871_Y),     .A(D2126_Y));
KC_NAND4_X1 D9894 ( .Y(D9894_Y), .D(D10621_Y), .C(D9891_Y),     .B(D9851_Y), .A(D9873_Y));
KC_NAND4_X1 D9893 ( .Y(D9893_Y), .D(D9910_Y), .C(D9855_Y), .B(D9854_Y),     .A(D8623_Y));
KC_NAND4_X1 D9874 ( .Y(D9874_Y), .D(D10627_Y), .C(D9865_Y),     .B(D9859_Y), .A(D9866_Y));
KC_NAND4_X1 D9871 ( .Y(D9871_Y), .D(D10622_Y), .C(D9867_Y),     .B(D9852_Y), .A(D9868_Y));
KC_NAND4_X1 D9870 ( .Y(D9870_Y), .D(D9912_Y), .C(D9861_Y), .B(D9853_Y),     .A(D9869_Y));
KC_NAND4_X1 D9862 ( .Y(D9862_Y), .D(D10624_Y), .C(D9864_Y),     .B(D9860_Y), .A(D9875_Y));
KC_NAND4_X1 D9823 ( .Y(D9823_Y), .D(D9847_Y), .C(D9805_Y), .B(D9821_Y),     .A(D9818_Y));
KC_NAND4_X1 D9822 ( .Y(D9822_Y), .D(D9848_Y), .C(D9800_Y), .B(D9816_Y),     .A(D9817_Y));
KC_NAND4_X1 D9820 ( .Y(D9820_Y), .D(D9845_Y), .C(D9799_Y), .B(D9815_Y),     .A(D9814_Y));
KC_NAND4_X1 D9811 ( .Y(D9811_Y), .D(D9844_Y), .C(D9803_Y), .B(D9813_Y),     .A(D9804_Y));
KC_NAND4_X1 D9810 ( .Y(D9810_Y), .D(D9846_Y), .C(D9806_Y), .B(D9819_Y),     .A(D9808_Y));
KC_NAND4_X1 D9809 ( .Y(D9809_Y), .D(D9843_Y), .C(D9801_Y), .B(D9812_Y),     .A(D9807_Y));
KC_NAND4_X1 D9678 ( .Y(D9678_Y), .D(D2088_Y), .C(D9677_Y), .B(D9665_Y),     .A(D9653_Y));
KC_NAND4_X1 D9671 ( .Y(D9671_Y), .D(D10434_Y), .C(D9679_Y),     .B(D9662_Y), .A(D9655_Y));
KC_NAND4_X1 D9670 ( .Y(D9670_Y), .D(D10433_Y), .C(D9680_Y),     .B(D9669_Y), .A(D9652_Y));
KC_NAND4_X1 D9668 ( .Y(D9668_Y), .D(D9619_Y), .C(D9676_Y), .B(D9663_Y),     .A(D9656_Y));
KC_NAND4_X1 D9667 ( .Y(D9667_Y), .D(D2089_Y), .C(D9675_Y), .B(D9659_Y),     .A(D9654_Y));
KC_NAND4_X1 D9666 ( .Y(D9666_Y), .D(D138_Y), .C(D9673_Y), .B(D9664_Y),     .A(D9650_Y));
KC_NAND4_X1 D9661 ( .Y(D9661_Y), .D(D2087_Y), .C(D9674_Y), .B(D9658_Y),     .A(D9651_Y));
KC_NAND4_X1 D9660 ( .Y(D9660_Y), .D(D9618_Y), .C(D9594_Y), .B(D9657_Y),     .A(D9649_Y));
KC_NAND4_X1 D9525 ( .Y(D9525_Y), .D(D1991_Y), .C(D9575_Q), .B(D9579_Q),     .A(D9544_Y));
KC_NAND4_X1 D9518 ( .Y(D9518_Y), .D(D9514_Y), .C(D9528_Y), .B(D9575_Q),     .A(D9544_Y));
KC_NAND4_X1 D9517 ( .Y(D9517_Y), .D(D9507_Y), .C(D643_Y), .B(D9578_Q),     .A(D9577_Q));
KC_NAND4_X1 D9515 ( .Y(D9515_Y), .D(D2101_Y), .C(D10265_Y),     .B(D9552_Y), .A(D9546_Y));
KC_NAND4_X1 D9505 ( .Y(D9505_Y), .D(D9501_Y), .C(D9528_Y), .B(D9514_Y),     .A(D9597_Y));
KC_NAND4_X1 D9411 ( .Y(D9411_Y), .D(D9462_Y), .C(D9461_Y), .B(D9466_Y),     .A(D9467_Y));
KC_NAND4_X1 D9410 ( .Y(D9410_Y), .D(D9465_Y), .C(D9464_Y), .B(D2074_Y),     .A(D9455_Y));
KC_NAND4_X1 D9401 ( .Y(D9401_Y), .D(D9419_Y), .C(D9400_Y), .B(D8083_Y),     .A(D714_Q));
KC_NAND4_X1 D9372 ( .Y(D9372_Y), .D(D6285_Y), .C(D6281_Y), .B(D9378_Y),     .A(D11660_Y));
KC_NAND4_X1 D9370 ( .Y(D9370_Y), .D(D9380_Y), .C(D9794_Y), .B(D9794_Y),     .A(D8056_Y));
KC_NAND4_X1 D9365 ( .Y(D9365_Y), .D(D10180_Y), .C(D6285_Y),     .B(D8015_Y), .A(D9378_Y));
KC_NAND4_X1 D9364 ( .Y(D9364_Y), .D(D4747_Y), .C(D263_Y), .B(D9368_Y),     .A(D10177_Y));
KC_NAND4_X1 D9363 ( .Y(D9363_Y), .D(D392_Y), .C(D7669_Y), .B(D6288_Y),     .A(D10177_Y));
KC_NAND4_X1 D9343 ( .Y(D9343_Y), .D(D4540_Y), .C(D837_Q), .B(D2103_Q),     .A(D486_Q));
KC_NAND4_X1 D9241 ( .Y(D9241_Y), .D(D1787_Y), .C(D7626_Y), .B(D9242_Y),     .A(D9258_Y));
KC_NAND4_X1 D9190 ( .Y(D9190_Y), .D(D9184_Y), .C(D9188_Y), .B(D9189_Y),     .A(D1996_Y));
KC_NAND4_X1 D9178 ( .Y(D9178_Y), .D(D9173_Y), .C(D9185_Y), .B(D9177_Y),     .A(D9232_Y));
KC_NAND4_X1 D9171 ( .Y(D9171_Y), .D(D9170_Y), .C(D9169_Y), .B(D9233_Y),     .A(D1999_Y));
KC_NAND4_X1 D9119 ( .Y(D9119_Y), .D(D9120_Y), .C(D7635_Y), .B(D9121_Y),     .A(D9121_Y));
KC_NAND4_X1 D9067 ( .Y(D9067_Y), .D(D7542_Y), .C(D59_Y), .B(D26_Y),     .A(D2005_Y));
KC_NAND4_X1 D9066 ( .Y(D9066_Y), .D(D7566_Y), .C(D9062_Y), .B(D9032_Y),     .A(D8982_Y));
KC_NAND4_X1 D9050 ( .Y(D9050_Y), .D(D9095_Y), .C(D7546_Y), .B(D9044_Y),     .A(D8961_Y));
KC_NAND4_X1 D9040 ( .Y(D9040_Y), .D(D2045_Y), .C(D7551_Y), .B(D9092_Y),     .A(D9036_Y));
KC_NAND4_X1 D8978 ( .Y(D8978_Y), .D(D9010_Y), .C(D9011_Y), .B(D9091_Y),     .A(D9009_Y));
KC_NAND4_X1 D8977 ( .Y(D8977_Y), .D(D9145_Y), .C(D2077_Y), .B(D9007_Y),     .A(D320_Y));
KC_NAND4_X1 D8975 ( .Y(D8975_Y), .D(D9004_Y), .C(D7528_Y), .B(D7525_Y),     .A(D9008_Y));
KC_NAND4_X1 D8962 ( .Y(D8962_Y), .D(D7491_Y), .C(D8963_Y), .B(D2010_Y),     .A(D8960_Y));
KC_NAND4_X1 D8922 ( .Y(D8922_Y), .D(D8848_Y), .C(D8916_Y), .B(D8925_Y),     .A(D8920_Y));
KC_NAND4_X1 D8915 ( .Y(D8915_Y), .D(D8912_Y), .C(D8913_Y), .B(D8924_Y),     .A(D8921_Y));
KC_NAND4_X1 D8875 ( .Y(D8875_Y), .D(D8871_Y), .C(D8872_Y), .B(D8873_Y),     .A(D8923_Y));
KC_NAND4_X1 D8868 ( .Y(D8868_Y), .D(D8870_Y), .C(D8863_Y), .B(D8867_Y),     .A(D8914_Y));
KC_NAND4_X1 D8862 ( .Y(D8862_Y), .D(D8927_Y), .C(D8850_Y), .B(D8856_Y),     .A(D8858_Y));
KC_NAND4_X1 D8761 ( .Y(D8761_Y), .D(D9981_Q), .C(D9980_Q), .B(D233_Q),     .A(D8823_Q));
KC_NAND4_X1 D8754 ( .Y(D8754_Y), .D(D8741_Y), .C(D8743_Y), .B(D2095_Y),     .A(D9480_Y));
KC_NAND4_X1 D8753 ( .Y(D8753_Y), .D(D8757_Y), .C(D8801_Y), .B(D8789_Y),     .A(D8793_Y));
KC_NAND4_X1 D8752 ( .Y(D8752_Y), .D(D2027_Y), .C(D7183_Y), .B(D2095_Y),     .A(D8747_Y));
KC_NAND4_X1 D8679 ( .Y(D8679_Y), .D(D8710_Y), .C(D188_Y), .B(D8683_Y),     .A(D188_Y));
KC_NAND4_X1 D8670 ( .Y(D8670_Y), .D(D8725_Y), .C(D8731_Y), .B(D8673_Y),     .A(D8723_Y));
KC_NAND4_X1 D8664 ( .Y(D8664_Y), .D(D227_Q), .C(D9950_Q), .B(D9941_Q),     .A(D8712_Q));
KC_NAND4_X1 D8610 ( .Y(D8610_Y), .D(D7086_Y), .C(D8617_Y), .B(D8647_Y),     .A(D7023_Y));
KC_NAND4_X1 D8609 ( .Y(D8609_Y), .D(D7091_Y), .C(D8612_Y), .B(D8646_Y),     .A(D7073_Y));
KC_NAND4_X1 D8417 ( .Y(D8417_Y), .D(D8200_Y), .C(D2267_Y), .B(D8416_Y),     .A(D8556_Y));
KC_NAND4_X1 D8409 ( .Y(D8409_Y), .D(D8075_Y), .C(D2266_Y), .B(D8407_Y),     .A(D8624_Y));
KC_NAND4_X1 D8399 ( .Y(D8399_Y), .D(D8096_Y), .C(D80_Y), .B(D8396_Y),     .A(D8554_Y));
KC_NAND4_X1 D8398 ( .Y(D8398_Y), .D(D8103_Y), .C(D2313_Y), .B(D8408_Y),     .A(D8625_Y));
KC_NAND4_X1 D8391 ( .Y(D8391_Y), .D(D8097_Y), .C(D12424_Y),     .B(D8373_Y), .A(D8555_Y));
KC_NAND4_X1 D8390 ( .Y(D8390_Y), .D(D8104_Y), .C(D12425_Y),     .B(D8389_Y), .A(D8621_Y));
KC_NAND4_X1 D8380 ( .Y(D8380_Y), .D(D8112_Y), .C(D12429_Y),     .B(D8379_Y), .A(D8553_Y));
KC_NAND4_X1 D8375 ( .Y(D8375_Y), .D(D8074_Y), .C(D2318_Y), .B(D8374_Y),     .A(D8613_Y));
KC_NAND4_X1 D8277 ( .Y(D8277_Y), .D(D8334_Y), .C(D11818_Y),     .B(D10843_Y), .A(D5334_Y));
KC_NAND4_X1 D8275 ( .Y(D8275_Y), .D(D8118_Y), .C(D12373_Y),     .B(D8271_Y), .A(D8615_Y));
KC_NAND4_X1 D8274 ( .Y(D8274_Y), .D(D8113_Y), .C(D864_Y), .B(D8347_Y),     .A(D8619_Y));
KC_NAND4_X1 D8273 ( .Y(D8273_Y), .D(D8335_Y), .C(D11816_Y),     .B(D10842_Y), .A(D5333_Y));
KC_NAND4_X1 D8272 ( .Y(D8272_Y), .D(D8333_Y), .C(D11817_Y),     .B(D2195_Y), .A(D5332_Y));
KC_NAND4_X1 D8270 ( .Y(D8270_Y), .D(D8332_Y), .C(D11832_Y),     .B(D10838_Y), .A(D859_Y));
KC_NAND4_X1 D8269 ( .Y(D8269_Y), .D(D8188_Y), .C(D12372_Y),     .B(D8268_Y), .A(D1829_Y));
KC_NAND4_X1 D8183 ( .Y(D8183_Y), .D(D8190_Y), .C(D8256_Y), .B(D8190_Y),     .A(D8219_Y));
KC_NAND4_X1 D8174 ( .Y(D8174_Y), .D(D1944_Q), .C(D8243_Q), .B(D8245_Q),     .A(D8244_Q));
KC_NAND4_X1 D8116 ( .Y(D8116_Y), .D(D8115_Y), .C(D8220_Y), .B(D1984_Y),     .A(D8221_Y));
KC_NAND4_X1 D7844 ( .Y(D7844_Y), .D(D7901_Y), .C(D7843_Y), .B(D7945_Y),     .A(D7875_Y));
KC_NAND4_X1 D7826 ( .Y(D7826_Y), .D(D7831_Y), .C(D7840_Y), .B(D1854_Y),     .A(D1917_Y));
KC_NAND4_X1 D7768 ( .Y(D7768_Y), .D(D9320_Y), .C(D12863_Y),     .B(D13288_Y), .A(D724_Y));
KC_NAND4_X1 D7765 ( .Y(D7765_Y), .D(D13171_Y), .C(D13289_Y),     .B(D13280_Q), .A(D13287_Y));
KC_NAND4_X1 D7764 ( .Y(D7764_Y), .D(D10155_Y), .C(D12762_Y),     .B(D12301_Y), .A(D725_Y));
KC_NAND4_X1 D7760 ( .Y(D7760_Y), .D(D12300_Y), .C(D12763_Y),     .B(D12761_Y), .A(D12764_Y));
KC_NAND4_X1 D7688 ( .Y(D7688_Y), .D(D7729_Y), .C(D7755_Y), .B(D7724_Y),     .A(D7725_Y));
KC_NAND4_X1 D7685 ( .Y(D7685_Y), .D(D7720_Y), .C(D7722_Y), .B(D7650_Y),     .A(D7726_Y));
KC_NAND4_X1 D7679 ( .Y(D7679_Y), .D(D10160_Y), .C(D12300_Y),     .B(D13287_Y), .A(D12762_Y));
KC_NAND4_X1 D7676 ( .Y(D7676_Y), .D(D7785_Y), .C(D9354_Y),     .B(D12761_Y), .A(D724_Y));
KC_NAND4_X1 D7675 ( .Y(D7675_Y), .D(D7717_Y), .C(D7714_Y), .B(D7715_Y),     .A(D7716_Y));
KC_NAND4_X1 D7673 ( .Y(D7673_Y), .D(D7735_Q), .C(D7734_Q), .B(D7736_Q),     .A(D7745_Q));
KC_NAND4_X1 D7622 ( .Y(D7622_Y), .D(D7689_Y), .C(D7677_Y),     .B(D13280_Q), .A(D280_Y));
KC_NAND4_X1 D7541 ( .Y(D7541_Y), .D(D7639_Y), .C(D1938_Y), .B(D7628_Y),     .A(D7572_Y));
KC_NAND4_X1 D7489 ( .Y(D7489_Y), .D(D6637_Y), .C(D1767_Y), .B(D1769_Y),     .A(D6157_Y));
KC_NAND4_X1 D7437 ( .Y(D7437_Y), .D(D1880_Y), .C(D5867_Y), .B(D7337_Y),     .A(D7480_Q));
KC_NAND4_X1 D7433 ( .Y(D7433_Y), .D(D5705_Y), .C(D7419_Y), .B(D287_Y),     .A(D6003_Y));
KC_NAND4_X1 D7432 ( .Y(D7432_Y), .D(D7444_Y), .C(D306_Y), .B(D8849_Y),     .A(D8965_Y));
KC_NAND4_X1 D7425 ( .Y(D7425_Y), .D(D7472_Y), .C(D7377_Y), .B(D7733_Q),     .A(D7446_Y));
KC_NAND4_X1 D7416 ( .Y(D7416_Y), .D(D6041_Y), .C(D5966_Y), .B(D5646_Y),     .A(D726_Y));
KC_NAND4_X1 D7355 ( .Y(D7355_Y), .D(D179_Y), .C(D5703_Y), .B(D5647_Y),     .A(D1736_Y));
KC_NAND4_X1 D7321 ( .Y(D7321_Y), .D(D5704_Y), .C(D7322_Y), .B(D7375_Y),     .A(D7314_Y));
KC_NAND4_X1 D7253 ( .Y(D7253_Y), .D(D7260_Y), .C(D7101_Y), .B(D7140_Y),     .A(D6333_Y));
KC_NAND4_X1 D7252 ( .Y(D7252_Y), .D(D7092_Y), .C(D6334_Y), .B(D6333_Y),     .A(D7141_Y));
KC_NAND4_X1 D7231 ( .Y(D7231_Y), .D(D8778_Y), .C(D9475_Y), .B(D7170_Y),     .A(D8760_Y));
KC_NAND4_X1 D7228 ( .Y(D7228_Y), .D(D7183_Y), .C(D8876_Y), .B(D9477_Y),     .A(D9480_Y));
KC_NAND4_X1 D7227 ( .Y(D7227_Y), .D(D8756_Y), .C(D8749_Y), .B(D8743_Y),     .A(D9477_Y));
KC_NAND4_X1 D7215 ( .Y(D7215_Y), .D(D1887_Y), .C(D7217_Y), .B(D8749_Y),     .A(D8812_Y));
KC_NAND4_X1 D7208 ( .Y(D7208_Y), .D(D202_Y), .C(D7215_Y), .B(D7216_Y),     .A(D7202_Y));
KC_NAND4_X1 D7201 ( .Y(D7201_Y), .D(D209_Y), .C(D9475_Y), .B(D2026_Y),     .A(D9476_Y));
KC_NAND4_X1 D7191 ( .Y(D7191_Y), .D(D7196_Y), .C(D7354_Y), .B(D7341_Y),     .A(D7310_Y));
KC_NAND4_X1 D7190 ( .Y(D7190_Y), .D(D7299_Y), .C(D5748_Y), .B(D1882_Y),     .A(D1725_Y));
KC_NAND4_X1 D7189 ( .Y(D7189_Y), .D(D7227_Y), .C(D7205_Y), .B(D9475_Y),     .A(D7222_Y));
KC_NAND4_X1 D7174 ( .Y(D7174_Y), .D(D202_Y), .C(D7227_Y), .B(D7176_Y),     .A(D211_Y));
KC_NAND4_X1 D7173 ( .Y(D7173_Y), .D(D7175_Y), .C(D7216_Y), .B(D7238_Y),     .A(D8788_Y));
KC_NAND4_X1 D7102 ( .Y(D7102_Y), .D(D7095_Y), .C(D7235_Y), .B(D7259_Y),     .A(D7105_Y));
KC_NAND4_X1 D7074 ( .Y(D7074_Y), .D(D7090_Y), .C(D8611_Y), .B(D8644_Y),     .A(D7065_Y));
KC_NAND4_X1 D7068 ( .Y(D7068_Y), .D(D7088_Y), .C(D8616_Y), .B(D8645_Y),     .A(D7066_Y));
KC_NAND4_X1 D7039 ( .Y(D7039_Y), .D(D7059_Y), .C(D7037_Y), .B(D7038_Y),     .A(D7031_Y));
KC_NAND4_X1 D7032 ( .Y(D7032_Y), .D(D7060_Y), .C(D7040_Y), .B(D7036_Y),     .A(D7034_Y));
KC_NAND4_X1 D7027 ( .Y(D7027_Y), .D(D7058_Y), .C(D7033_Y), .B(D7028_Y),     .A(D7067_Y));
KC_NAND4_X1 D7026 ( .Y(D7026_Y), .D(D7057_Y), .C(D7030_Y), .B(D7025_Y),     .A(D7070_Y));
KC_NAND4_X1 D7022 ( .Y(D7022_Y), .D(D7087_Y), .C(D8620_Y), .B(D8648_Y),     .A(D7020_Y));
KC_NAND4_X1 D7021 ( .Y(D7021_Y), .D(D7089_Y), .C(D1254_Y), .B(D7071_Y),     .A(D7072_Y));
KC_NAND4_X1 D6985 ( .Y(D6985_Y), .D(D1318_Y), .C(D6983_Y), .B(D62_Y),     .A(D1167_Y));
KC_NAND4_X1 D6981 ( .Y(D6981_Y), .D(D1319_Y), .C(D6979_Y), .B(D6980_Y),     .A(D6984_Y));
KC_NAND4_X1 D6918 ( .Y(D6918_Y), .D(D5535_Y), .C(D6988_Y), .B(D1080_Y),     .A(D5511_Y));
KC_NAND4_X1 D6872 ( .Y(D6872_Y), .D(D1789_Y), .C(D6865_Y), .B(D6834_Y),     .A(D5425_Y));
KC_NAND4_X1 D6871 ( .Y(D6871_Y), .D(D6906_Y), .C(D6849_Y), .B(D6846_Y),     .A(D6844_Y));
KC_NAND4_X1 D6867 ( .Y(D6867_Y), .D(D1788_Y), .C(D6850_Y), .B(D6841_Y),     .A(D6837_Y));
KC_NAND4_X1 D6866 ( .Y(D6866_Y), .D(D6905_Y), .C(D6852_Y), .B(D6835_Y),     .A(D6838_Y));
KC_NAND4_X1 D6859 ( .Y(D6859_Y), .D(D6907_Y), .C(D6851_Y), .B(D6845_Y),     .A(D971_Y));
KC_NAND4_X1 D6848 ( .Y(D6848_Y), .D(D6908_Y), .C(D6857_Y), .B(D6839_Y),     .A(D5424_Y));
KC_NAND4_X1 D6847 ( .Y(D6847_Y), .D(D6904_Y), .C(D6858_Y), .B(D6840_Y),     .A(D969_Y));
KC_NAND4_X1 D6725 ( .Y(D6725_Y), .D(D5330_Y), .C(D6724_Y), .B(D6723_Y),     .A(D6721_Y));
KC_NAND4_X1 D6717 ( .Y(D6717_Y), .D(D5329_Y), .C(D6722_Y), .B(D6715_Y),     .A(D6716_Y));
KC_NAND4_X1 D6709 ( .Y(D6709_Y), .D(D5328_Y), .C(D6704_Y), .B(D6712_Y),     .A(D6708_Y));
KC_NAND4_X1 D6707 ( .Y(D6707_Y), .D(D5327_Y), .C(D6705_Y), .B(D6714_Y),     .A(D6703_Y));
KC_NAND4_X1 D6698 ( .Y(D6698_Y), .D(D5326_Y), .C(D6701_Y), .B(D6690_Y),     .A(D6697_Y));
KC_NAND4_X1 D6694 ( .Y(D6694_Y), .D(D5325_Y), .C(D6700_Y), .B(D6683_Y),     .A(D6686_Y));
KC_NAND4_X1 D6693 ( .Y(D6693_Y), .D(D5324_Y), .C(D6696_Y), .B(D6687_Y),     .A(D6692_Y));
KC_NAND4_X1 D6688 ( .Y(D6688_Y), .D(D811_Y), .C(D6691_Y), .B(D6684_Y),     .A(D6685_Y));
KC_NAND4_X1 D6634 ( .Y(D6634_Y), .D(D5241_Y), .C(D6641_Y), .B(D1691_Y),     .A(D6628_Y));
KC_NAND4_X1 D6633 ( .Y(D6633_Y), .D(D5242_Y), .C(D6638_Y), .B(D6626_Y),     .A(D6630_Y));
KC_NAND4_X1 D6625 ( .Y(D6625_Y), .D(D5245_Y), .C(D6632_Y), .B(D6629_Y),     .A(D6623_Y));
KC_NAND4_X1 D6624 ( .Y(D6624_Y), .D(D5244_Y), .C(D6631_Y), .B(D6627_Y),     .A(D6622_Y));
KC_NAND4_X1 D6619 ( .Y(D6619_Y), .D(D5254_Y), .C(D6620_Y), .B(D6635_Y),     .A(D5202_Y));
KC_NAND4_X1 D6618 ( .Y(D6618_Y), .D(D5243_Y), .C(D6621_Y), .B(D6636_Y),     .A(D623_Y));
KC_NAND4_X1 D6589 ( .Y(D6589_Y), .D(D3698_Y), .C(D6581_Y), .B(D6587_Y),     .A(D6588_Y));
KC_NAND4_X1 D6585 ( .Y(D6585_Y), .D(D3693_Y), .C(D6572_Y), .B(D6583_Y),     .A(D6569_Y));
KC_NAND4_X1 D6584 ( .Y(D6584_Y), .D(D3694_Y), .C(D6582_Y), .B(D6590_Y),     .A(D551_Y));
KC_NAND4_X1 D6580 ( .Y(D6580_Y), .D(D3749_Y), .C(D6579_Y), .B(D6573_Y),     .A(D6577_Y));
KC_NAND4_X1 D6576 ( .Y(D6576_Y), .D(D1511_Y), .C(D6574_Y), .B(D6575_Y),     .A(D6578_Y));
KC_NAND4_X1 D6570 ( .Y(D6570_Y), .D(D3692_Y), .C(D6571_Y), .B(D6568_Y),     .A(D549_Y));
KC_NAND4_X1 D6290 ( .Y(D6290_Y), .D(D6339_Y), .C(D6319_Y), .B(D6320_Y),     .A(D6176_Y));
KC_NAND4_X1 D6215 ( .Y(D6215_Y), .D(D6217_Y), .C(D7731_Y), .B(D7701_Y),     .A(D7649_Y));
KC_NAND4_X1 D6138 ( .Y(D6138_Y), .D(D6181_Y), .C(D6155_Y), .B(D5930_Y),     .A(D6159_Y));
KC_NAND4_X1 D6132 ( .Y(D6132_Y), .D(D6178_Y), .C(D6180_Y), .B(D7784_Y),     .A(D6179_Y));
KC_NAND4_X1 D6085 ( .Y(D6085_Y), .D(D6637_Y), .C(D1767_Y), .B(D1769_Y),     .A(D6637_Y));
KC_NAND4_X1 D6084 ( .Y(D6084_Y), .D(D6102_Y), .C(D6101_Y), .B(D6165_Y),     .A(D322_Y));
KC_NAND4_X1 D6031 ( .Y(D6031_Y), .D(D253_Y), .C(D7321_Y), .B(D6082_Y),     .A(D7337_Y));
KC_NAND4_X1 D6030 ( .Y(D6030_Y), .D(D6025_Y), .C(D6013_Y), .B(D5841_Y),     .A(D5646_Y));
KC_NAND4_X1 D6029 ( .Y(D6029_Y), .D(D6047_Y), .C(D6069_Y), .B(D6034_Y),     .A(D5979_Y));
KC_NAND4_X1 D6017 ( .Y(D6017_Y), .D(D6002_Y), .C(D5641_Y), .B(D6049_Y),     .A(D6022_Y));
KC_NAND4_X1 D6016 ( .Y(D6016_Y), .D(D1581_Y), .C(D5954_Y), .B(D6077_Y),     .A(D4427_Y));
KC_NAND4_X1 D6005 ( .Y(D6005_Y), .D(D6012_Y), .C(D1713_Y), .B(D5954_Y),     .A(D7164_Y));
KC_NAND4_X1 D5999 ( .Y(D5999_Y), .D(D1713_Y), .C(D4416_Y), .B(D4408_Y),     .A(D235_Y));
KC_NAND4_X1 D5998 ( .Y(D5998_Y), .D(D8944_Y), .C(D229_Q), .B(D5693_Q),     .A(D4136_Q));
KC_NAND4_X1 D5997 ( .Y(D5997_Y), .D(D4421_Y), .C(D4417_Y), .B(D4235_Q),     .A(D4150_Y));
KC_NAND4_X1 D5996 ( .Y(D5996_Y), .D(D4431_Y), .C(D6000_Y), .B(D5962_Y),     .A(D5869_Y));
KC_NAND4_X1 D5995 ( .Y(D5995_Y), .D(D6065_Y), .C(D5869_Y), .B(D1708_Y),     .A(D5671_Y));
KC_NAND4_X1 D5991 ( .Y(D5991_Y), .D(D5967_Y), .C(D7984_Y), .B(D5877_Y),     .A(D6007_Y));
KC_NAND4_X1 D5961 ( .Y(D5961_Y), .D(D4294_Y), .C(D4412_Y), .B(D275_Y),     .A(D165_Y));
KC_NAND4_X1 D5951 ( .Y(D5951_Y), .D(D5792_Y), .C(D12305_Y),     .B(D6062_Y), .A(D275_Y));
KC_NAND4_X1 D5950 ( .Y(D5950_Y), .D(D4417_Y), .C(D7499_Y), .B(D5953_Y),     .A(D239_Q));
KC_NAND4_X1 D5892 ( .Y(D5892_Y), .D(D5885_Y), .C(D1736_Y), .B(D251_Y),     .A(D5916_Y));
KC_NAND4_X1 D5862 ( .Y(D5862_Y), .D(D7321_Y), .C(D7203_Y), .B(D1738_Y),     .A(D5860_Y));
KC_NAND4_X1 D5861 ( .Y(D5861_Y), .D(D5923_Y), .C(D5826_Y), .B(D5878_Y),     .A(D5860_Y));
KC_NAND4_X1 D5855 ( .Y(D5855_Y), .D(D7321_Y), .C(D7303_Y), .B(D1739_Y),     .A(D287_Y));
KC_NAND4_X1 D5854 ( .Y(D5854_Y), .D(D5844_Y), .C(D7339_Y), .B(D5843_Y),     .A(D5842_Y));
KC_NAND4_X1 D5853 ( .Y(D5853_Y), .D(D5926_Y), .C(D7100_Y), .B(D5710_Y),     .A(D7337_Y));
KC_NAND4_X1 D5845 ( .Y(D5845_Y), .D(D5920_Y), .C(D5893_Y), .B(D5943_Y),     .A(D7374_Y));
KC_NAND4_X1 D5750 ( .Y(D5750_Y), .D(D7286_Y), .C(D5797_Y), .B(D4321_Y),     .A(D5740_Y));
KC_NAND4_X1 D5735 ( .Y(D5735_Y), .D(D7211_Y), .C(D269_Y), .B(D5732_Y),     .A(D1725_Y));
KC_NAND4_X1 D5731 ( .Y(D5731_Y), .D(D7203_Y), .C(D4198_Y), .B(D5767_Y),     .A(D5817_Y));
KC_NAND4_X1 D5725 ( .Y(D5725_Y), .D(D5840_Y), .C(D7184_Y), .B(D4136_Q),     .A(D5693_Q));
KC_NAND4_X1 D5724 ( .Y(D5724_Y), .D(D7185_Y), .C(D5840_Y), .B(D5649_Y),     .A(D4226_Y));
KC_NAND4_X1 D5720 ( .Y(D5720_Y), .D(D5995_Y), .C(D5723_Y), .B(D5757_Y),     .A(D5764_Y));
KC_NAND4_X1 D5719 ( .Y(D5719_Y), .D(D4249_Y), .C(D5656_Y), .B(D5727_Y),     .A(D5718_Y));
KC_NAND4_X1 D5710 ( .Y(D5710_Y), .D(D4226_Y), .C(D1956_Y), .B(D7184_Y),     .A(D4119_Q));
KC_NAND4_X1 D5659 ( .Y(D5659_Y), .D(D5664_Y), .C(D5686_Q), .B(D5690_Q),     .A(D5691_Q));
KC_NAND4_X1 D5641 ( .Y(D5641_Y), .D(D5642_Y), .C(D7255_Y), .B(D7093_Y),     .A(D7256_Y));
KC_NAND4_X1 D5623 ( .Y(D5623_Y), .D(D5635_Y), .C(D5585_Y), .B(D5575_Y),     .A(D5619_Y));
KC_NAND4_X1 D5600 ( .Y(D5600_Y), .D(D5612_Y), .C(D5602_Y), .B(D5597_Y),     .A(D1541_Y));
KC_NAND4_X1 D5599 ( .Y(D5599_Y), .D(D5614_Y), .C(D5601_Y), .B(D5596_Y),     .A(D1542_Y));
KC_NAND4_X1 D5587 ( .Y(D5587_Y), .D(D5638_Y), .C(D5593_Y), .B(D5586_Y),     .A(D5580_Y));
KC_NAND4_X1 D5584 ( .Y(D5584_Y), .D(D5639_Y), .C(D5592_Y), .B(D5583_Y),     .A(D5615_Y));
KC_NAND4_X1 D5582 ( .Y(D5582_Y), .D(D5636_Y), .C(D5590_Y), .B(D5581_Y),     .A(D5621_Y));
KC_NAND4_X1 D5579 ( .Y(D5579_Y), .D(D5637_Y), .C(D5589_Y), .B(D5576_Y),     .A(D5622_Y));
KC_NAND4_X1 D5578 ( .Y(D5578_Y), .D(D5634_Y), .C(D5588_Y), .B(D5577_Y),     .A(D5618_Y));
KC_NAND4_X1 D5547 ( .Y(D5547_Y), .D(D5613_Y), .C(D5572_Y), .B(D1539_Y),     .A(D5545_Y));
KC_NAND4_X1 D5546 ( .Y(D5546_Y), .D(D5611_Y), .C(D5544_Y), .B(D1540_Y),     .A(D5548_Y));
KC_NAND4_X1 D5508 ( .Y(D5508_Y), .D(D5539_Y), .C(D1170_Y), .B(D5493_Y),     .A(D5512_Y));
KC_NAND4_X1 D5507 ( .Y(D5507_Y), .D(D5537_Y), .C(D5549_Y), .B(D1548_Y),     .A(D5514_Y));
KC_NAND4_X1 D5502 ( .Y(D5502_Y), .D(D5536_Y), .C(D5554_Y), .B(D1547_Y),     .A(D5515_Y));
KC_NAND4_X1 D5501 ( .Y(D5501_Y), .D(D5538_Y), .C(D5553_Y), .B(D1545_Y),     .A(D5513_Y));
KC_NAND4_X1 D5496 ( .Y(D5496_Y), .D(D1649_Y), .C(D5550_Y), .B(D1546_Y),     .A(D5499_Y));
KC_NAND4_X1 D5495 ( .Y(D5495_Y), .D(D5541_Y), .C(D5552_Y), .B(D1543_Y),     .A(D5516_Y));
KC_NAND4_X1 D5494 ( .Y(D5494_Y), .D(D1650_Y), .C(D5551_Y), .B(D1544_Y),     .A(D5506_Y));
KC_NAND4_X1 D5446 ( .Y(D5446_Y), .D(D3947_Y), .C(D5443_Y), .B(D3922_Y),     .A(D5444_Y));
KC_NAND4_X1 D5435 ( .Y(D5435_Y), .D(D3979_Y), .C(D5433_Y), .B(D5423_Y),     .A(D5421_Y));
KC_NAND4_X1 D5430 ( .Y(D5430_Y), .D(D3976_Y), .C(D5439_Y), .B(D63_Y),     .A(D1549_Y));
KC_NAND4_X1 D5429 ( .Y(D5429_Y), .D(D1510_Y), .C(D5434_Y), .B(D3895_Y),     .A(D5428_Y));
KC_NAND4_X1 D5420 ( .Y(D5420_Y), .D(D1507_Y), .C(D5438_Y), .B(D3893_Y),     .A(D5422_Y));
KC_NAND4_X1 D5418 ( .Y(D5418_Y), .D(D3882_Y), .C(D5337_Y), .B(D5335_Y),     .A(D5343_Y));
KC_NAND4_X1 D5366 ( .Y(D5366_Y), .D(D3884_Y), .C(D5367_Y), .B(D5351_Y),     .A(D5362_Y));
KC_NAND4_X1 D5365 ( .Y(D5365_Y), .D(D3885_Y), .C(D5364_Y), .B(D5352_Y),     .A(D5363_Y));
KC_NAND4_X1 D5339 ( .Y(D5339_Y), .D(D3883_Y), .C(D5336_Y), .B(D3831_Y),     .A(D5338_Y));
KC_NAND4_X1 D5293 ( .Y(D5293_Y), .D(D3745_Y), .C(D5290_Y), .B(D5279_Y),     .A(D5289_Y));
KC_NAND4_X1 D5288 ( .Y(D5288_Y), .D(D3748_Y), .C(D5285_Y), .B(D5271_Y),     .A(D5283_Y));
KC_NAND4_X1 D5277 ( .Y(D5277_Y), .D(D3747_Y), .C(D5275_Y), .B(D5272_Y),     .A(D5292_Y));
KC_NAND4_X1 D5276 ( .Y(D5276_Y), .D(D3828_Y), .C(D5286_Y), .B(D5274_Y),     .A(D5280_Y));
KC_NAND4_X1 D5268 ( .Y(D5268_Y), .D(D3823_Y), .C(D5257_Y), .B(D5269_Y),     .A(D5263_Y));
KC_NAND4_X1 D5258 ( .Y(D5258_Y), .D(D3820_Y), .C(D5255_Y), .B(D5264_Y),     .A(D5256_Y));
KC_NAND4_X1 D5213 ( .Y(D5213_Y), .D(D5246_Y), .C(D6639_Y), .B(D5206_Y),     .A(D5207_Y));
KC_NAND4_X1 D5180 ( .Y(D5180_Y), .D(D3699_Y), .C(D5175_Y), .B(D5177_Y),     .A(D5169_Y));
KC_NAND4_X1 D5174 ( .Y(D5174_Y), .D(D3697_Y), .C(D5167_Y), .B(D5178_Y),     .A(D5163_Y));
KC_NAND4_X1 D5173 ( .Y(D5173_Y), .D(D3695_Y), .C(D5170_Y), .B(D5144_Y),     .A(D5164_Y));
KC_NAND4_X1 D5172 ( .Y(D5172_Y), .D(D3696_Y), .C(D5161_Y), .B(D5176_Y),     .A(D6586_Y));
KC_NAND4_X1 D5171 ( .Y(D5171_Y), .D(D600_Y), .C(D5162_Y), .B(D5179_Y),     .A(D550_Y));
KC_NAND4_X1 D5166 ( .Y(D5166_Y), .D(D3689_Y), .C(D5168_Y), .B(D5143_Y),     .A(D5165_Y));
KC_NAND4_X1 D5160 ( .Y(D5160_Y), .D(D3690_Y), .C(D5156_Y), .B(D5152_Y),     .A(D5147_Y));
KC_NAND4_X1 D5159 ( .Y(D5159_Y), .D(D3691_Y), .C(D5151_Y), .B(D5149_Y),     .A(D5199_Y));
KC_NAND4_X1 D5155 ( .Y(D5155_Y), .D(D3687_Y), .C(D5153_Y), .B(D5150_Y),     .A(D5145_Y));
KC_NAND4_X1 D5154 ( .Y(D5154_Y), .D(D3688_Y), .C(D5158_Y), .B(D5157_Y),     .A(D5146_Y));
KC_NAND4_X1 D5017 ( .Y(D5017_Y), .D(D5014_Y), .C(D5092_Y), .B(D5026_Y),     .A(D5013_Y));
KC_NAND4_X1 D5016 ( .Y(D5016_Y), .D(D5058_Y), .C(D5018_Y), .B(D4912_Y),     .A(D5013_Y));
KC_NAND4_X1 D4994 ( .Y(D4994_Y), .D(D4998_Y), .C(D5082_Y), .B(D5015_Y),     .A(D5073_Y));
KC_NAND4_X1 D4993 ( .Y(D4993_Y), .D(D488_Y), .C(D5057_Y), .B(D3513_Y),     .A(D1560_Y));
KC_NAND4_X1 D4990 ( .Y(D4990_Y), .D(D4991_Y), .C(D5027_Y), .B(D4986_Y),     .A(D5070_Y));
KC_NAND4_X1 D4989 ( .Y(D4989_Y), .D(D5000_Y), .C(D5045_Y), .B(D4988_Y),     .A(D470_Y));
KC_NAND4_X1 D4984 ( .Y(D4984_Y), .D(D5045_Y), .C(D5079_Y), .B(D5093_Y),     .A(D5084_Y));
KC_NAND4_X1 D4890 ( .Y(D4890_Y), .D(D4933_Y), .C(D4896_Y), .B(D4880_Y),     .A(D4902_Y));
KC_NAND4_X1 D4864 ( .Y(D4864_Y), .D(D4928_Y), .C(D4932_Y), .B(D4870_Y),     .A(D3523_Y));
KC_NAND4_X1 D4863 ( .Y(D4863_Y), .D(D3470_Y), .C(D4930_Y), .B(D1446_Y),     .A(D4907_Y));
KC_NAND4_X1 D4773 ( .Y(D4773_Y), .D(D4818_Q), .C(D4820_Q), .B(D4821_Q),     .A(D4822_Q));
KC_NAND4_X1 D4765 ( .Y(D4765_Y), .D(D4811_Y), .C(D4820_Q), .B(D4821_Q),     .A(D4822_Q));
KC_NAND4_X1 D4689 ( .Y(D4689_Y), .D(D4575_Y), .C(D4688_Y), .B(D4578_Y),     .A(D4638_Q));
KC_NAND4_X1 D4677 ( .Y(D4677_Y), .D(D4708_Y), .C(D4707_Y), .B(D4678_Y),     .A(D4681_Y));
KC_NAND4_X1 D4676 ( .Y(D4676_Y), .D(D4686_Y), .C(D4679_Y), .B(D4732_Y),     .A(D4656_Y));
KC_NAND4_X1 D4675 ( .Y(D4675_Y), .D(D1668_Y), .C(D4660_Y), .B(D4674_Y),     .A(D3227_Y));
KC_NAND4_X1 D4662 ( .Y(D4662_Y), .D(D4617_Y), .C(D3219_Y), .B(D4658_Y),     .A(D4657_Y));
KC_NAND4_X1 D4496 ( .Y(D4496_Y), .D(D4505_Y), .C(D1648_Y), .B(D1578_Y),     .A(D1945_Y));
KC_NAND4_X1 D6 ( .Y(D6_Y), .D(D4387_Y), .C(D1632_Y), .B(D351_Y),     .A(D4474_Y));
KC_NAND4_X1 D4443 ( .Y(D4443_Y), .D(D4438_Y), .C(D1719_Y), .B(D239_Q),     .A(D8838_Y));
KC_NAND4_X1 D4442 ( .Y(D4442_Y), .D(D7467_Y), .C(D4472_Y), .B(D5988_Y),     .A(D6033_Y));
KC_NAND4_X1 D4437 ( .Y(D4437_Y), .D(D4440_Y), .C(D4412_Y), .B(D4427_Y),     .A(D239_Q));
KC_NAND4_X1 D4430 ( .Y(D4430_Y), .D(D5988_Y), .C(D5989_Y), .B(D4235_Q),     .A(D228_Q));
KC_NAND4_X1 D4429 ( .Y(D4429_Y), .D(D4471_Y), .C(D4473_Y), .B(D4475_Y),     .A(D4469_Y));
KC_NAND4_X1 D4353 ( .Y(D4353_Y), .D(D4360_Y), .C(D1592_Y), .B(D4332_Y),     .A(D4346_Y));
KC_NAND4_X1 D4333 ( .Y(D4333_Y), .D(D4329_Y), .C(D4374_Y), .B(D4336_Y),     .A(D4332_Y));
KC_NAND4_X1 D4322 ( .Y(D4322_Y), .D(D4339_Y), .C(D4328_Y), .B(D4338_Y),     .A(D4277_Y));
KC_NAND4_X1 D4307 ( .Y(D4307_Y), .D(D2829_Y), .C(D4399_Y), .B(D2831_Y),     .A(D4115_Y));
KC_NAND4_X1 D4298 ( .Y(D4298_Y), .D(D4294_Y), .C(D4421_Y), .B(D165_Y),     .A(D4150_Y));
KC_NAND4_X1 D4275 ( .Y(D4275_Y), .D(D4363_Y), .C(D5977_Y), .B(D6011_Y),     .A(D4179_Y));
KC_NAND4_X1 D4274 ( .Y(D4274_Y), .D(D4309_Y), .C(D7324_Y), .B(D4284_Y),     .A(D4304_Y));
KC_NAND4_X1 D4207 ( .Y(D4207_Y), .D(D4203_Y), .C(D5733_Y), .B(D4183_Y),     .A(D4210_Y));
KC_NAND4_X1 D4177 ( .Y(D4177_Y), .D(D4228_Y), .C(D4227_Y), .B(D203_Y),     .A(D4093_Y));
KC_NAND4_X1 D4170 ( .Y(D4170_Y), .D(D4337_Y), .C(D4362_Y), .B(D5708_Y),     .A(D4176_Y));
KC_NAND4_X1 D4169 ( .Y(D4169_Y), .D(D4162_Y), .C(D4355_Y), .B(D4401_Y),     .A(D4344_Y));
KC_NAND4_X1 D4101 ( .Y(D4101_Y), .D(D4110_Y), .C(D4123_Y), .B(D4109_Y),     .A(D4225_Y));
KC_NAND4_X1 D3924 ( .Y(D3924_Y), .D(D3950_Y), .C(D3908_Y), .B(D3918_Y),     .A(D1410_Y));
KC_NAND4_X1 D3923 ( .Y(D3923_Y), .D(D3949_Y), .C(D3951_Y), .B(D3921_Y),     .A(D3917_Y));
KC_NAND4_X1 D3916 ( .Y(D3916_Y), .D(D1508_Y), .C(D3901_Y), .B(D3902_Y),     .A(D3911_Y));
KC_NAND4_X1 D3915 ( .Y(D3915_Y), .D(D1509_Y), .C(D3907_Y), .B(D3912_Y),     .A(D3910_Y));
KC_NAND4_X1 D3906 ( .Y(D3906_Y), .D(D3946_Y), .C(D3904_Y), .B(D3897_Y),     .A(D3900_Y));
KC_NAND4_X1 D3903 ( .Y(D3903_Y), .D(D3945_Y), .C(D3905_Y), .B(D3898_Y),     .A(D3896_Y));
KC_NAND4_X1 D3830 ( .Y(D3830_Y), .D(D3825_Y), .C(D3789_Y), .B(D3779_Y),     .A(D3772_Y));
KC_NAND4_X1 D3792 ( .Y(D3792_Y), .D(D3826_Y), .C(D3790_Y), .B(D3777_Y),     .A(D3773_Y));
KC_NAND4_X1 D3783 ( .Y(D3783_Y), .D(D3824_Y), .C(D3788_Y), .B(D3780_Y),     .A(D3786_Y));
KC_NAND4_X1 D3776 ( .Y(D3776_Y), .D(D3822_Y), .C(D732_Y), .B(D3770_Y),     .A(D3771_Y));
KC_NAND4_X1 D3769 ( .Y(D3769_Y), .D(D3821_Y), .C(D731_Y), .B(D3767_Y),     .A(D3765_Y));
KC_NAND4_X1 D3514 ( .Y(D3514_Y), .D(D3519_Y), .C(D3515_Y), .B(D5011_Y),     .A(D3512_Y));
KC_NAND4_X1 D3507 ( .Y(D3507_Y), .D(D3571_Y), .C(D3571_Y), .B(D3571_Y),     .A(D3545_Y));
KC_NAND4_X1 D3445 ( .Y(D3445_Y), .D(D3432_Y), .C(D4913_Y), .B(D3373_Q),     .A(D3479_Y));
KC_NAND4_X1 D3436 ( .Y(D3436_Y), .D(D4893_Y), .C(D4912_Y), .B(D3435_Y),     .A(D3412_Y));
KC_NAND4_X1 D3425 ( .Y(D3425_Y), .D(D3473_Y), .C(D3495_Y), .B(D3417_Y),     .A(D4943_Y));
KC_NAND4_X1 D3320 ( .Y(D3320_Y), .D(D3317_Y), .C(D3275_Y), .B(D3208_Y),     .A(D3369_Y));
KC_NAND4_X1 D3319 ( .Y(D3319_Y), .D(D3317_Y), .C(D3329_Y), .B(D3369_Y),     .A(D3387_Q));
KC_NAND4_X1 D3228 ( .Y(D3228_Y), .D(D3293_Y), .C(D3380_Y), .B(D3143_Y),     .A(D3348_Y));
KC_NAND4_X1 D3212 ( .Y(D3212_Y), .D(D4617_Y), .C(D4710_Y), .B(D1427_Y),     .A(D3214_Y));
KC_NAND4_X1 D3148 ( .Y(D3148_Y), .D(D1432_Y), .C(D3144_Y), .B(D3187_Q),     .A(D3188_Q));
KC_NAND4_X1 D3137 ( .Y(D3137_Y), .D(D3138_Y), .C(D3190_Q), .B(D3187_Q),     .A(D3189_Q));
KC_NAND4_X1 D3124 ( .Y(D3124_Y), .D(D3134_Y), .C(D3139_Y), .B(D1430_Y),     .A(D3189_Q));
KC_NAND4_X1 D3116 ( .Y(D3116_Y), .D(D1430_Y), .C(D3185_Q), .B(D3188_Q),     .A(D3130_Y));
KC_NAND4_X1 D3105 ( .Y(D3105_Y), .D(D1429_Y), .C(D4573_Y), .B(D3199_Y),     .A(D3126_Y));
KC_NAND4_X1 D3104 ( .Y(D3104_Y), .D(D4770_Y), .C(D3124_Y), .B(D3183_Y),     .A(D3111_Y));
KC_NAND4_X1 D3096 ( .Y(D3096_Y), .D(D3118_Y), .C(D3116_Y), .B(D3117_Y),     .A(D3126_Y));
KC_NAND4_X1 D3018 ( .Y(D3018_Y), .D(D3015_Y), .C(D3041_Y), .B(D3084_Q),     .A(D3079_Q));
KC_NAND4_X1 D3012 ( .Y(D3012_Y), .D(D3039_Y), .C(D3079_Q), .B(D1515_Q),     .A(D3080_Q));
KC_NAND4_X1 D3010 ( .Y(D3010_Y), .D(D3036_Y), .C(D3050_Y), .B(D3011_Y),     .A(D6255_Y));
KC_NAND4_X1 D2938 ( .Y(D2938_Y), .D(D2953_Y), .C(D2990_Y), .B(D2991_Y),     .A(D2982_Y));
KC_NAND4_X1 D2931 ( .Y(D2931_Y), .D(D2941_Y), .C(D2894_Y), .B(D2987_Y),     .A(D1435_Y));
KC_NAND4_X1 D2924 ( .Y(D2924_Y), .D(D2940_Y), .C(D2894_Y), .B(D2986_Y),     .A(D1435_Y));
KC_NAND4_X1 D2923 ( .Y(D2923_Y), .D(D2945_Y), .C(D2894_Y), .B(D1490_Y),     .A(D1435_Y));
KC_NAND4_X1 D2849 ( .Y(D2849_Y), .D(D2808_Y), .C(D2848_Y), .B(D1437_Y),     .A(D1441_Y));
KC_NAND4_X1 D2845 ( .Y(D2845_Y), .D(D2823_Y), .C(D2887_Q), .B(D2890_Q),     .A(D2888_Q));
KC_NAND4_X1 D2832 ( .Y(D2832_Y), .D(D2993_Y), .C(D16788_Y),     .B(D16787_Y), .A(D16786_Y));
KC_NAND4_X1 D2830 ( .Y(D2830_Y), .D(D2932_Y), .C(D2855_Y), .B(D2867_Y),     .A(D2880_Y));
KC_NAND4_X1 D2818 ( .Y(D2818_Y), .D(D14580_Y), .C(D16785_Y),     .B(D14583_Y), .A(D16783_Y));
KC_NAND4_X1 D2817 ( .Y(D2817_Y), .D(D2994_Y), .C(D16782_Y),     .B(D2992_Y), .A(D16784_Y));
KC_NAND4_X1 D2769 ( .Y(D2769_Y), .D(D2770_Y), .C(D2780_Y), .B(D2798_Q),     .A(D2797_Q));
KC_NAND4_X1 D2765 ( .Y(D2765_Y), .D(D2768_Y), .C(D2780_Y), .B(D2798_Q),     .A(D2799_Q));
KC_NAND4_X1 D2751 ( .Y(D2751_Y), .D(D2758_Y), .C(D2848_Y), .B(D2833_Y),     .A(D2757_Y));
KC_NAND4_X1 D2738 ( .Y(D2738_Y), .D(D2739_Y), .C(D2795_Q), .B(D2796_Q),     .A(D2782_Y));
KC_NAND4_X1 D2737 ( .Y(D2737_Y), .D(D2740_Y), .C(D2796_Q), .B(D2782_Y),     .A(D2794_Q));
KC_NAND4_X1 D2736 ( .Y(D2736_Y), .D(D2739_Y), .C(D2768_Y), .B(D2795_Q),     .A(D2799_Q));
KC_NAND4_X1 D2661 ( .Y(D2661_Y), .D(D89_Y), .C(D16192_Y), .B(D2659_Y),     .A(D2628_Y));
KC_NAND4_X1 D2494 ( .Y(D2494_Y), .D(D14206_Y), .C(D14210_Y),     .B(D2488_Y), .A(D14121_Y));
KC_NAND4_X1 D2493 ( .Y(D2493_Y), .D(D14217_Y), .C(D14209_Y),     .B(D2489_Y), .A(D14119_Y));
KC_NAND4_X1 D2486 ( .Y(D2486_Y), .D(D14198_Y), .C(D14279_Y),     .B(D14199_Y), .A(D2485_Y));
KC_NAND4_X1 D2425 ( .Y(D2425_Y), .D(D2380_Y), .C(D13633_Y),     .B(D13628_Y), .A(D13598_Y));
KC_NAND4_X1 D2419 ( .Y(D2419_Y), .D(D13655_Y), .C(D13664_Y),     .B(D13665_Y), .A(D13666_Y));
KC_NAND4_X1 D2406 ( .Y(D2406_Y), .D(D13954_Y), .C(D2404_Y),     .B(D13277_Y), .A(D13877_Y));
KC_NAND4_X1 D2362 ( .Y(D2362_Y), .D(D7670_Y), .C(D7669_Y), .B(D2343_Y),     .A(D12188_Y));
KC_NAND4_X1 D2321 ( .Y(D2321_Y), .D(D13049_Y), .C(D12938_Y),     .B(D12477_Y), .A(D2319_Y));
KC_NAND4_X1 D2306 ( .Y(D2306_Y), .D(D6281_Y), .C(D12207_Y),     .B(D12206_Y), .A(D11657_Y));
KC_NAND4_X1 D2276 ( .Y(D2276_Y), .D(D11928_Y), .C(D11898_Y),     .B(D11895_Y), .A(D11896_Y));
KC_NAND4_X1 D2270 ( .Y(D2270_Y), .D(D11984_Y), .C(D11886_Y),     .B(D2265_Y), .A(D11889_Y));
KC_NAND4_X1 D2269 ( .Y(D2269_Y), .D(D11983_Y), .C(D2314_Y),     .B(D11943_Y), .A(D11882_Y));
KC_NAND4_X1 D2200 ( .Y(D2200_Y), .D(D10893_Y), .C(D2197_Y),     .B(D2199_Y), .A(D10930_Y));
KC_NAND4_X1 D2188 ( .Y(D2188_Y), .D(D11405_Y), .C(D2186_Y),     .B(D10976_Y), .A(D2187_Y));
KC_NAND4_X1 D2132 ( .Y(D2132_Y), .D(D139_Y), .C(D10532_Y), .B(D2128_Y),     .A(D10534_Y));
KC_NAND4_X1 D2131 ( .Y(D2131_Y), .D(D2226_Y), .C(D10539_Y),     .B(D2130_Y), .A(D10527_Y));
KC_NAND4_X1 D2121 ( .Y(D2121_Y), .D(D8948_Y), .C(D9017_Y), .B(D9016_Y),     .A(D2086_Y));
KC_NAND4_X1 D2023 ( .Y(D2023_Y), .D(D8907_Y), .C(D8846_Y), .B(D8852_Y),     .A(D8911_Y));
KC_NAND4_X1 D2022 ( .Y(D2022_Y), .D(D8910_Y), .C(D2024_Y), .B(D289_Y),     .A(D2018_Y));
KC_NAND4_X1 D2021 ( .Y(D2021_Y), .D(D8853_Y), .C(D8845_Y), .B(D8847_Y),     .A(D8909_Y));
KC_NAND4_X1 D2020 ( .Y(D2020_Y), .D(D7445_Y), .C(D8849_Y), .B(D8926_Y),     .A(D2019_Y));
KC_NAND4_X1 D2012 ( .Y(D2012_Y), .D(D7568_Y), .C(D2011_Y), .B(D2006_Y),     .A(D8981_Y));
KC_NAND4_X1 D1982 ( .Y(D1982_Y), .D(D9573_Y), .C(D9521_Y), .B(D9549_Y),     .A(D1987_Y));
KC_NAND4_X1 D1876 ( .Y(D1876_Y), .D(D1879_Y), .C(D5828_Y), .B(D4434_Y),     .A(D1877_Y));
KC_NAND4_X1 D1851 ( .Y(D1851_Y), .D(D1860_Y), .C(D467_Y), .B(D7951_Y),     .A(D1917_Y));
KC_NAND4_X1 D1834 ( .Y(D1834_Y), .D(D8195_Y), .C(D12442_Y),     .B(D1833_Y), .A(D8614_Y));
KC_NAND4_X1 D1718 ( .Y(D1718_Y), .D(D213_Y), .C(D214_Y), .B(D7438_Y),     .A(D6019_Y));
KC_NAND4_X1 D1717 ( .Y(D1717_Y), .D(D4285_Y), .C(D1876_Y), .B(D7371_Y),     .A(D1585_Y));
KC_NAND4_X1 D1716 ( .Y(D1716_Y), .D(D5941_Y), .C(D1876_Y), .B(D5957_Y),     .A(D5985_Y));
KC_NAND4_X1 D1681 ( .Y(D1681_Y), .D(D7061_Y), .C(D1679_Y), .B(D7041_Y),     .A(D6978_Y));
KC_NAND4_X1 D1680 ( .Y(D1680_Y), .D(D7062_Y), .C(D1678_Y), .B(D7063_Y),     .A(D6982_Y));
KC_NAND4_X1 D1580 ( .Y(D1580_Y), .D(D4565_Y), .C(D4519_Y), .B(D4423_Y),     .A(D4559_Y));
KC_NAND4_X1 D1571 ( .Y(D1571_Y), .D(D4575_Y), .C(D4589_Y), .B(D4737_Y),     .A(D4640_Q));
KC_NAND4_X1 D1557 ( .Y(D1557_Y), .D(D5247_Y), .C(D6640_Y), .B(D5148_Y),     .A(D5208_Y));
KC_NAND4_X1 D1553 ( .Y(D1553_Y), .D(D3977_Y), .C(D5426_Y), .B(D1551_Y),     .A(D1550_Y));
KC_NAND4_X1 D1552 ( .Y(D1552_Y), .D(D3978_Y), .C(D5427_Y), .B(D967_Y),     .A(D5519_Y));
KC_NAND4_X1 D1434 ( .Y(D1434_Y), .D(D16779_Y), .C(D14578_Y),     .B(D2874_Y), .A(D15246_Y));
KC_NAND4_X1 D1433 ( .Y(D1433_Y), .D(D2952_Y), .C(D2952_Y), .B(D2903_Y),     .A(D2996_Y));
KC_NAND4_X1 D1429 ( .Y(D1429_Y), .D(D1432_Y), .C(D3146_Y), .B(D3138_Y),     .A(D3187_Q));
KC_NAND4_X1 D1342 ( .Y(D1342_Y), .D(D16660_Q), .C(D1320_Q),     .B(D16667_Y), .A(D16647_Y));
KC_NAND4_X1 D1276 ( .Y(D1276_Y), .D(D16426_Y), .C(D16380_Y),     .B(D16459_Q), .A(D1324_Q));
KC_NAND4_X1 D1275 ( .Y(D1275_Y), .D(D14425_Y), .C(D15169_Y),     .B(D15174_Y), .A(D14426_Y));
KC_NAND4_X1 D1273 ( .Y(D1273_Y), .D(D16443_Y), .C(D16380_Y),     .B(D1322_Q), .A(D1324_Q));
KC_NAND4_X1 D1271 ( .Y(D1271_Y), .D(D16443_Y), .C(D16414_Y),     .B(D16435_Y), .A(D1322_Q));
KC_NAND4_X1 D1270 ( .Y(D1270_Y), .D(D15999_Q), .C(D16012_Q),     .B(D15997_Q), .A(D16008_Q));
KC_NAND4_X1 D1264 ( .Y(D1264_Y), .D(D13129_Y), .C(D13102_Y),     .B(D1265_Y), .A(D12558_Y));
KC_NAND4_X1 D1255 ( .Y(D1255_Y), .D(D9911_Y), .C(D8618_Y), .B(D9857_Y),     .A(D1257_Y));
KC_NAND4_X1 D1252 ( .Y(D1252_Y), .D(D1370_Y), .C(D9856_Y), .B(D8649_Y),     .A(D8622_Y));
KC_NAND4_X1 D1179 ( .Y(D1179_Y), .D(D15722_Y), .C(D15945_Y),     .B(D15211_Y), .A(D15180_Y));
KC_NAND4_X1 D1177 ( .Y(D1177_Y), .D(D14321_Y), .C(D1277_Y),     .B(D14317_Y), .A(D14337_Y));
KC_NAND4_X1 D1095 ( .Y(D1095_Y), .D(D15809_Y), .C(D2594_Y),     .B(D15834_Y), .A(D15043_Y));
KC_NAND4_X1 D1092 ( .Y(D1092_Y), .D(D14303_Q), .C(D14306_Q),     .B(D14240_Q), .A(D14302_Q));
KC_NAND4_X1 D1087 ( .Y(D1087_Y), .D(D11988_Y), .C(D12482_Y),     .B(D11944_Y), .A(D11881_Y));
KC_NAND4_X1 D976 ( .Y(D976_Y), .D(D3948_Y), .C(D5445_Y), .B(D3909_Y),     .A(D5448_Y));
KC_NAND4_X1 D970 ( .Y(D970_Y), .D(D781_Y), .C(D8364_Y), .B(D8364_Y),     .A(D8364_Y));
KC_NAND4_X1 D872 ( .Y(D872_Y), .D(D14908_Y), .C(D14866_Y),     .B(D14128_Y), .A(D14851_Y));
KC_NAND4_X1 D741 ( .Y(D741_Y), .D(D9533_Y), .C(D8147_Q), .B(D9534_Y),     .A(D9544_Y));
KC_NAND4_X1 D740 ( .Y(D740_Y), .D(D3744_Y), .C(D5291_Y), .B(D5281_Y),     .A(D3794_Y));
KC_NAND4_X1 D739 ( .Y(D739_Y), .D(D8095_Y), .C(D824_Q), .B(D9526_Y),     .A(D9534_Y));
KC_NAND4_X1 D737 ( .Y(D737_Y), .D(D3746_Y), .C(D5282_Y), .B(D735_Y),     .A(D3787_Y));
KC_NAND4_X1 D558 ( .Y(D558_Y), .D(D11648_Y), .C(D11649_Y),     .B(D11653_Y), .A(D12197_Y));
KC_NAND4_X1 D496 ( .Y(D496_Y), .D(D12172_Y), .C(D12650_Y), .B(D510_Y),     .A(D12649_Y));
KC_NAND4_X1 D495 ( .Y(D495_Y), .D(D12643_Y), .C(D12233_Y),     .B(D12634_Y), .A(D12636_Y));
KC_NAND4_X1 D466 ( .Y(D466_Y), .D(D7919_Y), .C(D4981_Y), .B(D5096_Y),     .A(D3633_Y));
KC_NAND4_X1 D399 ( .Y(D399_Y), .D(D3306_Y), .C(D4911_Y), .B(D3446_Y),     .A(D3375_Q));
KC_NAND4_X1 D307 ( .Y(D307_Y), .D(D310_Y), .C(D4500_Y), .B(D3018_Y),     .A(D4502_Y));
KC_NAND4_X1 D284 ( .Y(D284_Y), .D(D8992_Y), .C(D7423_Y), .B(D8943_Y),     .A(D2076_Y));
KC_NAND4_X1 D244 ( .Y(D244_Y), .D(D7327_Y), .C(D5864_Y), .B(D5866_Y),     .A(D213_Y));
KC_NAND4_X1 D214 ( .Y(D214_Y), .D(D7107_Y), .C(D7254_Y), .B(D7255_Y),     .A(D7141_Y));
KC_NAND4_X1 D202 ( .Y(D202_Y), .D(D2027_Y), .C(D7183_Y), .B(D209_Y),     .A(D8741_Y));
KC_NAND4_X1 D67 ( .Y(D67_Y), .D(D2041_Y), .C(D2117_Y), .B(D9529_Y),     .A(D9483_Y));
KC_NOR2_X1 D16652 ( .Y(D16652_Y), .B(D16660_Q), .A(D1320_Q));
KC_NOR2_X1 D16622 ( .Y(D16622_Y), .B(D16570_Y), .A(D1320_Q));
KC_NOR2_X1 D16607 ( .Y(D16607_Y), .B(D16603_Y), .A(D16611_Q));
KC_NOR2_X1 D16603 ( .Y(D16603_Y), .B(D16600_Y), .A(D16595_Y));
KC_NOR2_X1 D16602 ( .Y(D16602_Y), .B(D16573_Y), .A(D16613_Q));
KC_NOR2_X1 D16572 ( .Y(D16572_Y), .B(D16613_Q), .A(D1374_Q));
KC_NOR2_X1 D16569 ( .Y(D16569_Y), .B(D16596_Y), .A(D16573_Y));
KC_NOR2_X1 D16563 ( .Y(D16563_Y), .B(D1340_Y), .A(D16561_Y));
KC_NOR2_X1 D16540 ( .Y(D16540_Y), .B(D16624_Y), .A(D16560_Y));
KC_NOR2_X1 D16539 ( .Y(D16539_Y), .B(D16535_Y), .A(D16556_Q));
KC_NOR2_X1 D16538 ( .Y(D16538_Y), .B(D16543_Y), .A(D16557_Q));
KC_NOR2_X1 D16534 ( .Y(D16534_Y), .B(D16771_Y), .A(D1385_Q));
KC_NOR2_X1 D16532 ( .Y(D16532_Y), .B(D16533_Y), .A(D7609_Y));
KC_NOR2_X1 D16530 ( .Y(D16530_Y), .B(D16550_Y), .A(D16654_Y));
KC_NOR2_X1 D16528 ( .Y(D16528_Y), .B(D16558_Q), .A(D16557_Q));
KC_NOR2_X1 D16522 ( .Y(D16522_Y), .B(D16496_Y), .A(D16521_Y));
KC_NOR2_X1 D16521 ( .Y(D16521_Y), .B(D16491_Y), .A(D16529_Y));
KC_NOR2_X1 D16499 ( .Y(D16499_Y), .B(D16488_Y), .A(D16536_Y));
KC_NOR2_X1 D16498 ( .Y(D16498_Y), .B(D16514_Y), .A(D16497_Y));
KC_NOR2_X1 D16497 ( .Y(D16497_Y), .B(D16500_Y), .A(D16771_Y));
KC_NOR2_X1 D16493 ( .Y(D16493_Y), .B(D16487_Y), .A(D16771_Y));
KC_NOR2_X1 D16484 ( .Y(D16484_Y), .B(D13988_Y), .A(D14651_Y));
KC_NOR2_X1 D16467 ( .Y(D16467_Y), .B(D13392_Y), .A(D16418_Y));
KC_NOR2_X1 D16465 ( .Y(D16465_Y), .B(D16407_Y), .A(D16462_Y));
KC_NOR2_X1 D16441 ( .Y(D16441_Y), .B(D16431_Y), .A(D16470_Q));
KC_NOR2_X1 D16436 ( .Y(D16436_Y), .B(D16459_Q), .A(D1324_Q));
KC_NOR2_X1 D16435 ( .Y(D16435_Y), .B(D16433_Y), .A(D16473_Q));
KC_NOR2_X1 D16434 ( .Y(D16434_Y), .B(D16439_Y), .A(D16433_Y));
KC_NOR2_X1 D16415 ( .Y(D16415_Y), .B(D16424_Y), .A(D16448_Y));
KC_NOR2_X1 D16414 ( .Y(D16414_Y), .B(D16438_Y), .A(D16444_Y));
KC_NOR2_X1 D16413 ( .Y(D16413_Y), .B(D16418_Y), .A(D16415_Y));
KC_NOR2_X1 D16412 ( .Y(D16412_Y), .B(D16431_Y), .A(D16443_Y));
KC_NOR2_X1 D16411 ( .Y(D16411_Y), .B(D16442_Y), .A(D16412_Y));
KC_NOR2_X1 D16372 ( .Y(D16372_Y), .B(D16458_Y), .A(D15475_Y));
KC_NOR2_X1 D16249 ( .Y(D16249_Y), .B(D16255_Y), .A(D7609_Y));
KC_NOR2_X1 D16248 ( .Y(D16248_Y), .B(D16260_Y), .A(D16245_Y));
KC_NOR2_X1 D16117 ( .Y(D16117_Y), .B(D16119_Y), .A(D16114_Y));
KC_NOR2_X1 D16116 ( .Y(D16116_Y), .B(D2591_Y), .A(D15270_Y));
KC_NOR2_X1 D16062 ( .Y(D16062_Y), .B(D16094_Y), .A(D16059_Y));
KC_NOR2_X1 D16057 ( .Y(D16057_Y), .B(D16043_Y), .A(D16094_Y));
KC_NOR2_X1 D16052 ( .Y(D16052_Y), .B(D16058_Y), .A(D16054_Y));
KC_NOR2_X1 D16051 ( .Y(D16051_Y), .B(D16094_Y), .A(D15335_Y));
KC_NOR2_X1 D16047 ( .Y(D16047_Y), .B(D16065_Y), .A(D16054_Y));
KC_NOR2_X1 D15968 ( .Y(D15968_Y), .B(D15962_Y), .A(D15935_S));
KC_NOR2_X1 D15963 ( .Y(D15963_Y), .B(D15964_Y), .A(D16012_Q));
KC_NOR2_X1 D15962 ( .Y(D15962_Y), .B(D15960_Y), .A(D15999_Q));
KC_NOR2_X1 D15900 ( .Y(D15900_Y), .B(D15899_Y), .A(D1229_Q));
KC_NOR2_X1 D15892 ( .Y(D15892_Y), .B(D15896_Y), .A(D15997_Q));
KC_NOR2_X1 D15891 ( .Y(D15891_Y), .B(D15892_Y), .A(D15939_S));
KC_NOR2_X1 D15889 ( .Y(D15889_Y), .B(D15900_Y), .A(D15857_S));
KC_NOR2_X1 D15731 ( .Y(D15731_Y), .B(D1070_Q), .A(D15728_Y));
KC_NOR2_X1 D15634 ( .Y(D15634_Y), .B(D14563_Y), .A(D15611_Y));
KC_NOR2_X1 D15616 ( .Y(D15616_Y), .B(D15611_Y), .A(D14830_Y));
KC_NOR2_X1 D15540 ( .Y(D15540_Y), .B(D15350_Y), .A(D15367_Y));
KC_NOR2_X1 D15539 ( .Y(D15539_Y), .B(D15531_Y), .A(D16200_Y));
KC_NOR2_X1 D15538 ( .Y(D15538_Y), .B(D15531_Y), .A(D8889_Y));
KC_NOR2_X1 D15537 ( .Y(D15537_Y), .B(D15362_Y), .A(D15349_Y));
KC_NOR2_X1 D15533 ( .Y(D15533_Y), .B(D15561_Y), .A(D15515_Y));
KC_NOR2_X1 D15532 ( .Y(D15532_Y), .B(D15362_Y), .A(D15359_Y));
KC_NOR2_X1 D15529 ( .Y(D15529_Y), .B(D15531_Y), .A(D15607_Y));
KC_NOR2_X1 D15528 ( .Y(D15528_Y), .B(D15531_Y), .A(D16132_Y));
KC_NOR2_X1 D15522 ( .Y(D15522_Y), .B(D16226_Q), .A(D15563_Y));
KC_NOR2_X1 D15506 ( .Y(D15506_Y), .B(D15611_Y), .A(D15607_Y));
KC_NOR2_X1 D15505 ( .Y(D15505_Y), .B(D816_Q), .A(D16242_Q));
KC_NOR2_X1 D15501 ( .Y(D15501_Y), .B(D15503_Y), .A(D15500_Y));
KC_NOR2_X1 D15500 ( .Y(D15500_Y), .B(D15476_Y), .A(D16242_Q));
KC_NOR2_X1 D15491 ( .Y(D15491_Y), .B(D16272_Y), .A(D15502_Y));
KC_NOR2_X1 D15490 ( .Y(D15490_Y), .B(D12140_Y), .A(D15562_Y));
KC_NOR2_X1 D15481 ( .Y(D15481_Y), .B(D14728_Y), .A(D15620_Y));
KC_NOR2_X1 D15480 ( .Y(D15480_Y), .B(D15469_Y), .A(D15562_Y));
KC_NOR2_X1 D15479 ( .Y(D15479_Y), .B(D14728_Y), .A(D15611_Y));
KC_NOR2_X1 D15478 ( .Y(D15478_Y), .B(D15470_Y), .A(D2604_Y));
KC_NOR2_X1 D15474 ( .Y(D15474_Y), .B(D16272_Y), .A(D15475_Y));
KC_NOR2_X1 D15464 ( .Y(D15464_Y), .B(D15470_Y), .A(D15480_Y));
KC_NOR2_X1 D15463 ( .Y(D15463_Y), .B(D15611_Y), .A(D12140_Y));
KC_NOR2_X1 D15406 ( .Y(D15406_Y), .B(D15267_Y), .A(D16056_Y));
KC_NOR2_X1 D15405 ( .Y(D15405_Y), .B(D15267_Y), .A(D564_Y));
KC_NOR2_X1 D15402 ( .Y(D15402_Y), .B(D15348_Y), .A(D15367_Y));
KC_NOR2_X1 D15372 ( .Y(D15372_Y), .B(D14625_Y), .A(D15514_Y));
KC_NOR2_X1 D15371 ( .Y(D15371_Y), .B(D15611_Y), .A(D12214_Y));
KC_NOR2_X1 D15359 ( .Y(D15359_Y), .B(D15375_Y), .A(D15563_Y));
KC_NOR2_X1 D15349 ( .Y(D15349_Y), .B(D14625_Y), .A(D15563_Y));
KC_NOR2_X1 D15348 ( .Y(D15348_Y), .B(D14625_Y), .A(D15611_Y));
KC_NOR2_X1 D15339 ( .Y(D15339_Y), .B(D15309_Y), .A(D15326_Y));
KC_NOR2_X1 D15338 ( .Y(D15338_Y), .B(D2654_Y), .A(D15339_Y));
KC_NOR2_X1 D15311 ( .Y(D15311_Y), .B(D15269_Y), .A(D574_Y));
KC_NOR2_X1 D15309 ( .Y(D15309_Y), .B(D15262_Y), .A(D15280_Y));
KC_NOR2_X1 D15308 ( .Y(D15308_Y), .B(D15300_Y), .A(D15310_Y));
KC_NOR2_X1 D15307 ( .Y(D15307_Y), .B(D15289_Y), .A(D15310_Y));
KC_NOR2_X1 D15305 ( .Y(D15305_Y), .B(D15394_Y), .A(D16067_Y));
KC_NOR2_X1 D15304 ( .Y(D15304_Y), .B(D15394_Y), .A(D570_Y));
KC_NOR2_X1 D15303 ( .Y(D15303_Y), .B(D570_Y), .A(D15306_Y));
KC_NOR2_X1 D15301 ( .Y(D15301_Y), .B(D16067_Y), .A(D15306_Y));
KC_NOR2_X1 D15297 ( .Y(D15297_Y), .B(D15302_Y), .A(D15276_Y));
KC_NOR2_X1 D15296 ( .Y(D15296_Y), .B(D15302_Y), .A(D15277_Y));
KC_NOR2_X1 D15295 ( .Y(D15295_Y), .B(D15288_Y), .A(D15284_Y));
KC_NOR2_X1 D15292 ( .Y(D15292_Y), .B(D15289_Y), .A(D15276_Y));
KC_NOR2_X1 D15287 ( .Y(D15287_Y), .B(D15300_Y), .A(D15276_Y));
KC_NOR2_X1 D15286 ( .Y(D15286_Y), .B(D15300_Y), .A(D15277_Y));
KC_NOR2_X1 D15285 ( .Y(D15285_Y), .B(D15289_Y), .A(D15277_Y));
KC_NOR2_X1 D15284 ( .Y(D15284_Y), .B(D15279_Y), .A(D16090_Y));
KC_NOR2_X1 D15283 ( .Y(D15283_Y), .B(D16088_Y), .A(D15290_Y));
KC_NOR2_X1 D15282 ( .Y(D15282_Y), .B(D15262_Y), .A(D16089_Y));
KC_NOR2_X1 D15275 ( .Y(D15275_Y), .B(D15300_Y), .A(D15278_Y));
KC_NOR2_X1 D15274 ( .Y(D15274_Y), .B(D15289_Y), .A(D15278_Y));
KC_NOR2_X1 D15273 ( .Y(D15273_Y), .B(D16053_Y), .A(D16090_Y));
KC_NOR2_X1 D15272 ( .Y(D15272_Y), .B(D15290_Y), .A(D16053_Y));
KC_NOR2_X1 D15242 ( .Y(D15242_Y), .B(D15243_Y), .A(D15258_Y));
KC_NOR2_X1 D15225 ( .Y(D15225_Y), .B(D15224_Y), .A(D16008_Q));
KC_NOR2_X1 D15223 ( .Y(D15223_Y), .B(D15225_Y), .A(D15126_S));
KC_NOR2_X1 D15182 ( .Y(D15182_Y), .B(D15971_Y), .A(D15993_Q));
KC_NOR2_X1 D15176 ( .Y(D15176_Y), .B(D15110_Y), .A(D16011_Q));
KC_NOR2_X1 D15166 ( .Y(D15166_Y), .B(D15182_Y), .A(D15942_S));
KC_NOR2_X1 D15105 ( .Y(D15105_Y), .B(D15176_Y), .A(D15127_S));
KC_NOR2_X1 D15100 ( .Y(D15100_Y), .B(D15101_Y), .A(D16009_Q));
KC_NOR2_X1 D15098 ( .Y(D15098_Y), .B(D15100_Y), .A(D15071_S));
KC_NOR2_X1 D15041 ( .Y(D15041_Y), .B(D1095_Y), .A(D15022_Y));
KC_NOR2_X1 D15024 ( .Y(D15024_Y), .B(D15042_Y), .A(D15037_Y));
KC_NOR2_X1 D14958 ( .Y(D14958_Y), .B(D14952_Y), .A(D14820_Y));
KC_NOR2_X1 D14954 ( .Y(D14954_Y), .B(D14940_Y), .A(D14835_Y));
KC_NOR2_X1 D14945 ( .Y(D14945_Y), .B(D14266_Q), .A(D14946_Y));
KC_NOR2_X1 D14936 ( .Y(D14936_Y), .B(D15720_Y), .A(D14924_Y));
KC_NOR2_X1 D14932 ( .Y(D14932_Y), .B(D14929_Y), .A(D14836_Y));
KC_NOR2_X1 D14920 ( .Y(D14920_Y), .B(D15714_Y), .A(D14921_Y));
KC_NOR2_X1 D14853 ( .Y(D14853_Y), .B(D14854_Y), .A(D13156_Y));
KC_NOR2_X1 D14850 ( .Y(D14850_Y), .B(D14854_Y), .A(D6111_Y));
KC_NOR2_X1 D14846 ( .Y(D14846_Y), .B(D14854_Y), .A(D16080_Y));
KC_NOR2_X1 D14840 ( .Y(D14840_Y), .B(D14854_Y), .A(D14830_Y));
KC_NOR2_X1 D14829 ( .Y(D14829_Y), .B(D14563_Y), .A(D15562_Y));
KC_NOR2_X1 D14813 ( .Y(D14813_Y), .B(D16226_Q), .A(D15562_Y));
KC_NOR2_X1 D14750 ( .Y(D14750_Y), .B(D14564_Y), .A(D15563_Y));
KC_NOR2_X1 D14743 ( .Y(D14743_Y), .B(D16524_Y), .A(D14665_Y));
KC_NOR2_X1 D14742 ( .Y(D14742_Y), .B(D13935_Y), .A(D13392_Y));
KC_NOR2_X1 D14734 ( .Y(D14734_Y), .B(D13330_Y), .A(D16263_Y));
KC_NOR2_X1 D14715 ( .Y(D14715_Y), .B(D14714_Y), .A(D13963_Y));
KC_NOR2_X1 D14714 ( .Y(D14714_Y), .B(D13973_Y), .A(D645_Y));
KC_NOR2_X1 D14654 ( .Y(D14654_Y), .B(D13971_Y), .A(D16117_Y));
KC_NOR2_X1 D14635 ( .Y(D14635_Y), .B(D13952_Y), .A(D13997_Q));
KC_NOR2_X1 D14634 ( .Y(D14634_Y), .B(D721_Q), .A(D722_Q));
KC_NOR2_X1 D14627 ( .Y(D14627_Y), .B(D14652_Y), .A(D14641_Y));
KC_NOR2_X1 D14624 ( .Y(D14624_Y), .B(D12214_Y), .A(D15563_Y));
KC_NOR2_X1 D14539 ( .Y(D14539_Y), .B(D14534_Y), .A(D14543_Y));
KC_NOR2_X1 D14530 ( .Y(D14530_Y), .B(D14528_Y), .A(D14531_Y));
KC_NOR2_X1 D14529 ( .Y(D14529_Y), .B(D14557_Y), .A(D14518_Q));
KC_NOR2_X1 D14528 ( .Y(D14528_Y), .B(D14544_Y), .A(D14557_Y));
KC_NOR2_X1 D14500 ( .Y(D14500_Y), .B(D14501_Y), .A(D2512_Y));
KC_NOR2_X1 D14499 ( .Y(D14499_Y), .B(D14497_Y), .A(D2512_Y));
KC_NOR2_X1 D14483 ( .Y(D14483_Y), .B(D14485_Y), .A(D14478_Y));
KC_NOR2_X1 D14479 ( .Y(D14479_Y), .B(D15161_Y), .A(D1380_Q));
KC_NOR2_X1 D14451 ( .Y(D14451_Y), .B(D14453_Y), .A(D15235_Q));
KC_NOR2_X1 D14443 ( .Y(D14443_Y), .B(D14417_Y), .A(D14496_Q));
KC_NOR2_X1 D14412 ( .Y(D14412_Y), .B(D14415_Y), .A(D14452_Y));
KC_NOR2_X1 D14403 ( .Y(D14403_Y), .B(D14404_Y), .A(D14400_Y));
KC_NOR2_X1 D14399 ( .Y(D14399_Y), .B(D1268_Y), .A(D14493_Q));
KC_NOR2_X1 D14358 ( .Y(D14358_Y), .B(D14438_Y), .A(D16014_Q));
KC_NOR2_X1 D14353 ( .Y(D14353_Y), .B(D14344_Y), .A(D14354_Y));
KC_NOR2_X1 D14352 ( .Y(D14352_Y), .B(D14350_Y), .A(D15230_Q));
KC_NOR2_X1 D14334 ( .Y(D14334_Y), .B(D14335_Y), .A(D1379_Q));
KC_NOR2_X1 D14322 ( .Y(D14322_Y), .B(D14360_Y), .A(D14359_Y));
KC_NOR2_X1 D14276 ( .Y(D14276_Y), .B(D14290_Y), .A(D14277_Y));
KC_NOR2_X1 D14220 ( .Y(D14220_Y), .B(D14133_Y), .A(D874_Y));
KC_NOR2_X1 D14130 ( .Y(D14130_Y), .B(D14018_Y), .A(D14134_Y));
KC_NOR2_X1 D14129 ( .Y(D14129_Y), .B(D14137_Y), .A(D13379_Y));
KC_NOR2_X1 D14126 ( .Y(D14126_Y), .B(D14132_Y), .A(D13379_Y));
KC_NOR2_X1 D14113 ( .Y(D14113_Y), .B(D14018_Y), .A(D14133_Y));
KC_NOR2_X1 D14046 ( .Y(D14046_Y), .B(D15508_Y), .A(D13947_Y));
KC_NOR2_X1 D14038 ( .Y(D14038_Y), .B(D14045_Y), .A(D14097_Y));
KC_NOR2_X1 D14034 ( .Y(D14034_Y), .B(D14045_Y), .A(D14065_Y));
KC_NOR2_X1 D14033 ( .Y(D14033_Y), .B(D2478_Y), .A(D14065_Y));
KC_NOR2_X1 D14029 ( .Y(D14029_Y), .B(D14038_Y), .A(D14034_Y));
KC_NOR2_X1 D14009 ( .Y(D14009_Y), .B(D14018_Y), .A(D14137_Y));
KC_NOR2_X1 D14008 ( .Y(D14008_Y), .B(D13313_Y), .A(D14018_Y));
KC_NOR2_X1 D13955 ( .Y(D13955_Y), .B(D13186_Y), .A(D7609_Y));
KC_NOR2_X1 D13950 ( .Y(D13950_Y), .B(D15394_Y), .A(D16226_Q));
KC_NOR2_X1 D13946 ( .Y(D13946_Y), .B(D637_Y), .A(D14619_Y));
KC_NOR2_X1 D13945 ( .Y(D13945_Y), .B(D14629_Y), .A(D14689_Q));
KC_NOR2_X1 D13937 ( .Y(D13937_Y), .B(D13941_Y), .A(D13936_Y));
KC_NOR2_X1 D13932 ( .Y(D13932_Y), .B(D13926_Y), .A(D14616_Y));
KC_NOR2_X1 D13929 ( .Y(D13929_Y), .B(D16559_Y), .A(D13936_Y));
KC_NOR2_X1 D13928 ( .Y(D13928_Y), .B(D13964_Y), .A(D13929_Y));
KC_NOR2_X1 D13902 ( .Y(D13902_Y), .B(D2408_Y), .A(D7668_Y));
KC_NOR2_X1 D13778 ( .Y(D13778_Y), .B(D14405_Y), .A(D14445_Y));
KC_NOR2_X1 D13723 ( .Y(D13723_Y), .B(D10266_Y), .A(D13769_Y));
KC_NOR2_X1 D13722 ( .Y(D13722_Y), .B(D14329_Y), .A(D13726_Y));
KC_NOR2_X1 D13668 ( .Y(D13668_Y), .B(D13672_Y), .A(D13770_Q));
KC_NOR2_X1 D13663 ( .Y(D13663_Y), .B(D13656_Y), .A(D13536_Y));
KC_NOR2_X1 D13662 ( .Y(D13662_Y), .B(D14222_Y), .A(D13536_Y));
KC_NOR2_X1 D13566 ( .Y(D13566_Y), .B(D12955_Y), .A(D13559_Y));
KC_NOR2_X1 D13553 ( .Y(D13553_Y), .B(D13549_Y), .A(D13338_Y));
KC_NOR2_X1 D13552 ( .Y(D13552_Y), .B(D2430_Y), .A(D13559_Y));
KC_NOR2_X1 D13540 ( .Y(D13540_Y), .B(D14132_Y), .A(D874_Y));
KC_NOR2_X1 D13539 ( .Y(D13539_Y), .B(D13297_Y), .A(D13559_Y));
KC_NOR2_X1 D13538 ( .Y(D13538_Y), .B(D13295_Y), .A(D13559_Y));
KC_NOR2_X1 D13535 ( .Y(D13535_Y), .B(D13472_Y), .A(D962_Y));
KC_NOR2_X1 D13532 ( .Y(D13532_Y), .B(D13472_Y), .A(D13531_Y));
KC_NOR2_X1 D13531 ( .Y(D13531_Y), .B(D13330_Y), .A(D14137_Y));
KC_NOR2_X1 D13529 ( .Y(D13529_Y), .B(D13472_Y), .A(D13528_Y));
KC_NOR2_X1 D13528 ( .Y(D13528_Y), .B(D13330_Y), .A(D14134_Y));
KC_NOR2_X1 D13471 ( .Y(D13471_Y), .B(D7669_Y), .A(D13338_Y));
KC_NOR2_X1 D13464 ( .Y(D13464_Y), .B(D13470_Y), .A(D13477_Y));
KC_NOR2_X1 D13454 ( .Y(D13454_Y), .B(D13448_Y), .A(D13323_Y));
KC_NOR2_X1 D13443 ( .Y(D13443_Y), .B(D866_Y), .A(D13536_Y));
KC_NOR2_X1 D13442 ( .Y(D13442_Y), .B(D13448_Y), .A(D13536_Y));
KC_NOR2_X1 D13441 ( .Y(D13441_Y), .B(D13559_Y), .A(D2429_Y));
KC_NOR2_X1 D13435 ( .Y(D13435_Y), .B(D13421_Y), .A(D13409_Y));
KC_NOR2_X1 D13417 ( .Y(D13417_Y), .B(D2433_Y), .A(D13559_Y));
KC_NOR2_X1 D13410 ( .Y(D13410_Y), .B(D812_Y), .A(D13977_Y));
KC_NOR2_X1 D13354 ( .Y(D13354_Y), .B(D13221_Y), .A(D13348_Y));
KC_NOR2_X1 D13353 ( .Y(D13353_Y), .B(D13269_Q), .A(D13267_Q));
KC_NOR2_X1 D13352 ( .Y(D13352_Y), .B(D13358_Y), .A(D13267_Q));
KC_NOR2_X1 D13337 ( .Y(D13337_Y), .B(D13369_Y), .A(D13365_Y));
KC_NOR2_X1 D13336 ( .Y(D13336_Y), .B(D13395_Q), .A(D13396_Q));
KC_NOR2_X1 D13335 ( .Y(D13335_Y), .B(D13395_Q), .A(D13346_Y));
KC_NOR2_X1 D13329 ( .Y(D13329_Y), .B(D7609_Y), .A(D13337_Y));
KC_NOR2_X1 D13328 ( .Y(D13328_Y), .B(D12816_Y), .A(D12756_Q));
KC_NOR2_X1 D13327 ( .Y(D13327_Y), .B(D13356_Y), .A(D13357_Y));
KC_NOR2_X1 D13326 ( .Y(D13326_Y), .B(D13389_Y), .A(D10207_Y));
KC_NOR2_X1 D13325 ( .Y(D13325_Y), .B(D13356_Y), .A(D13339_Y));
KC_NOR2_X1 D13318 ( .Y(D13318_Y), .B(D2312_Y), .A(D2353_Y));
KC_NOR2_X1 D13317 ( .Y(D13317_Y), .B(D7670_Y), .A(D2353_Y));
KC_NOR2_X1 D13316 ( .Y(D13316_Y), .B(D161_Y), .A(D12241_Y));
KC_NOR2_X1 D13315 ( .Y(D13315_Y), .B(D7668_Y), .A(D12241_Y));
KC_NOR2_X1 D13314 ( .Y(D13314_Y), .B(D14017_Y), .A(D14665_Y));
KC_NOR2_X1 D13312 ( .Y(D13312_Y), .B(D13334_Y), .A(D13977_Y));
KC_NOR2_X1 D13311 ( .Y(D13311_Y), .B(D12279_Q), .A(D12277_Q));
KC_NOR2_X1 D13306 ( .Y(D13306_Y), .B(D2343_Y), .A(D12241_Y));
KC_NOR2_X1 D13305 ( .Y(D13305_Y), .B(D13474_Y), .A(D13306_Y));
KC_NOR2_X1 D13299 ( .Y(D13299_Y), .B(D13296_Y), .A(D13298_Y));
KC_NOR2_X1 D13298 ( .Y(D13298_Y), .B(D13474_Y), .A(D13478_Y));
KC_NOR2_X1 D13297 ( .Y(D13297_Y), .B(D13301_Y), .A(D7668_Y));
KC_NOR2_X1 D13296 ( .Y(D13296_Y), .B(D13474_Y), .A(D13315_Y));
KC_NOR2_X1 D13295 ( .Y(D13295_Y), .B(D13301_Y), .A(D2343_Y));
KC_NOR2_X1 D13294 ( .Y(D13294_Y), .B(D13475_Y), .A(D2343_Y));
KC_NOR2_X1 D13293 ( .Y(D13293_Y), .B(D7668_Y), .A(D12732_Y));
KC_NOR2_X1 D13292 ( .Y(D13292_Y), .B(D13302_Y), .A(D12279_Q));
KC_NOR2_X1 D13233 ( .Y(D13233_Y), .B(D13364_Y), .A(D13246_Y));
KC_NOR2_X1 D13229 ( .Y(D13229_Y), .B(D2407_Y), .A(D12191_Y));
KC_NOR2_X1 D13221 ( .Y(D13221_Y), .B(D13361_Y), .A(D15508_Y));
KC_NOR2_X1 D13218 ( .Y(D13218_Y), .B(D2362_Y), .A(D12191_Y));
KC_NOR2_X1 D13184 ( .Y(D13184_Y), .B(D2408_Y), .A(D2343_Y));
KC_NOR2_X1 D12949 ( .Y(D12949_Y), .B(D12963_Y), .A(D12931_Y));
KC_NOR2_X1 D12944 ( .Y(D12944_Y), .B(D13010_Y), .A(D13338_Y));
KC_NOR2_X1 D12939 ( .Y(D12939_Y), .B(D13536_Y), .A(D12872_Y));
KC_NOR2_X1 D12891 ( .Y(D12891_Y), .B(D12909_Y), .A(D13392_Y));
KC_NOR2_X1 D12889 ( .Y(D12889_Y), .B(D13501_Y), .A(D12861_Y));
KC_NOR2_X1 D12885 ( .Y(D12885_Y), .B(D12908_Y), .A(D13392_Y));
KC_NOR2_X1 D12884 ( .Y(D12884_Y), .B(D12910_Y), .A(D13392_Y));
KC_NOR2_X1 D12883 ( .Y(D12883_Y), .B(D12911_Y), .A(D13392_Y));
KC_NOR2_X1 D12882 ( .Y(D12882_Y), .B(D2400_Y), .A(D13392_Y));
KC_NOR2_X1 D12881 ( .Y(D12881_Y), .B(D852_Q), .A(D814_Q));
KC_NOR2_X1 D12877 ( .Y(D12877_Y), .B(D956_Q), .A(D146_Q));
KC_NOR2_X1 D12872 ( .Y(D12872_Y), .B(D12899_Y), .A(D2395_Y));
KC_NOR2_X1 D12812 ( .Y(D12812_Y), .B(D12844_Y), .A(D13392_Y));
KC_NOR2_X1 D12811 ( .Y(D12811_Y), .B(D12841_Y), .A(D13392_Y));
KC_NOR2_X1 D12804 ( .Y(D12804_Y), .B(D12754_Q), .A(D12704_Y));
KC_NOR2_X1 D12803 ( .Y(D12803_Y), .B(D12805_Y), .A(D12858_Q));
KC_NOR2_X1 D12802 ( .Y(D12802_Y), .B(D12862_Y), .A(D13392_Y));
KC_NOR2_X1 D12789 ( .Y(D12789_Y), .B(D12855_Q), .A(D12856_Q));
KC_NOR2_X1 D12783 ( .Y(D12783_Y), .B(D15498_Y), .A(D13361_Y));
KC_NOR2_X1 D12782 ( .Y(D12782_Y), .B(D12810_Y), .A(D13361_Y));
KC_NOR2_X1 D12781 ( .Y(D12781_Y), .B(D12785_Y), .A(D13372_Y));
KC_NOR2_X1 D12780 ( .Y(D12780_Y), .B(D13361_Y), .A(D12795_Y));
KC_NOR2_X1 D12779 ( .Y(D12779_Y), .B(D14730_Y), .A(D13361_Y));
KC_NOR2_X1 D12721 ( .Y(D12721_Y), .B(D12751_Y), .A(D12713_Y));
KC_NOR2_X1 D12719 ( .Y(D12719_Y), .B(D12250_Y), .A(D12298_Y));
KC_NOR2_X1 D12707 ( .Y(D12707_Y), .B(D12700_Y), .A(D699_Q));
KC_NOR2_X1 D12698 ( .Y(D12698_Y), .B(D12753_Q), .A(D12756_Q));
KC_NOR2_X1 D12695 ( .Y(D12695_Y), .B(D13344_Y), .A(D13349_Y));
KC_NOR2_X1 D12694 ( .Y(D12694_Y), .B(D13373_Y), .A(D13344_Y));
KC_NOR2_X1 D12692 ( .Y(D12692_Y), .B(D12722_Y), .A(D14785_Y));
KC_NOR2_X1 D12660 ( .Y(D12660_Y), .B(D12733_Y), .A(D12756_Q));
KC_NOR2_X1 D12659 ( .Y(D12659_Y), .B(D2361_Y), .A(D12191_Y));
KC_NOR2_X1 D12323 ( .Y(D12323_Y), .B(D12355_Q), .A(D843_Q));
KC_NOR2_X1 D12312 ( .Y(D12312_Y), .B(D12316_Y), .A(D12782_Y));
KC_NOR2_X1 D12256 ( .Y(D12256_Y), .B(D12209_Y), .A(D12819_Y));
KC_NOR2_X1 D12254 ( .Y(D12254_Y), .B(D2306_Y), .A(D2358_Y));
KC_NOR2_X1 D12253 ( .Y(D12253_Y), .B(D12297_Y), .A(D12819_Y));
KC_NOR2_X1 D12252 ( .Y(D12252_Y), .B(D12251_Y), .A(D12819_Y));
KC_NOR2_X1 D12251 ( .Y(D12251_Y), .B(D12362_Y), .A(D12801_Y));
KC_NOR2_X1 D12250 ( .Y(D12250_Y), .B(D2306_Y), .A(D12190_Y));
KC_NOR2_X1 D12249 ( .Y(D12249_Y), .B(D717_Q), .A(D12356_Q));
KC_NOR2_X1 D12247 ( .Y(D12247_Y), .B(D12705_Y), .A(D12279_Q));
KC_NOR2_X1 D12245 ( .Y(D12245_Y), .B(D12701_Y), .A(D12279_Q));
KC_NOR2_X1 D12239 ( .Y(D12239_Y), .B(D2329_Y), .A(D12185_Q));
KC_NOR2_X1 D12207 ( .Y(D12207_Y), .B(D1954_Y), .A(D14806_Y));
KC_NOR2_X1 D12206 ( .Y(D12206_Y), .B(D10179_Y), .A(D11660_Y));
KC_NOR2_X1 D12202 ( .Y(D12202_Y), .B(D9371_Y), .A(D2353_Y));
KC_NOR2_X1 D12198 ( .Y(D12198_Y), .B(D12200_Y), .A(D7782_Y));
KC_NOR2_X1 D12193 ( .Y(D12193_Y), .B(D11655_Y), .A(D11657_Y));
KC_NOR2_X1 D12188 ( .Y(D12188_Y), .B(D12205_Y), .A(D9371_Y));
KC_NOR2_X1 D12187 ( .Y(D12187_Y), .B(D12192_Y), .A(D12191_Y));
KC_NOR2_X1 D12184 ( .Y(D12184_Y), .B(D12178_Q), .A(D11183_Y));
KC_NOR2_X1 D12026 ( .Y(D12026_Y), .B(D12030_Y), .A(D12013_Y));
KC_NOR2_X1 D12025 ( .Y(D12025_Y), .B(D11963_Y), .A(D12017_Y));
KC_NOR2_X1 D12024 ( .Y(D12024_Y), .B(D12030_Y), .A(D12027_Y));
KC_NOR2_X1 D12023 ( .Y(D12023_Y), .B(D12031_Y), .A(D12027_Y));
KC_NOR2_X1 D12016 ( .Y(D12016_Y), .B(D12032_Y), .A(D12027_Y));
KC_NOR2_X1 D12015 ( .Y(D12015_Y), .B(D12032_Y), .A(D12013_Y));
KC_NOR2_X1 D12012 ( .Y(D12012_Y), .B(D11965_Y), .A(D12017_Y));
KC_NOR2_X1 D12011 ( .Y(D12011_Y), .B(D12031_Y), .A(D12013_Y));
KC_NOR2_X1 D12010 ( .Y(D12010_Y), .B(D11964_Y), .A(D12017_Y));
KC_NOR2_X1 D11953 ( .Y(D11953_Y), .B(D11962_Y), .A(D11945_Y));
KC_NOR2_X1 D11952 ( .Y(D11952_Y), .B(D11904_Y), .A(D11941_Y));
KC_NOR2_X1 D11951 ( .Y(D11951_Y), .B(D11959_Y), .A(D11946_Y));
KC_NOR2_X1 D11950 ( .Y(D11950_Y), .B(D11960_Y), .A(D11945_Y));
KC_NOR2_X1 D11949 ( .Y(D11949_Y), .B(D11961_Y), .A(D11955_Y));
KC_NOR2_X1 D11948 ( .Y(D11948_Y), .B(D11962_Y), .A(D11955_Y));
KC_NOR2_X1 D11615 ( .Y(D11615_Y), .B(D8903_Y), .A(D11672_Q));
KC_NOR2_X1 D11551 ( .Y(D11551_Y), .B(D6792_Y), .A(D5214_Y));
KC_NOR2_X1 D11546 ( .Y(D11546_Y), .B(D6792_Y), .A(D5214_Y));
KC_NOR2_X1 D11363 ( .Y(D11363_Y), .B(D6792_Y), .A(D5214_Y));
KC_NOR2_X1 D11145 ( .Y(D11145_Y), .B(D6792_Y), .A(D5214_Y));
KC_NOR2_X1 D10917 ( .Y(D10917_Y), .B(D10937_Y), .A(D10972_Y));
KC_NOR2_X1 D10913 ( .Y(D10913_Y), .B(D10987_Y), .A(D10967_Y));
KC_NOR2_X1 D10912 ( .Y(D10912_Y), .B(D10987_Y), .A(D10905_Y));
KC_NOR2_X1 D10904 ( .Y(D10904_Y), .B(D10986_Y), .A(D10967_Y));
KC_NOR2_X1 D10903 ( .Y(D10903_Y), .B(D10937_Y), .A(D10936_Y));
KC_NOR2_X1 D10902 ( .Y(D10902_Y), .B(D10986_Y), .A(D10905_Y));
KC_NOR2_X1 D10856 ( .Y(D10856_Y), .B(D2146_Y), .A(D2135_Y));
KC_NOR2_X1 D10854 ( .Y(D10854_Y), .B(D6792_Y), .A(D5214_Y));
KC_NOR2_X1 D10757 ( .Y(D10757_Y), .B(D10771_Y), .A(D10664_Y));
KC_NOR2_X1 D10750 ( .Y(D10750_Y), .B(D10768_Y), .A(D10734_Y));
KC_NOR2_X1 D10749 ( .Y(D10749_Y), .B(D10771_Y), .A(D10734_Y));
KC_NOR2_X1 D10745 ( .Y(D10745_Y), .B(D10763_Y), .A(D10729_Y));
KC_NOR2_X1 D10743 ( .Y(D10743_Y), .B(D10763_Y), .A(D10747_Y));
KC_NOR2_X1 D10742 ( .Y(D10742_Y), .B(D10761_Y), .A(D10747_Y));
KC_NOR2_X1 D10672 ( .Y(D10672_Y), .B(D10764_Y), .A(D10734_Y));
KC_NOR2_X1 D10663 ( .Y(D10663_Y), .B(D10764_Y), .A(D10664_Y));
KC_NOR2_X1 D10541 ( .Y(D10541_Y), .B(D10486_Y), .A(D10536_Y));
KC_NOR2_X1 D10535 ( .Y(D10535_Y), .B(D10485_Y), .A(D10536_Y));
KC_NOR2_X1 D10520 ( .Y(D10520_Y), .B(D10458_Y), .A(D8365_Y));
KC_NOR2_X1 D10463 ( .Y(D10463_Y), .B(D10464_Y), .A(D8365_Y));
KC_NOR2_X1 D10462 ( .Y(D10462_Y), .B(D10466_Y), .A(D8365_Y));
KC_NOR2_X1 D10457 ( .Y(D10457_Y), .B(D10459_Y), .A(D8365_Y));
KC_NOR2_X1 D10456 ( .Y(D10456_Y), .B(D10460_Y), .A(D8365_Y));
KC_NOR2_X1 D10450 ( .Y(D10450_Y), .B(D10452_Y), .A(D8365_Y));
KC_NOR2_X1 D10449 ( .Y(D10449_Y), .B(D10451_Y), .A(D8365_Y));
KC_NOR2_X1 D10448 ( .Y(D10448_Y), .B(D10447_Y), .A(D8365_Y));
KC_NOR2_X1 D10394 ( .Y(D10394_Y), .B(D1107_Y), .A(D10967_Y));
KC_NOR2_X1 D10195 ( .Y(D10195_Y), .B(D10310_Y), .A(D10214_Y));
KC_NOR2_X1 D10168 ( .Y(D10168_Y), .B(D10027_Y), .A(D2162_Y));
KC_NOR2_X1 D10167 ( .Y(D10167_Y), .B(D2086_Y), .A(D2162_Y));
KC_NOR2_X1 D10104 ( .Y(D10104_Y), .B(D9175_Y), .A(D1711_Y));
KC_NOR2_X1 D10099 ( .Y(D10099_Y), .B(D10067_Y), .A(D10098_Y));
KC_NOR2_X1 D10098 ( .Y(D10098_Y), .B(D10088_Y), .A(D10070_Y));
KC_NOR2_X1 D10083 ( .Y(D10083_Y), .B(D10091_Y), .A(D10090_Y));
KC_NOR2_X1 D10079 ( .Y(D10079_Y), .B(D2122_Y), .A(D10093_Y));
KC_NOR2_X1 D10078 ( .Y(D10078_Y), .B(D374_Y), .A(D10075_Y));
KC_NOR2_X1 D10077 ( .Y(D10077_Y), .B(D10100_Y), .A(D10075_Y));
KC_NOR2_X1 D10074 ( .Y(D10074_Y), .B(D368_Y), .A(D10075_Y));
KC_NOR2_X1 D10073 ( .Y(D10073_Y), .B(D10077_Y), .A(D10070_Y));
KC_NOR2_X1 D10072 ( .Y(D10072_Y), .B(D10087_Y), .A(D10074_Y));
KC_NOR2_X1 D10070 ( .Y(D10070_Y), .B(D10100_Y), .A(D10068_Y));
KC_NOR2_X1 D10067 ( .Y(D10067_Y), .B(D368_Y), .A(D10068_Y));
KC_NOR2_X1 D9967 ( .Y(D9967_Y), .B(D9922_Y), .A(D9973_Y));
KC_NOR2_X1 D9966 ( .Y(D9966_Y), .B(D9962_Y), .A(D9972_Y));
KC_NOR2_X1 D9965 ( .Y(D9965_Y), .B(D9922_Y), .A(D9971_Y));
KC_NOR2_X1 D9964 ( .Y(D9964_Y), .B(D9922_Y), .A(D9972_Y));
KC_NOR2_X1 D9963 ( .Y(D9963_Y), .B(D9962_Y), .A(D9973_Y));
KC_NOR2_X1 D9962 ( .Y(D9962_Y), .B(D8768_Y), .A(D201_Y));
KC_NOR2_X1 D9959 ( .Y(D9959_Y), .B(D8737_Y), .A(D8768_Y));
KC_NOR2_X1 D9958 ( .Y(D9958_Y), .B(D8737_Y), .A(D9961_Y));
KC_NOR2_X1 D9957 ( .Y(D9957_Y), .B(D8737_Y), .A(D9960_Y));
KC_NOR2_X1 D9956 ( .Y(D9956_Y), .B(D9962_Y), .A(D223_Y));
KC_NOR2_X1 D9955 ( .Y(D9955_Y), .B(D9962_Y), .A(D9971_Y));
KC_NOR2_X1 D9925 ( .Y(D9925_Y), .B(D9927_Y), .A(D9940_Y));
KC_NOR2_X1 D9922 ( .Y(D9922_Y), .B(D7781_Y), .A(D201_Y));
KC_NOR2_X1 D9751 ( .Y(D9751_Y), .B(D9750_Y), .A(D8365_Y));
KC_NOR2_X1 D9749 ( .Y(D9749_Y), .B(D9682_Y), .A(D8365_Y));
KC_NOR2_X1 D9748 ( .Y(D9748_Y), .B(D8503_Y), .A(D8365_Y));
KC_NOR2_X1 D9747 ( .Y(D9747_Y), .B(D9752_Y), .A(D8365_Y));
KC_NOR2_X1 D9745 ( .Y(D9745_Y), .B(D9744_Y), .A(D8365_Y));
KC_NOR2_X1 D9734 ( .Y(D9734_Y), .B(D9740_Y), .A(D8422_Y));
KC_NOR2_X1 D9732 ( .Y(D9732_Y), .B(D9736_Y), .A(D8365_Y));
KC_NOR2_X1 D9731 ( .Y(D9731_Y), .B(D9727_Y), .A(D8422_Y));
KC_NOR2_X1 D9730 ( .Y(D9730_Y), .B(D9733_Y), .A(D8422_Y));
KC_NOR2_X1 D9729 ( .Y(D9729_Y), .B(D9741_Y), .A(D8422_Y));
KC_NOR2_X1 D9725 ( .Y(D9725_Y), .B(D8542_Y), .A(D8534_Y));
KC_NOR2_X1 D9599 ( .Y(D9599_Y), .B(D2061_Y), .A(D9504_Y));
KC_NOR2_X1 D9598 ( .Y(D9598_Y), .B(D9496_Y), .A(D9494_Y));
KC_NOR2_X1 D9534 ( .Y(D9534_Y), .B(D9575_Q), .A(D9576_Q));
KC_NOR2_X1 D9533 ( .Y(D9533_Y), .B(D1988_Y), .A(D9579_Q));
KC_NOR2_X1 D9532 ( .Y(D9532_Y), .B(D1897_Y), .A(D1984_Y));
KC_NOR2_X1 D9530 ( .Y(D9530_Y), .B(D9394_Y), .A(D8105_Y));
KC_NOR2_X1 D9526 ( .Y(D9526_Y), .B(D9547_Y), .A(D9574_Q));
KC_NOR2_X1 D9519 ( .Y(D9519_Y), .B(D9398_Y), .A(D9558_Y));
KC_NOR2_X1 D9507 ( .Y(D9507_Y), .B(D9527_Y), .A(D9579_Q));
KC_NOR2_X1 D9506 ( .Y(D9506_Y), .B(D9501_Y), .A(D9514_Y));
KC_NOR2_X1 D9491 ( .Y(D9491_Y), .B(D10193_Y), .A(D10194_Y));
KC_NOR2_X1 D9490 ( .Y(D9490_Y), .B(D9418_Y), .A(D9491_Y));
KC_NOR2_X1 D9487 ( .Y(D9487_Y), .B(D9411_Y), .A(D9410_Y));
KC_NOR2_X1 D9486 ( .Y(D9486_Y), .B(D2063_Y), .A(D9487_Y));
KC_NOR2_X1 D9408 ( .Y(D9408_Y), .B(D9484_Y), .A(D9463_Y));
KC_NOR2_X1 D9402 ( .Y(D9402_Y), .B(D8079_Y), .A(D8221_Y));
KC_NOR2_X1 D9390 ( .Y(D9390_Y), .B(D622_Y), .A(D9405_Y));
KC_NOR2_X1 D9368 ( .Y(D9368_Y), .B(D2042_Y), .A(D6288_Y));
KC_NOR2_X1 D9237 ( .Y(D9237_Y), .B(D2001_Y), .A(D417_Y));
KC_NOR2_X1 D9191 ( .Y(D9191_Y), .B(D9101_Y), .A(D1711_Y));
KC_NOR2_X1 D9187 ( .Y(D9187_Y), .B(D7683_Y), .A(D1711_Y));
KC_NOR2_X1 D9182 ( .Y(D9182_Y), .B(D9180_Y), .A(D1711_Y));
KC_NOR2_X1 D9179 ( .Y(D9179_Y), .B(D382_Y), .A(D9268_Y));
KC_NOR2_X1 D9174 ( .Y(D9174_Y), .B(D9215_Q), .A(D421_Q));
KC_NOR2_X1 D9117 ( .Y(D9117_Y), .B(D2099_Y), .A(D7500_Y));
KC_NOR2_X1 D9112 ( .Y(D9112_Y), .B(D9113_Y), .A(D1904_Y));
KC_NOR2_X1 D9111 ( .Y(D9111_Y), .B(D2099_Y), .A(D9057_Y));
KC_NOR2_X1 D9106 ( .Y(D9106_Y), .B(D2099_Y), .A(D338_Y));
KC_NOR2_X1 D9104 ( .Y(D9104_Y), .B(D10068_Y), .A(D374_Y));
KC_NOR2_X1 D9068 ( .Y(D9068_Y), .B(D5705_Y), .A(D1711_Y));
KC_NOR2_X1 D9054 ( .Y(D9054_Y), .B(D5705_Y), .A(D7500_Y));
KC_NOR2_X1 D9029 ( .Y(D9029_Y), .B(D9145_Y), .A(D2077_Y));
KC_NOR2_X1 D9028 ( .Y(D9028_Y), .B(D9007_Y), .A(D320_Y));
KC_NOR2_X1 D8974 ( .Y(D8974_Y), .B(D8970_Y), .A(D7361_Y));
KC_NOR2_X1 D8969 ( .Y(D8969_Y), .B(D9064_Y), .A(D7361_Y));
KC_NOR2_X1 D8876 ( .Y(D8876_Y), .B(D9481_Y), .A(D2095_Y));
KC_NOR2_X1 D8874 ( .Y(D8874_Y), .B(D8864_Y), .A(D8899_Q));
KC_NOR2_X1 D8869 ( .Y(D8869_Y), .B(D8860_Y), .A(D8898_Q));
KC_NOR2_X1 D8859 ( .Y(D8859_Y), .B(D8919_Y), .A(D8824_Q));
KC_NOR2_X1 D8762 ( .Y(D8762_Y), .B(D215_Y), .A(D7460_Y));
KC_NOR2_X1 D8750 ( .Y(D8750_Y), .B(D8791_Y), .A(D2028_Y));
KC_NOR2_X1 D8747 ( .Y(D8747_Y), .B(D8877_Y), .A(D8748_Y));
KC_NOR2_X1 D8746 ( .Y(D8746_Y), .B(D5725_Y), .A(D8815_Y));
KC_NOR2_X1 D8745 ( .Y(D8745_Y), .B(D5725_Y), .A(D2160_Y));
KC_NOR2_X1 D8741 ( .Y(D8741_Y), .B(D8744_Y), .A(D9479_Y));
KC_NOR2_X1 D8735 ( .Y(D8735_Y), .B(D5725_Y), .A(D7185_Y));
KC_NOR2_X1 D8677 ( .Y(D8677_Y), .B(D8728_Y), .A(D8674_Y));
KC_NOR2_X1 D8667 ( .Y(D8667_Y), .B(D8769_Y), .A(D9923_Y));
KC_NOR2_X1 D8563 ( .Y(D8563_Y), .B(D8564_Y), .A(D8422_Y));
KC_NOR2_X1 D8495 ( .Y(D8495_Y), .B(D8501_Y), .A(D8422_Y));
KC_NOR2_X1 D8491 ( .Y(D8491_Y), .B(D8493_Y), .A(D8422_Y));
KC_NOR2_X1 D8490 ( .Y(D8490_Y), .B(D8494_Y), .A(D8422_Y));
KC_NOR2_X1 D8489 ( .Y(D8489_Y), .B(D8492_Y), .A(D8422_Y));
KC_NOR2_X1 D8486 ( .Y(D8486_Y), .B(D8488_Y), .A(D8422_Y));
KC_NOR2_X1 D8483 ( .Y(D8483_Y), .B(D8482_Y), .A(D8422_Y));
KC_NOR2_X1 D8480 ( .Y(D8480_Y), .B(D8481_Y), .A(D8422_Y));
KC_NOR2_X1 D8479 ( .Y(D8479_Y), .B(D1832_Y), .A(D8422_Y));
KC_NOR2_X1 D8418 ( .Y(D8418_Y), .B(D9369_Y), .A(D7668_Y));
KC_NOR2_X1 D8415 ( .Y(D8415_Y), .B(D8018_Y), .A(D2353_Y));
KC_NOR2_X1 D8410 ( .Y(D8410_Y), .B(D1993_Y), .A(D2343_Y));
KC_NOR2_X1 D8401 ( .Y(D8401_Y), .B(D9369_Y), .A(D2343_Y));
KC_NOR2_X1 D8400 ( .Y(D8400_Y), .B(D8405_Y), .A(D8388_Y));
KC_NOR2_X1 D8384 ( .Y(D8384_Y), .B(D8368_Y), .A(D8387_Y));
KC_NOR2_X1 D8383 ( .Y(D8383_Y), .B(D8419_Y), .A(D8388_Y));
KC_NOR2_X1 D8382 ( .Y(D8382_Y), .B(D8414_Y), .A(D8405_Y));
KC_NOR2_X1 D8381 ( .Y(D8381_Y), .B(D8392_Y), .A(D6787_Y));
KC_NOR2_X1 D8376 ( .Y(D8376_Y), .B(D8504_Y), .A(D8395_Y));
KC_NOR2_X1 D8372 ( .Y(D8372_Y), .B(D9643_Y), .A(D8365_Y));
KC_NOR2_X1 D8367 ( .Y(D8367_Y), .B(D8366_Y), .A(D8365_Y));
KC_NOR2_X1 D8286 ( .Y(D8286_Y), .B(D1993_Y), .A(D7668_Y));
KC_NOR2_X1 D8279 ( .Y(D8279_Y), .B(D8018_Y), .A(D7669_Y));
KC_NOR2_X1 D8278 ( .Y(D8278_Y), .B(D8350_Y), .A(D8048_Y));
KC_NOR2_X1 D8266 ( .Y(D8266_Y), .B(D8175_Y), .A(D854_Y));
KC_NOR2_X1 D8202 ( .Y(D8202_Y), .B(D8249_Q), .A(D8247_Q));
KC_NOR2_X1 D8201 ( .Y(D8201_Y), .B(D8250_Q), .A(D8248_Q));
KC_NOR2_X1 D8184 ( .Y(D8184_Y), .B(D8199_Y), .A(D8186_Y));
KC_NOR2_X1 D8177 ( .Y(D8177_Y), .B(D8186_Y), .A(D7974_Y));
KC_NOR2_X1 D8111 ( .Y(D8111_Y), .B(D9390_Y), .A(D8120_Y));
KC_NOR2_X1 D8108 ( .Y(D8108_Y), .B(D8117_Y), .A(D9551_Y));
KC_NOR2_X1 D8107 ( .Y(D8107_Y), .B(D8098_Y), .A(D8105_Y));
KC_NOR2_X1 D8106 ( .Y(D8106_Y), .B(D9437_Y), .A(D8108_Y));
KC_NOR2_X1 D8105 ( .Y(D8105_Y), .B(D8109_Y), .A(D4137_Q));
KC_NOR2_X1 D8099 ( .Y(D8099_Y), .B(D8077_Y), .A(D8221_Y));
KC_NOR2_X1 D8098 ( .Y(D8098_Y), .B(D8115_Y), .A(D9407_Y));
KC_NOR2_X1 D8087 ( .Y(D8087_Y), .B(D8083_Y), .A(D8079_Y));
KC_NOR2_X1 D8086 ( .Y(D8086_Y), .B(D8088_Y), .A(D8138_Y));
KC_NOR2_X1 D8078 ( .Y(D8078_Y), .B(D8120_Y), .A(D8093_Y));
KC_NOR2_X1 D8077 ( .Y(D8077_Y), .B(D8194_Y), .A(D8201_Y));
KC_NOR2_X1 D8076 ( .Y(D8076_Y), .B(D8147_Q), .A(D7478_Q));
KC_NOR2_X1 D8019 ( .Y(D8019_Y), .B(D8044_Y), .A(D620_Y));
KC_NOR2_X1 D8013 ( .Y(D8013_Y), .B(D8015_Y), .A(D8016_Y));
KC_NOR2_X1 D8005 ( .Y(D8005_Y), .B(D8121_Y), .A(D8007_Y));
KC_NOR2_X1 D8001 ( .Y(D8001_Y), .B(D9363_Y), .A(D9372_Y));
KC_NOR2_X1 D7986 ( .Y(D7986_Y), .B(D7925_Y), .A(D7946_Y));
KC_NOR2_X1 D7948 ( .Y(D7948_Y), .B(D1940_Q), .A(D7949_Y));
KC_NOR2_X1 D7945 ( .Y(D7945_Y), .B(D7932_Y), .A(D7936_Y));
KC_NOR2_X1 D7944 ( .Y(D7944_Y), .B(D7936_Y), .A(D7933_Y));
KC_NOR2_X1 D7943 ( .Y(D7943_Y), .B(D7946_Y), .A(D7924_Y));
KC_NOR2_X1 D7942 ( .Y(D7942_Y), .B(D152_Q), .A(D1940_Q));
KC_NOR2_X1 D7936 ( .Y(D7936_Y), .B(D7946_Y), .A(D7923_Y));
KC_NOR2_X1 D7935 ( .Y(D7935_Y), .B(D7937_Y), .A(D7923_Y));
KC_NOR2_X1 D7934 ( .Y(D7934_Y), .B(D7986_Y), .A(D1852_Y));
KC_NOR2_X1 D7933 ( .Y(D7933_Y), .B(D7925_Y), .A(D7938_Y));
KC_NOR2_X1 D7932 ( .Y(D7932_Y), .B(D7924_Y), .A(D7937_Y));
KC_NOR2_X1 D7929 ( .Y(D7929_Y), .B(D7938_Y), .A(D7923_Y));
KC_NOR2_X1 D7921 ( .Y(D7921_Y), .B(D7924_Y), .A(D7938_Y));
KC_NOR2_X1 D7920 ( .Y(D7920_Y), .B(D7922_Y), .A(D7937_Y));
KC_NOR2_X1 D7919 ( .Y(D7919_Y), .B(D7925_Y), .A(D7937_Y));
KC_NOR2_X1 D7916 ( .Y(D7916_Y), .B(D7937_Y), .A(D7917_Y));
KC_NOR2_X1 D7915 ( .Y(D7915_Y), .B(D7922_Y), .A(D7938_Y));
KC_NOR2_X1 D7912 ( .Y(D7912_Y), .B(D7975_Y), .A(D7837_Y));
KC_NOR2_X1 D7911 ( .Y(D7911_Y), .B(D7922_Y), .A(D7937_Y));
KC_NOR2_X1 D7857 ( .Y(D7857_Y), .B(D7859_Y), .A(D7885_Q));
KC_NOR2_X1 D7855 ( .Y(D7855_Y), .B(D7852_Y), .A(D7883_Q));
KC_NOR2_X1 D7851 ( .Y(D7851_Y), .B(D7580_Y), .A(D7887_Q));
KC_NOR2_X1 D7846 ( .Y(D7846_Y), .B(D7886_Q), .A(D480_Q));
KC_NOR2_X1 D7845 ( .Y(D7845_Y), .B(D7854_Y), .A(D7889_Q));
KC_NOR2_X1 D7841 ( .Y(D7841_Y), .B(D7829_Y), .A(D7888_Q));
KC_NOR2_X1 D7828 ( .Y(D7828_Y), .B(D7831_Y), .A(D7839_Y));
KC_NOR2_X1 D7827 ( .Y(D7827_Y), .B(D7955_Y), .A(D7925_Y));
KC_NOR2_X1 D7769 ( .Y(D7769_Y), .B(D7766_Y), .A(D272_Y));
KC_NOR2_X1 D7766 ( .Y(D7766_Y), .B(D7765_Y), .A(D10154_Y));
KC_NOR2_X1 D7761 ( .Y(D7761_Y), .B(D7796_Y), .A(D7804_Y));
KC_NOR2_X1 D7692 ( .Y(D7692_Y), .B(D10142_Y), .A(D346_Y));
KC_NOR2_X1 D7691 ( .Y(D7691_Y), .B(D10142_Y), .A(D7563_Y));
KC_NOR2_X1 D7690 ( .Y(D7690_Y), .B(D7784_Y), .A(D346_Y));
KC_NOR2_X1 D7689 ( .Y(D7689_Y), .B(D7784_Y), .A(D723_Q));
KC_NOR2_X1 D7686 ( .Y(D7686_Y), .B(D9268_Y), .A(D7564_Y));
KC_NOR2_X1 D7682 ( .Y(D7682_Y), .B(D9354_Y), .A(D7564_Y));
KC_NOR2_X1 D7678 ( .Y(D7678_Y), .B(D13288_Y), .A(D481_Y));
KC_NOR2_X1 D7677 ( .Y(D7677_Y), .B(D7679_Y), .A(D7676_Y));
KC_NOR2_X1 D7638 ( .Y(D7638_Y), .B(D6097_Y), .A(D1713_Y));
KC_NOR2_X1 D7636 ( .Y(D7636_Y), .B(D10162_Y), .A(D7564_Y));
KC_NOR2_X1 D7631 ( .Y(D7631_Y), .B(D6096_Y), .A(D1787_Y));
KC_NOR2_X1 D7630 ( .Y(D7630_Y), .B(D9354_Y), .A(D7563_Y));
KC_NOR2_X1 D7628 ( .Y(D7628_Y), .B(D7713_Y), .A(D7564_Y));
KC_NOR2_X1 D7627 ( .Y(D7627_Y), .B(D10142_Y), .A(D7564_Y));
KC_NOR2_X1 D7626 ( .Y(D7626_Y), .B(D10159_Y), .A(D346_Y));
KC_NOR2_X1 D7625 ( .Y(D7625_Y), .B(D7648_Y), .A(D6250_Y));
KC_NOR2_X1 D7623 ( .Y(D7623_Y), .B(D9268_Y), .A(D7563_Y));
KC_NOR2_X1 D7562 ( .Y(D7562_Y), .B(D7587_Q), .A(D7586_Q));
KC_NOR2_X1 D7561 ( .Y(D7561_Y), .B(D10159_Y), .A(D7564_Y));
KC_NOR2_X1 D7558 ( .Y(D7558_Y), .B(D7730_Y), .A(D7563_Y));
KC_NOR2_X1 D7557 ( .Y(D7557_Y), .B(D9269_Y), .A(D346_Y));
KC_NOR2_X1 D7556 ( .Y(D7556_Y), .B(D7730_Y), .A(D346_Y));
KC_NOR2_X1 D7554 ( .Y(D7554_Y), .B(D10159_Y), .A(D7563_Y));
KC_NOR2_X1 D7553 ( .Y(D7553_Y), .B(D10160_Y), .A(D7564_Y));
KC_NOR2_X1 D7550 ( .Y(D7550_Y), .B(D9354_Y), .A(D346_Y));
KC_NOR2_X1 D7549 ( .Y(D7549_Y), .B(D9269_Y), .A(D7564_Y));
KC_NOR2_X1 D7548 ( .Y(D7548_Y), .B(D10160_Y), .A(D346_Y));
KC_NOR2_X1 D7547 ( .Y(D7547_Y), .B(D10160_Y), .A(D7563_Y));
KC_NOR2_X1 D7543 ( .Y(D7543_Y), .B(D7615_Q), .A(D7614_Q));
KC_NOR2_X1 D7499 ( .Y(D7499_Y), .B(D6097_Y), .A(D8838_Y));
KC_NOR2_X1 D7494 ( .Y(D7494_Y), .B(D5705_Y), .A(D7503_Y));
KC_NOR2_X1 D10 ( .Y(D10_Y), .B(D7480_Q), .A(D9473_Y));
KC_NOR2_X1 D9 ( .Y(D9_Y), .B(D6061_Y), .A(D10_Y));
KC_NOR2_X1 D7439 ( .Y(D7439_Y), .B(D7318_Y), .A(D7164_Y));
KC_NOR2_X1 D7438 ( .Y(D7438_Y), .B(D5828_Y), .A(D6045_Y));
KC_NOR2_X1 D7434 ( .Y(D7434_Y), .B(D7451_Y), .A(D7361_Y));
KC_NOR2_X1 D7426 ( .Y(D7426_Y), .B(D6073_Q), .A(D8153_Y));
KC_NOR2_X1 D7423 ( .Y(D7423_Y), .B(D5998_Y), .A(D7465_Y));
KC_NOR2_X1 D7422 ( .Y(D7422_Y), .B(D6003_Y), .A(D7480_Q));
KC_NOR2_X1 D7418 ( .Y(D7418_Y), .B(D5961_Y), .A(D7296_Y));
KC_NOR2_X1 D7417 ( .Y(D7417_Y), .B(D7505_Y), .A(D5826_Y));
KC_NOR2_X1 D7357 ( .Y(D7357_Y), .B(D1908_Y), .A(D7406_Y));
KC_NOR2_X1 D7356 ( .Y(D7356_Y), .B(D5846_Y), .A(D5703_Y));
KC_NOR2_X1 D7349 ( .Y(D7349_Y), .B(D7215_Y), .A(D7199_Y));
KC_NOR2_X1 D7348 ( .Y(D7348_Y), .B(D214_Y), .A(D4444_Y));
KC_NOR2_X1 D7347 ( .Y(D7347_Y), .B(D7215_Y), .A(D7319_Y));
KC_NOR2_X1 D7345 ( .Y(D7345_Y), .B(D5825_Y), .A(D7460_Y));
KC_NOR2_X1 D7342 ( .Y(D7342_Y), .B(D5647_Y), .A(D7376_Y));
KC_NOR2_X1 D7333 ( .Y(D7333_Y), .B(D4448_Y), .A(D214_Y));
KC_NOR2_X1 D7326 ( .Y(D7326_Y), .B(D7233_Y), .A(D7263_Y));
KC_NOR2_X1 D7325 ( .Y(D7325_Y), .B(D1877_Y), .A(D5851_Y));
KC_NOR2_X1 D7322 ( .Y(D7322_Y), .B(D7355_Y), .A(D7433_Y));
KC_NOR2_X1 D7320 ( .Y(D7320_Y), .B(D272_Y), .A(D7_Y));
KC_NOR2_X1 D7315 ( .Y(D7315_Y), .B(D5703_Y), .A(D7361_Y));
KC_NOR2_X1 D7314 ( .Y(D7314_Y), .B(D5677_Y), .A(D5698_Y));
KC_NOR2_X1 D7313 ( .Y(D7313_Y), .B(D7314_Y), .A(D7460_Y));
KC_NOR2_X1 D7304 ( .Y(D7304_Y), .B(D7248_Y), .A(D7303_Y));
KC_NOR2_X1 D7257 ( .Y(D7257_Y), .B(D6333_Y), .A(D7101_Y));
KC_NOR2_X1 D7256 ( .Y(D7256_Y), .B(D6333_Y), .A(D7141_Y));
KC_NOR2_X1 D7255 ( .Y(D7255_Y), .B(D7260_Y), .A(D7140_Y));
KC_NOR2_X1 D7254 ( .Y(D7254_Y), .B(D7104_Y), .A(D6334_Y));
KC_NOR2_X1 D7251 ( .Y(D7251_Y), .B(D2027_Y), .A(D8756_Y));
KC_NOR2_X1 D7243 ( .Y(D7243_Y), .B(D7279_Y), .A(D7104_Y));
KC_NOR2_X1 D7242 ( .Y(D7242_Y), .B(D6470_Y), .A(D7140_Y));
KC_NOR2_X1 D7241 ( .Y(D7241_Y), .B(D6334_Y), .A(D7097_Y));
KC_NOR2_X1 D7234 ( .Y(D7234_Y), .B(D7303_Y), .A(D7152_Q));
KC_NOR2_X1 D7233 ( .Y(D7233_Y), .B(D7247_Y), .A(D7253_Y));
KC_NOR2_X1 D7232 ( .Y(D7232_Y), .B(D7247_Y), .A(D7273_Y));
KC_NOR2_X1 D7210 ( .Y(D7210_Y), .B(D7252_Y), .A(D7246_Y));
KC_NOR2_X1 D7209 ( .Y(D7209_Y), .B(D1887_Y), .A(D9479_Y));
KC_NOR2_X1 D7205 ( .Y(D7205_Y), .B(D7218_Y), .A(D220_Y));
KC_NOR2_X1 D7195 ( .Y(D7195_Y), .B(D7203_Y), .A(D8776_Y));
KC_NOR2_X1 D7194 ( .Y(D7194_Y), .B(D7172_Y), .A(D7212_Y));
KC_NOR2_X1 D7193 ( .Y(D7193_Y), .B(D5647_Y), .A(D1740_Y));
KC_NOR2_X1 D7192 ( .Y(D7192_Y), .B(D2053_Y), .A(D7203_Y));
KC_NOR2_X1 D7177 ( .Y(D7177_Y), .B(D7250_Y), .A(D7253_Y));
KC_NOR2_X1 D7167 ( .Y(D7167_Y), .B(D7180_Y), .A(D9481_Y));
KC_NOR2_X1 D7166 ( .Y(D7166_Y), .B(D7172_Y), .A(D7167_Y));
KC_NOR2_X1 D7116 ( .Y(D7116_Y), .B(D7144_Q), .A(D7146_Q));
KC_NOR2_X1 D7114 ( .Y(D7114_Y), .B(D8706_Y), .A(D5682_Y));
KC_NOR2_X1 D7110 ( .Y(D7110_Y), .B(D7111_Y), .A(D7112_Y));
KC_NOR2_X1 D7108 ( .Y(D7108_Y), .B(D7124_Y), .A(D5672_Y));
KC_NOR2_X1 D7093 ( .Y(D7093_Y), .B(D7137_Y), .A(D7106_Y));
KC_NOR2_X1 D7092 ( .Y(D7092_Y), .B(D7099_Y), .A(D189_Y));
KC_NOR2_X1 D6991 ( .Y(D6991_Y), .B(D6944_Y), .A(D6935_Y));
KC_NOR2_X1 D6937 ( .Y(D6937_Y), .B(D6936_Y), .A(D8395_Y));
KC_NOR2_X1 D6930 ( .Y(D6930_Y), .B(D8542_Y), .A(D1743_Y));
KC_NOR2_X1 D6926 ( .Y(D6926_Y), .B(D6925_Y), .A(D8395_Y));
KC_NOR2_X1 D6921 ( .Y(D6921_Y), .B(D6944_Y), .A(D6923_Y));
KC_NOR2_X1 D6920 ( .Y(D6920_Y), .B(D6922_Y), .A(D8395_Y));
KC_NOR2_X1 D6919 ( .Y(D6919_Y), .B(D6938_Y), .A(D8542_Y));
KC_NOR2_X1 D6915 ( .Y(D6915_Y), .B(D6942_Y), .A(D6935_Y));
KC_NOR2_X1 D6869 ( .Y(D6869_Y), .B(D992_Y), .A(D6854_Y));
KC_NOR2_X1 D6868 ( .Y(D6868_Y), .B(D992_Y), .A(D6855_Y));
KC_NOR2_X1 D6863 ( .Y(D6863_Y), .B(D6881_Y), .A(D6854_Y));
KC_NOR2_X1 D6862 ( .Y(D6862_Y), .B(D5451_Y), .A(D5442_Y));
KC_NOR2_X1 D6861 ( .Y(D6861_Y), .B(D6881_Y), .A(D6855_Y));
KC_NOR2_X1 D6860 ( .Y(D6860_Y), .B(D6882_Y), .A(D6855_Y));
KC_NOR2_X1 D6856 ( .Y(D6856_Y), .B(D1846_Y), .A(D813_Y));
KC_NOR2_X1 D6853 ( .Y(D6853_Y), .B(D6882_Y), .A(D6854_Y));
KC_NOR2_X1 D6789 ( .Y(D6789_Y), .B(D1824_Y), .A(D1932_Y));
KC_NOR2_X1 D6785 ( .Y(D6785_Y), .B(D6766_Y), .A(D1932_Y));
KC_NOR2_X1 D6695 ( .Y(D6695_Y), .B(D5294_Y), .A(D5267_Y));
KC_NOR2_X1 D6689 ( .Y(D6689_Y), .B(D1598_Y), .A(D5260_Y));
KC_NOR2_X1 D6515 ( .Y(D6515_Y), .B(D6519_Y), .A(D6512_Y));
KC_NOR2_X1 D6514 ( .Y(D6514_Y), .B(D1694_Y), .A(D1786_Q));
KC_NOR2_X1 D6513 ( .Y(D6513_Y), .B(D6553_Q), .A(D6554_Q));
KC_NOR2_X1 D6511 ( .Y(D6511_Y), .B(D6514_Y), .A(D6555_Q));
KC_NOR2_X1 D6446 ( .Y(D6446_Y), .B(D3408_Y), .A(D1415_Y));
KC_NOR2_X1 D6445 ( .Y(D6445_Y), .B(D4889_Y), .A(D4865_Y));
KC_NOR2_X1 D6444 ( .Y(D6444_Y), .B(D6481_Q), .A(D485_Q));
KC_NOR2_X1 D6441 ( .Y(D6441_Y), .B(D7856_Y), .A(D479_Q));
KC_NOR2_X1 D6436 ( .Y(D6436_Y), .B(D6437_Y), .A(D6464_Y));
KC_NOR2_X1 D6432 ( .Y(D6432_Y), .B(D3647_Q), .A(D6491_Q));
KC_NOR2_X1 D6431 ( .Y(D6431_Y), .B(D6491_Q), .A(D6486_Q));
KC_NOR2_X1 D6426 ( .Y(D6426_Y), .B(D6427_Y), .A(D6431_Y));
KC_NOR2_X1 D6421 ( .Y(D6421_Y), .B(D5031_Y), .A(D4865_Y));
KC_NOR2_X1 D6420 ( .Y(D6420_Y), .B(D7918_Y), .A(D7935_Y));
KC_NOR2_X1 D6367 ( .Y(D6367_Y), .B(D6365_Y), .A(D446_Q));
KC_NOR2_X1 D6365 ( .Y(D6365_Y), .B(D441_Y), .A(D445_Q));
KC_NOR2_X1 D6364 ( .Y(D6364_Y), .B(D6411_Y), .A(D4951_Y));
KC_NOR2_X1 D6308 ( .Y(D6308_Y), .B(D10158_Y), .A(D346_Y));
KC_NOR2_X1 D6307 ( .Y(D6307_Y), .B(D7713_Y), .A(D346_Y));
KC_NOR2_X1 D6306 ( .Y(D6306_Y), .B(D10158_Y), .A(D7563_Y));
KC_NOR2_X1 D6305 ( .Y(D6305_Y), .B(D10161_Y), .A(D7563_Y));
KC_NOR2_X1 D6304 ( .Y(D6304_Y), .B(D7784_Y), .A(D7563_Y));
KC_NOR2_X1 D6303 ( .Y(D6303_Y), .B(D6302_Y), .A(D6354_Y));
KC_NOR2_X1 D6302 ( .Y(D6302_Y), .B(D6354_Y), .A(D6330_Y));
KC_NOR2_X1 D6301 ( .Y(D6301_Y), .B(D7713_Y), .A(D7563_Y));
KC_NOR2_X1 D6297 ( .Y(D6297_Y), .B(D10161_Y), .A(D7564_Y));
KC_NOR2_X1 D6296 ( .Y(D6296_Y), .B(D10158_Y), .A(D7564_Y));
KC_NOR2_X1 D6232 ( .Y(D6232_Y), .B(D481_Y), .A(D7564_Y));
KC_NOR2_X1 D6230 ( .Y(D6230_Y), .B(D9266_Y), .A(D7563_Y));
KC_NOR2_X1 D6225 ( .Y(D6225_Y), .B(D7784_Y), .A(D7564_Y));
KC_NOR2_X1 D6220 ( .Y(D6220_Y), .B(D6241_Y), .A(D6249_Y));
KC_NOR2_X1 D6216 ( .Y(D6216_Y), .B(D6211_Y), .A(D1945_Y));
KC_NOR2_X1 D6210 ( .Y(D6210_Y), .B(D10161_Y), .A(D346_Y));
KC_NOR2_X1 D6144 ( .Y(D6144_Y), .B(D7730_Y), .A(D7564_Y));
KC_NOR2_X1 D6143 ( .Y(D6143_Y), .B(D10157_Y), .A(D7563_Y));
KC_NOR2_X1 D6142 ( .Y(D6142_Y), .B(D10157_Y), .A(D346_Y));
KC_NOR2_X1 D6141 ( .Y(D6141_Y), .B(D10157_Y), .A(D7564_Y));
KC_NOR2_X1 D6140 ( .Y(D6140_Y), .B(D9266_Y), .A(D7564_Y));
KC_NOR2_X1 D6139 ( .Y(D6139_Y), .B(D7785_Y), .A(D346_Y));
KC_NOR2_X1 D6137 ( .Y(D6137_Y), .B(D9269_Y), .A(D7563_Y));
KC_NOR2_X1 D6136 ( .Y(D6136_Y), .B(D10162_Y), .A(D346_Y));
KC_NOR2_X1 D6135 ( .Y(D6135_Y), .B(D9266_Y), .A(D346_Y));
KC_NOR2_X1 D6133 ( .Y(D6133_Y), .B(D6154_Y), .A(D6134_Y));
KC_NOR2_X1 D6095 ( .Y(D6095_Y), .B(D5990_Y), .A(D7629_Y));
KC_NOR2_X1 D6090 ( .Y(D6090_Y), .B(D1787_Y), .A(D1713_Y));
KC_NOR2_X1 D6033 ( .Y(D6033_Y), .B(D5685_Y), .A(D1872_Y));
KC_NOR2_X1 D6032 ( .Y(D6032_Y), .B(D7305_Y), .A(D6037_Y));
KC_NOR2_X1 D6028 ( .Y(D6028_Y), .B(D6037_Y), .A(D203_Y));
KC_NOR2_X1 D6020 ( .Y(D6020_Y), .B(D4437_Y), .A(D4439_Y));
KC_NOR2_X1 D6019 ( .Y(D6019_Y), .B(D5872_Y), .A(D5877_Y));
KC_NOR2_X1 D6018 ( .Y(D6018_Y), .B(D5950_Y), .A(D6022_Y));
KC_NOR2_X1 D6014 ( .Y(D6014_Y), .B(D287_Y), .A(D7480_Q));
KC_NOR2_X1 D6008 ( .Y(D6008_Y), .B(D5745_Y), .A(D6010_Y));
KC_NOR2_X1 D6007 ( .Y(D6007_Y), .B(D5999_Y), .A(D4425_Y));
KC_NOR2_X1 D6006 ( .Y(D6006_Y), .B(D6048_Y), .A(D213_Y));
KC_NOR2_X1 D6003 ( .Y(D6003_Y), .B(D6039_Y), .A(D5646_Y));
KC_NOR2_X1 D6000 ( .Y(D6000_Y), .B(D4415_Y), .A(D5973_Y));
KC_NOR2_X1 D5984 ( .Y(D5984_Y), .B(D4410_Y), .A(D6097_Y));
KC_NOR2_X1 D5983 ( .Y(D5983_Y), .B(D5973_Y), .A(D6113_Y));
KC_NOR2_X1 D5982 ( .Y(D5982_Y), .B(D5971_Y), .A(D5981_Y));
KC_NOR2_X1 D5981 ( .Y(D5981_Y), .B(D4419_Y), .A(D290_Y));
KC_NOR2_X1 D5980 ( .Y(D5980_Y), .B(D4410_Y), .A(D6044_Y));
KC_NOR2_X1 D5971 ( .Y(D5971_Y), .B(D5974_Y), .A(D4410_Y));
KC_NOR2_X1 D5970 ( .Y(D5970_Y), .B(D5975_Y), .A(D4409_Y));
KC_NOR2_X1 D5969 ( .Y(D5969_Y), .B(D5973_Y), .A(D1713_Y));
KC_NOR2_X1 D5968 ( .Y(D5968_Y), .B(D6041_Y), .A(D1872_Y));
KC_NOR2_X1 D5967 ( .Y(D5967_Y), .B(D6075_Y), .A(D7469_Y));
KC_NOR2_X1 D5962 ( .Y(D5962_Y), .B(D165_Y), .A(D5958_Y));
KC_NOR2_X1 D5954 ( .Y(D5954_Y), .B(D4405_Y), .A(D239_Q));
KC_NOR2_X1 D5953 ( .Y(D5953_Y), .B(D4413_Y), .A(D5958_Y));
KC_NOR2_X1 D5952 ( .Y(D5952_Y), .B(D5805_Y), .A(D6108_Y));
KC_NOR2_X1 D5882 ( .Y(D5882_Y), .B(D7419_Y), .A(D4350_Y));
KC_NOR2_X1 D5881 ( .Y(D5881_Y), .B(D5876_Y), .A(D5856_Y));
KC_NOR2_X1 D5880 ( .Y(D5880_Y), .B(D7334_Y), .A(D4488_Q));
KC_NOR2_X1 D5872 ( .Y(D5872_Y), .B(D1592_Y), .A(D5756_Y));
KC_NOR2_X1 D5871 ( .Y(D5871_Y), .B(D4349_Y), .A(D5756_Y));
KC_NOR2_X1 D5870 ( .Y(D5870_Y), .B(D5874_Y), .A(D5867_Y));
KC_NOR2_X1 D5869 ( .Y(D5869_Y), .B(D7246_Y), .A(D5651_Y));
KC_NOR2_X1 D5863 ( .Y(D5863_Y), .B(D5867_Y), .A(D7376_Y));
KC_NOR2_X1 D5859 ( .Y(D5859_Y), .B(D1723_Y), .A(D247_Y));
KC_NOR2_X1 D5856 ( .Y(D5856_Y), .B(D1612_Y), .A(D5973_Y));
KC_NOR2_X1 D5839 ( .Y(D5839_Y), .B(D5896_Y), .A(D5838_Y));
KC_NOR2_X1 D5838 ( .Y(D5838_Y), .B(D4448_Y), .A(D5857_Y));
KC_NOR2_X1 D5837 ( .Y(D5837_Y), .B(D5888_Y), .A(D6001_Y));
KC_NOR2_X1 D5835 ( .Y(D5835_Y), .B(D7319_Y), .A(D5857_Y));
KC_NOR2_X1 D5833 ( .Y(D5833_Y), .B(D5830_Y), .A(D7376_Y));
KC_NOR2_X1 D5827 ( .Y(D5827_Y), .B(D4285_Y), .A(D7376_Y));
KC_NOR2_X1 D5760 ( .Y(D5760_Y), .B(D5847_Y), .A(D5763_Y));
KC_NOR2_X1 D5752 ( .Y(D5752_Y), .B(D6024_Y), .A(D5685_Y));
KC_NOR2_X1 D5751 ( .Y(D5751_Y), .B(D5741_Y), .A(D7263_Y));
KC_NOR2_X1 D5742 ( .Y(D5742_Y), .B(D5883_Y), .A(D5684_Y));
KC_NOR2_X1 D5741 ( .Y(D5741_Y), .B(D5746_Y), .A(D213_Y));
KC_NOR2_X1 D5737 ( .Y(D5737_Y), .B(D7500_Y), .A(D1736_Y));
KC_NOR2_X1 D5736 ( .Y(D5736_Y), .B(D6072_Y), .A(D1739_Y));
KC_NOR2_X1 D5726 ( .Y(D5726_Y), .B(D5722_Y), .A(D4136_Q));
KC_NOR2_X1 D5714 ( .Y(D5714_Y), .B(D5729_Y), .A(D14_Y));
KC_NOR2_X1 D5667 ( .Y(D5667_Y), .B(D5669_Y), .A(D5689_Q));
KC_NOR2_X1 D5666 ( .Y(D5666_Y), .B(D5686_Q), .A(D5690_Q));
KC_NOR2_X1 D5660 ( .Y(D5660_Y), .B(D5689_Q), .A(D5687_Q));
KC_NOR2_X1 D5657 ( .Y(D5657_Y), .B(D5655_Y), .A(D5688_Q));
KC_NOR2_X1 D5653 ( .Y(D5653_Y), .B(D5691_Q), .A(D5655_Y));
KC_NOR2_X1 D5652 ( .Y(D5652_Y), .B(D5668_Y), .A(D5664_Y));
KC_NOR2_X1 D5646 ( .Y(D5646_Y), .B(D5663_Y), .A(D5676_Y));
KC_NOR2_X1 D5645 ( .Y(D5645_Y), .B(D7266_Y), .A(D7376_Y));
KC_NOR2_X1 D5644 ( .Y(D5644_Y), .B(D5654_Y), .A(D5676_Y));
KC_NOR2_X1 D5543 ( .Y(D5543_Y), .B(D5523_Y), .A(D5520_Y));
KC_NOR2_X1 D5509 ( .Y(D5509_Y), .B(D5523_Y), .A(D5510_Y));
KC_NOR2_X1 D5498 ( .Y(D5498_Y), .B(D5521_Y), .A(D5510_Y));
KC_NOR2_X1 D5497 ( .Y(D5497_Y), .B(D5521_Y), .A(D5520_Y));
KC_NOR2_X1 D5440 ( .Y(D5440_Y), .B(D5452_Y), .A(D5441_Y));
KC_NOR2_X1 D5437 ( .Y(D5437_Y), .B(D5453_Y), .A(D5441_Y));
KC_NOR2_X1 D5436 ( .Y(D5436_Y), .B(D5453_Y), .A(D5442_Y));
KC_NOR2_X1 D5356 ( .Y(D5356_Y), .B(D5375_Y), .A(D5358_Y));
KC_NOR2_X1 D5355 ( .Y(D5355_Y), .B(D5373_Y), .A(D5361_Y));
KC_NOR2_X1 D5354 ( .Y(D5354_Y), .B(D5374_Y), .A(D5361_Y));
KC_NOR2_X1 D5353 ( .Y(D5353_Y), .B(D5374_Y), .A(D5358_Y));
KC_NOR2_X1 D5349 ( .Y(D5349_Y), .B(D5378_Y), .A(D5341_Y));
KC_NOR2_X1 D5348 ( .Y(D5348_Y), .B(D5371_Y), .A(D5341_Y));
KC_NOR2_X1 D5347 ( .Y(D5347_Y), .B(D5371_Y), .A(D5357_Y));
KC_NOR2_X1 D5346 ( .Y(D5346_Y), .B(D5378_Y), .A(D5357_Y));
KC_NOR2_X1 D5345 ( .Y(D5345_Y), .B(D5370_Y), .A(D5357_Y));
KC_NOR2_X1 D5344 ( .Y(D5344_Y), .B(D5373_Y), .A(D5358_Y));
KC_NOR2_X1 D5340 ( .Y(D5340_Y), .B(D5370_Y), .A(D5341_Y));
KC_NOR2_X1 D5266 ( .Y(D5266_Y), .B(D1599_Y), .A(D5267_Y));
KC_NOR2_X1 D5265 ( .Y(D5265_Y), .B(D1599_Y), .A(D5260_Y));
KC_NOR2_X1 D5038 ( .Y(D5038_Y), .B(D4902_Y), .A(D3371_Y));
KC_NOR2_X1 D5037 ( .Y(D5037_Y), .B(D4882_Y), .A(D1537_Y));
KC_NOR2_X1 D5036 ( .Y(D5036_Y), .B(D1570_Y), .A(D3498_Y));
KC_NOR2_X1 D5029 ( .Y(D5029_Y), .B(D4889_Y), .A(D5023_Y));
KC_NOR2_X1 D5028 ( .Y(D5028_Y), .B(D1570_Y), .A(D3499_Y));
KC_NOR2_X1 D5009 ( .Y(D5009_Y), .B(D5020_Y), .A(D4911_Y));
KC_NOR2_X1 D5008 ( .Y(D5008_Y), .B(D5021_Y), .A(D5023_Y));
KC_NOR2_X1 D4996 ( .Y(D4996_Y), .B(D5004_Y), .A(D3599_Y));
KC_NOR2_X1 D4995 ( .Y(D4995_Y), .B(D3420_Y), .A(D4865_Y));
KC_NOR2_X1 D4920 ( .Y(D4920_Y), .B(D3388_Q), .A(D3498_Y));
KC_NOR2_X1 D4913 ( .Y(D4913_Y), .B(D3400_Y), .A(D3388_Q));
KC_NOR2_X1 D4908 ( .Y(D4908_Y), .B(D4926_Y), .A(D3416_Y));
KC_NOR2_X1 D4907 ( .Y(D4907_Y), .B(D3388_Q), .A(D3484_Q));
KC_NOR2_X1 D4906 ( .Y(D4906_Y), .B(D3371_Y), .A(D3499_Y));
KC_NOR2_X1 D4900 ( .Y(D4900_Y), .B(D3599_Y), .A(D1537_Y));
KC_NOR2_X1 D4892 ( .Y(D4892_Y), .B(D7966_Q), .A(D7968_Q));
KC_NOR2_X1 D4891 ( .Y(D4891_Y), .B(D3400_Y), .A(D1537_Y));
KC_NOR2_X1 D4887 ( .Y(D4887_Y), .B(D4925_Y), .A(D3400_Y));
KC_NOR2_X1 D4886 ( .Y(D4886_Y), .B(D3499_Y), .A(D4867_Y));
KC_NOR2_X1 D4885 ( .Y(D4885_Y), .B(D4868_Y), .A(D4926_Y));
KC_NOR2_X1 D4877 ( .Y(D4877_Y), .B(D4922_Y), .A(D3400_Y));
KC_NOR2_X1 D4876 ( .Y(D4876_Y), .B(D4889_Y), .A(D4911_Y));
KC_NOR2_X1 D4875 ( .Y(D4875_Y), .B(D4960_Y), .A(D4925_Y));
KC_NOR2_X1 D4874 ( .Y(D4874_Y), .B(D3498_Y), .A(D3499_Y));
KC_NOR2_X1 D4873 ( .Y(D4873_Y), .B(D4869_Y), .A(D3371_Y));
KC_NOR2_X1 D4872 ( .Y(D4872_Y), .B(D3388_Q), .A(D3499_Y));
KC_NOR2_X1 D4871 ( .Y(D4871_Y), .B(D1567_Y), .A(D3498_Y));
KC_NOR2_X1 D4777 ( .Y(D4777_Y), .B(D3163_Y), .A(D4821_Q));
KC_NOR2_X1 D4776 ( .Y(D4776_Y), .B(D3163_Y), .A(D4822_Q));
KC_NOR2_X1 D4775 ( .Y(D4775_Y), .B(D4776_Y), .A(D4777_Y));
KC_NOR2_X1 D4774 ( .Y(D4774_Y), .B(D3258_Y), .A(D3284_Y));
KC_NOR2_X1 D4766 ( .Y(D4766_Y), .B(D413_Y), .A(D4819_Q));
KC_NOR2_X1 D4752 ( .Y(D4752_Y), .B(D4753_Y), .A(D4783_Y));
KC_NOR2_X1 D4737 ( .Y(D4737_Y), .B(D4696_Y), .A(D4736_Y));
KC_NOR2_X1 D4736 ( .Y(D4736_Y), .B(D3126_Y), .A(D1607_Y));
KC_NOR2_X1 D4694 ( .Y(D4694_Y), .B(D4636_Q), .A(D4637_Q));
KC_NOR2_X1 D4687 ( .Y(D4687_Y), .B(D4591_Y), .A(D369_Y));
KC_NOR2_X1 D4679 ( .Y(D4679_Y), .B(D4704_Y), .A(D4738_Y));
KC_NOR2_X1 D4678 ( .Y(D4678_Y), .B(D4705_Y), .A(D4738_Y));
KC_NOR2_X1 D4670 ( .Y(D4670_Y), .B(D1622_Y), .A(D4672_Y));
KC_NOR2_X1 D4665 ( .Y(D4665_Y), .B(D4672_Y), .A(D1622_Y));
KC_NOR2_X1 D4657 ( .Y(D4657_Y), .B(D3203_Y), .A(D4591_Y));
KC_NOR2_X1 D4656 ( .Y(D4656_Y), .B(D3203_Y), .A(D3298_Y));
KC_NOR2_X1 D4655 ( .Y(D4655_Y), .B(D3097_Y), .A(D4591_Y));
KC_NOR2_X1 D4597 ( .Y(D4597_Y), .B(D4650_Y), .A(D4640_Q));
KC_NOR2_X1 D4595 ( .Y(D4595_Y), .B(D4586_Y), .A(D4637_Q));
KC_NOR2_X1 D4594 ( .Y(D4594_Y), .B(D4586_Y), .A(D4581_Y));
KC_NOR2_X1 D4593 ( .Y(D4593_Y), .B(D166_Y), .A(D4629_Y));
KC_NOR2_X1 D4592 ( .Y(D4592_Y), .B(D4594_Y), .A(D4637_Q));
KC_NOR2_X1 D4590 ( .Y(D4590_Y), .B(D3150_Y), .A(D3131_Y));
KC_NOR2_X1 D4578 ( .Y(D4578_Y), .B(D4579_Y), .A(D4640_Q));
KC_NOR2_X1 D4574 ( .Y(D4574_Y), .B(D4585_Y), .A(D3112_Y));
KC_NOR2_X1 D4508 ( .Y(D4508_Y), .B(D4509_Y), .A(D3026_Y));
KC_NOR2_X1 D4503 ( .Y(D4503_Y), .B(D4509_Y), .A(D3020_Y));
KC_NOR2_X1 D4502 ( .Y(D4502_Y), .B(D3038_Y), .A(D4508_Y));
KC_NOR2_X1 D4501 ( .Y(D4501_Y), .B(D1515_Q), .A(D3080_Q));
KC_NOR2_X1 D4497 ( .Y(D4497_Y), .B(D4528_Y), .A(D4508_Y));
KC_NOR2_X1 D4444 ( .Y(D4444_Y), .B(D4434_Y), .A(D4116_Y));
KC_NOR2_X1 D4438 ( .Y(D4438_Y), .B(D4440_Y), .A(D228_Q));
KC_NOR2_X1 D4431 ( .Y(D4431_Y), .B(D4416_Y), .A(D1713_Y));
KC_NOR2_X1 D4424 ( .Y(D4424_Y), .B(D4422_Y), .A(D239_Q));
KC_NOR2_X1 D4418 ( .Y(D4418_Y), .B(D165_Y), .A(D4294_Y));
KC_NOR2_X1 D4414 ( .Y(D4414_Y), .B(D4743_Q), .A(D4516_Y));
KC_NOR2_X1 D4408 ( .Y(D4408_Y), .B(D8313_Q), .A(D228_Q));
KC_NOR2_X1 D4357 ( .Y(D4357_Y), .B(D4359_Y), .A(D4131_Y));
KC_NOR2_X1 D4356 ( .Y(D4356_Y), .B(D4316_Y), .A(D4349_Y));
KC_NOR2_X1 D4355 ( .Y(D4355_Y), .B(D4384_Y), .A(D4402_Y));
KC_NOR2_X1 D4354 ( .Y(D4354_Y), .B(D4306_Y), .A(D4291_Y));
KC_NOR2_X1 D4346 ( .Y(D4346_Y), .B(D4335_Y), .A(D4402_Y));
KC_NOR2_X1 D4345 ( .Y(D4345_Y), .B(D5651_Y), .A(D4301_Y));
KC_NOR2_X1 D4336 ( .Y(D4336_Y), .B(D5890_Y), .A(D4340_Y));
KC_NOR2_X1 D4335 ( .Y(D4335_Y), .B(D4338_Y), .A(D4349_Y));
KC_NOR2_X1 D4334 ( .Y(D4334_Y), .B(D5928_Y), .A(D4373_Y));
KC_NOR2_X1 D4313 ( .Y(D4313_Y), .B(D1721_Y), .A(D5990_Y));
KC_NOR2_X1 D4312 ( .Y(D4312_Y), .B(D4300_Y), .A(D4381_Y));
KC_NOR2_X1 D4311 ( .Y(D4311_Y), .B(D4282_Y), .A(D4306_Y));
KC_NOR2_X1 D4308 ( .Y(D4308_Y), .B(D4392_Y), .A(D4366_Y));
KC_NOR2_X1 D4301 ( .Y(D4301_Y), .B(D1629_Y), .A(D148_Q));
KC_NOR2_X1 D4300 ( .Y(D4300_Y), .B(D4303_Y), .A(D4301_Y));
KC_NOR2_X1 D4299 ( .Y(D4299_Y), .B(D4350_Y), .A(D4304_Y));
KC_NOR2_X1 D4291 ( .Y(D4291_Y), .B(D4449_Y), .A(D4447_Y));
KC_NOR2_X1 D4290 ( .Y(D4290_Y), .B(D1721_Y), .A(D286_Y));
KC_NOR2_X1 D4289 ( .Y(D4289_Y), .B(D4327_Y), .A(D148_Q));
KC_NOR2_X1 D4288 ( .Y(D4288_Y), .B(D4282_Y), .A(D1629_Y));
KC_NOR2_X1 D4287 ( .Y(D4287_Y), .B(D6070_Y), .A(D5837_Y));
KC_NOR2_X1 D4277 ( .Y(D4277_Y), .B(D4465_Y), .A(D4380_Y));
KC_NOR2_X1 D4276 ( .Y(D4276_Y), .B(D7316_Y), .A(D4414_Y));
KC_NOR2_X1 D4204 ( .Y(D4204_Y), .B(D4118_Q), .A(D4122_Q));
KC_NOR2_X1 D4196 ( .Y(D4196_Y), .B(D5847_Y), .A(D1722_Y));
KC_NOR2_X1 D4186 ( .Y(D4186_Y), .B(D5752_Y), .A(D4178_Y));
KC_NOR2_X1 D4178 ( .Y(D4178_Y), .B(D4374_Y), .A(D5867_Y));
KC_NOR2_X1 D4171 ( .Y(D4171_Y), .B(D4358_Y), .A(D4304_Y));
KC_NOR2_X1 D4099 ( .Y(D4099_Y), .B(D7783_Y), .A(D16135_Y));
KC_NOR2_X1 D4095 ( .Y(D4095_Y), .B(D4102_Y), .A(D4120_Q));
KC_NOR2_X1 D4093 ( .Y(D4093_Y), .B(D4231_Y), .A(D4127_Y));
KC_NOR2_X1 D4092 ( .Y(D4092_Y), .B(D4197_Y), .A(D4121_Q));
KC_NOR2_X1 D3841 ( .Y(D3841_Y), .B(D6260_Y), .A(D497_Y));
KC_NOR2_X1 D3713 ( .Y(D3713_Y), .B(D6792_Y), .A(D5214_Y));
KC_NOR2_X1 D3600 ( .Y(D3600_Y), .B(D1474_Y), .A(D3646_Q));
KC_NOR2_X1 D3535 ( .Y(D3535_Y), .B(D1526_Y), .A(D3554_Y));
KC_NOR2_X1 D3532 ( .Y(D3532_Y), .B(D3550_Y), .A(D4897_Y));
KC_NOR2_X1 D3531 ( .Y(D3531_Y), .B(D3405_Y), .A(D3388_Q));
KC_NOR2_X1 D3527 ( .Y(D3527_Y), .B(D4911_Y), .A(D3526_Y));
KC_NOR2_X1 D3526 ( .Y(D3526_Y), .B(D3525_Y), .A(D3522_Y));
KC_NOR2_X1 D3525 ( .Y(D3525_Y), .B(D1570_Y), .A(D3576_Q));
KC_NOR2_X1 D3501 ( .Y(D3501_Y), .B(D3516_Y), .A(D5020_Y));
KC_NOR2_X1 D3446 ( .Y(D3446_Y), .B(D3448_Y), .A(D3416_Y));
KC_NOR2_X1 D3442 ( .Y(D3442_Y), .B(D3415_Y), .A(D4923_Y));
KC_NOR2_X1 D3437 ( .Y(D3437_Y), .B(D3599_Y), .A(D3498_Y));
KC_NOR2_X1 D3426 ( .Y(D3426_Y), .B(D3371_Y), .A(D3599_Y));
KC_NOR2_X1 D3419 ( .Y(D3419_Y), .B(D3428_Y), .A(D3477_Y));
KC_NOR2_X1 D3413 ( .Y(D3413_Y), .B(D3428_Y), .A(D4915_Y));
KC_NOR2_X1 D3410 ( .Y(D3410_Y), .B(D3405_Y), .A(D4867_Y));
KC_NOR2_X1 D3409 ( .Y(D3409_Y), .B(D4960_Y), .A(D3477_Y));
KC_NOR2_X1 D3408 ( .Y(D3408_Y), .B(D3516_Y), .A(D4882_Y));
KC_NOR2_X1 D3330 ( .Y(D3330_Y), .B(D3320_Y), .A(D3332_Y));
KC_NOR2_X1 D3329 ( .Y(D3329_Y), .B(D3332_Y), .A(D3208_Y));
KC_NOR2_X1 D3324 ( .Y(D3324_Y), .B(D406_Y), .A(D7641_Y));
KC_NOR2_X1 D3323 ( .Y(D3323_Y), .B(D3317_Y), .A(D3275_Y));
KC_NOR2_X1 D3322 ( .Y(D3322_Y), .B(D3318_Y), .A(D3347_Y));
KC_NOR2_X1 D3321 ( .Y(D3321_Y), .B(D1453_Y), .A(D3349_Y));
KC_NOR2_X1 D3314 ( .Y(D3314_Y), .B(D3315_Y), .A(D3377_Y));
KC_NOR2_X1 D3311 ( .Y(D3311_Y), .B(D3338_Y), .A(D3376_Q));
KC_NOR2_X1 D3308 ( .Y(D3308_Y), .B(D3375_Q), .A(D3373_Q));
KC_NOR2_X1 D3238 ( .Y(D3238_Y), .B(D1425_Y), .A(D3283_Q));
KC_NOR2_X1 D3233 ( .Y(D3233_Y), .B(D1423_Y), .A(D3282_Q));
KC_NOR2_X1 D3232 ( .Y(D3232_Y), .B(D3281_Q), .A(D3282_Q));
KC_NOR2_X1 D3231 ( .Y(D3231_Y), .B(D3137_Y), .A(D3234_Y));
KC_NOR2_X1 D3205 ( .Y(D3205_Y), .B(D3215_Y), .A(D3368_Y));
KC_NOR2_X1 D3204 ( .Y(D3204_Y), .B(D3052_Y), .A(D3383_Q));
KC_NOR2_X1 D3203 ( .Y(D3203_Y), .B(D3320_Y), .A(D3206_Y));
KC_NOR2_X1 D3150 ( .Y(D3150_Y), .B(D3152_Y), .A(D1457_Y));
KC_NOR2_X1 D3149 ( .Y(D3149_Y), .B(D3146_Y), .A(D3186_Q));
KC_NOR2_X1 D3140 ( .Y(D3140_Y), .B(D1458_Y), .A(D3188_Q));
KC_NOR2_X1 D3139 ( .Y(D3139_Y), .B(D3188_Q), .A(D3144_Y));
KC_NOR2_X1 D3138 ( .Y(D3138_Y), .B(D3145_Y), .A(D3186_Q));
KC_NOR2_X1 D3131 ( .Y(D3131_Y), .B(D3132_Y), .A(D3148_Y));
KC_NOR2_X1 D3130 ( .Y(D3130_Y), .B(D3186_Q), .A(D3189_Q));
KC_NOR2_X1 D3129 ( .Y(D3129_Y), .B(D3134_Y), .A(D3189_Q));
KC_NOR2_X1 D3128 ( .Y(D3128_Y), .B(D3192_Y), .A(D3132_Y));
KC_NOR2_X1 D3127 ( .Y(D3127_Y), .B(D3192_Y), .A(D3133_Y));
KC_NOR2_X1 D3126 ( .Y(D3126_Y), .B(D3135_Y), .A(D3131_Y));
KC_NOR2_X1 D3125 ( .Y(D3125_Y), .B(D3148_Y), .A(D3133_Y));
KC_NOR2_X1 D3123 ( .Y(D3123_Y), .B(D3182_Y), .A(D3170_Y));
KC_NOR2_X1 D3122 ( .Y(D3122_Y), .B(D3182_Y), .A(D3170_Y));
KC_NOR2_X1 D3117 ( .Y(D3117_Y), .B(D3119_Y), .A(D3150_Y));
KC_NOR2_X1 D3112 ( .Y(D3112_Y), .B(D3165_Y), .A(D3172_Y));
KC_NOR2_X1 D3106 ( .Y(D3106_Y), .B(D3159_Y), .A(D3127_Y));
KC_NOR2_X1 D3101 ( .Y(D3101_Y), .B(D3100_Y), .A(D7641_Y));
KC_NOR2_X1 D3098 ( .Y(D3098_Y), .B(D1429_Y), .A(D3234_Y));
KC_NOR2_X1 D3097 ( .Y(D3097_Y), .B(D3234_Y), .A(D3116_Y));
KC_NOR2_X1 D3025 ( .Y(D3025_Y), .B(D3079_Q), .A(D3078_Q));
KC_NOR2_X1 D3024 ( .Y(D3024_Y), .B(D3043_Y), .A(D1516_Q));
KC_NOR2_X1 D2904 ( .Y(D2904_Y), .B(D2996_Y), .A(D2954_Y));
KC_NOR2_X1 D2843 ( .Y(D2843_Y), .B(D2839_Y), .A(D2847_Y));
KC_NOR2_X1 D2842 ( .Y(D2842_Y), .B(D2843_Y), .A(D2888_Q));
KC_NOR2_X1 D2837 ( .Y(D2837_Y), .B(D2804_Y), .A(D2887_Q));
KC_NOR2_X1 D2836 ( .Y(D2836_Y), .B(D2890_Q), .A(D2888_Q));
KC_NOR2_X1 D2834 ( .Y(D2834_Y), .B(D2775_Y), .A(D2750_Y));
KC_NOR2_X1 D2833 ( .Y(D2833_Y), .B(D2817_Y), .A(D2832_Y));
KC_NOR2_X1 D2828 ( .Y(D2828_Y), .B(D2876_Y), .A(D2804_Y));
KC_NOR2_X1 D2827 ( .Y(D2827_Y), .B(D2778_Y), .A(D2750_Y));
KC_NOR2_X1 D2823 ( .Y(D2823_Y), .B(D2885_Q), .A(D2884_Q));
KC_NOR2_X1 D2822 ( .Y(D2822_Y), .B(D2825_Y), .A(D2826_Y));
KC_NOR2_X1 D2819 ( .Y(D2819_Y), .B(D2765_Y), .A(D2836_Y));
KC_NOR2_X1 D2813 ( .Y(D2813_Y), .B(D2760_Y), .A(D2812_Y));
KC_NOR2_X1 D2812 ( .Y(D2812_Y), .B(D2845_Y), .A(D2778_Y));
KC_NOR2_X1 D2762 ( .Y(D2762_Y), .B(D2752_Y), .A(D2764_Y));
KC_NOR2_X1 D2761 ( .Y(D2761_Y), .B(D2745_Y), .A(D2795_Q));
KC_NOR2_X1 D2760 ( .Y(D2760_Y), .B(D2745_Y), .A(D2799_Q));
KC_NOR2_X1 D2756 ( .Y(D2756_Y), .B(D2886_Q), .A(D2801_Q));
KC_NOR2_X1 D2755 ( .Y(D2755_Y), .B(D2757_Y), .A(D1441_Y));
KC_NOR2_X1 D2752 ( .Y(D2752_Y), .B(D2755_Y), .A(D2816_Q));
KC_NOR2_X1 D2749 ( .Y(D2749_Y), .B(D2858_Y), .A(D2766_Y));
KC_NOR2_X1 D2660 ( .Y(D2660_Y), .B(D2658_Y), .A(D16597_Y));
KC_NOR2_X1 D2659 ( .Y(D2659_Y), .B(D16277_Y), .A(D16275_Y));
KC_NOR2_X1 D2658 ( .Y(D2658_Y), .B(D15475_Y), .A(D16192_Y));
KC_NOR2_X1 D2657 ( .Y(D2657_Y), .B(D16264_Y), .A(D16277_Y));
KC_NOR2_X1 D2656 ( .Y(D2656_Y), .B(D16257_Y), .A(D13392_Y));
KC_NOR2_X1 D2618 ( .Y(D2618_Y), .B(D15289_Y), .A(D15306_Y));
KC_NOR2_X1 D2615 ( .Y(D2615_Y), .B(D16275_Y), .A(D16271_Y));
KC_NOR2_X1 D2614 ( .Y(D2614_Y), .B(D15479_Y), .A(D15484_Y));
KC_NOR2_X1 D2605 ( .Y(D2605_Y), .B(D15483_Y), .A(D15484_Y));
KC_NOR2_X1 D2604 ( .Y(D2604_Y), .B(D14728_Y), .A(D15562_Y));
KC_NOR2_X1 D2589 ( .Y(D2589_Y), .B(D15394_Y), .A(D16068_Y));
KC_NOR2_X1 D2588 ( .Y(D2588_Y), .B(D2591_Y), .A(D15279_Y));
KC_NOR2_X1 D2587 ( .Y(D2587_Y), .B(D15394_Y), .A(D2654_Y));
KC_NOR2_X1 D2545 ( .Y(D2545_Y), .B(D2546_Y), .A(D2512_Y));
KC_NOR2_X1 D2544 ( .Y(D2544_Y), .B(D2563_Y), .A(D14567_Y));
KC_NOR2_X1 D2536 ( .Y(D2536_Y), .B(D952_Q), .A(D2538_Y));
KC_NOR2_X1 D2528 ( .Y(D2528_Y), .B(D15887_Y), .A(D15031_Y));
KC_NOR2_X1 D2496 ( .Y(D2496_Y), .B(D14018_Y), .A(D14132_Y));
KC_NOR2_X1 D2492 ( .Y(D2492_Y), .B(D14133_Y), .A(D13379_Y));
KC_NOR2_X1 D2491 ( .Y(D2491_Y), .B(D14134_Y), .A(D13379_Y));
KC_NOR2_X1 D2434 ( .Y(D2434_Y), .B(D13305_Y), .A(D13298_Y));
KC_NOR2_X1 D2433 ( .Y(D2433_Y), .B(D13321_Y), .A(D13308_Y));
KC_NOR2_X1 D2432 ( .Y(D2432_Y), .B(D13410_Y), .A(D13314_Y));
KC_NOR2_X1 D2431 ( .Y(D2431_Y), .B(D12732_Y), .A(D2343_Y));
KC_NOR2_X1 D2430 ( .Y(D2430_Y), .B(D13308_Y), .A(D13309_Y));
KC_NOR2_X1 D2429 ( .Y(D2429_Y), .B(D13322_Y), .A(D13308_Y));
KC_NOR2_X1 D2418 ( .Y(D2418_Y), .B(D14200_Y), .A(D13536_Y));
KC_NOR2_X1 D2417 ( .Y(D2417_Y), .B(D13536_Y), .A(D12889_Y));
KC_NOR2_X1 D2416 ( .Y(D2416_Y), .B(D13665_Y), .A(D13536_Y));
KC_NOR2_X1 D2405 ( .Y(D2405_Y), .B(D12720_Y), .A(D7670_Y));
KC_NOR2_X1 D2378 ( .Y(D2378_Y), .B(D12842_Y), .A(D13392_Y));
KC_NOR2_X1 D2363 ( .Y(D2363_Y), .B(D2343_Y), .A(D2312_Y));
KC_NOR2_X1 D2360 ( .Y(D2360_Y), .B(D12664_Y), .A(D2379_Y));
KC_NOR2_X1 D2326 ( .Y(D2326_Y), .B(D12316_Y), .A(D12780_Y));
KC_NOR2_X1 D2325 ( .Y(D2325_Y), .B(D12316_Y), .A(D12783_Y));
KC_NOR2_X1 D2310 ( .Y(D2310_Y), .B(D11657_Y), .A(D10179_Y));
KC_NOR2_X1 D2309 ( .Y(D2309_Y), .B(D12196_Y), .A(D7668_Y));
KC_NOR2_X1 D2308 ( .Y(D2308_Y), .B(D12196_Y), .A(D6287_Y));
KC_NOR2_X1 D2307 ( .Y(D2307_Y), .B(D12196_Y), .A(D7670_Y));
KC_NOR2_X1 D2273 ( .Y(D2273_Y), .B(D11960_Y), .A(D11955_Y));
KC_NOR2_X1 D2272 ( .Y(D2272_Y), .B(D1108_Y), .A(D11941_Y));
KC_NOR2_X1 D2271 ( .Y(D2271_Y), .B(D11961_Y), .A(D11945_Y));
KC_NOR2_X1 D2190 ( .Y(D2190_Y), .B(D10988_Y), .A(D10936_Y));
KC_NOR2_X1 D2189 ( .Y(D2189_Y), .B(D10988_Y), .A(D10972_Y));
KC_NOR2_X1 D2184 ( .Y(D2184_Y), .B(D10989_Y), .A(D10972_Y));
KC_NOR2_X1 D2183 ( .Y(D2183_Y), .B(D10989_Y), .A(D10936_Y));
KC_NOR2_X1 D2137 ( .Y(D2137_Y), .B(D10045_Y), .A(D2162_Y));
KC_NOR2_X1 D2026 ( .Y(D2026_Y), .B(D8748_Y), .A(D9482_Y));
KC_NOR2_X1 D2025 ( .Y(D2025_Y), .B(D8918_Y), .A(D305_Q));
KC_NOR2_X1 D2015 ( .Y(D2015_Y), .B(D9072_Y), .A(D7361_Y));
KC_NOR2_X1 D2007 ( .Y(D2007_Y), .B(D9115_Y), .A(D2008_Y));
KC_NOR2_X1 D1984 ( .Y(D1984_Y), .B(D1988_Y), .A(D9471_Q));
KC_NOR2_X1 D1983 ( .Y(D1983_Y), .B(D9550_Y), .A(D9432_Y));
KC_NOR2_X1 D1981 ( .Y(D1981_Y), .B(D9645_Y), .A(D8365_Y));
KC_NOR2_X1 D1980 ( .Y(D1980_Y), .B(D9681_Y), .A(D8365_Y));
KC_NOR2_X1 D1979 ( .Y(D1979_Y), .B(D9726_Y), .A(D8365_Y));
KC_NOR2_X1 D1886 ( .Y(D1886_Y), .B(D355_Y), .A(D7227_Y));
KC_NOR2_X1 D1883 ( .Y(D1883_Y), .B(D7359_Y), .A(D7295_Y));
KC_NOR2_X1 D1878 ( .Y(D1878_Y), .B(D1753_Y), .A(D1906_Y));
KC_NOR2_X1 D1877 ( .Y(D1877_Y), .B(D1880_Y), .A(D7334_Y));
KC_NOR2_X1 D1870 ( .Y(D1870_Y), .B(D6083_Y), .A(D6001_Y));
KC_NOR2_X1 D1869 ( .Y(D1869_Y), .B(D6083_Y), .A(D1709_Y));
KC_NOR2_X1 D1868 ( .Y(D1868_Y), .B(D1963_Y), .A(D6083_Y));
KC_NOR2_X1 D1864 ( .Y(D1864_Y), .B(D1904_Y), .A(D2008_Y));
KC_NOR2_X1 D1863 ( .Y(D1863_Y), .B(D9268_Y), .A(D346_Y));
KC_NOR2_X1 D1854 ( .Y(D1854_Y), .B(D1850_Y), .A(D7932_Y));
KC_NOR2_X1 D1853 ( .Y(D1853_Y), .B(D7923_Y), .A(D531_Q));
KC_NOR2_X1 D1852 ( .Y(D1852_Y), .B(D7955_Y), .A(D7923_Y));
KC_NOR2_X1 D1847 ( .Y(D1847_Y), .B(D8017_Y), .A(D7668_Y));
KC_NOR2_X1 D1843 ( .Y(D1843_Y), .B(D8102_Y), .A(D8007_Y));
KC_NOR2_X1 D1827 ( .Y(D1827_Y), .B(D1935_Y), .A(D105_Y));
KC_NOR2_X1 D1740 ( .Y(D1740_Y), .B(D5852_Y), .A(D247_Y));
KC_NOR2_X1 D1728 ( .Y(D1728_Y), .B(D5886_Y), .A(D1739_Y));
KC_NOR2_X1 D1727 ( .Y(D1727_Y), .B(D7211_Y), .A(D7334_Y));
KC_NOR2_X1 D1726 ( .Y(D1726_Y), .B(D1728_Y), .A(D7469_Y));
KC_NOR2_X1 D1719 ( .Y(D1719_Y), .B(D5857_Y), .A(D6113_Y));
KC_NOR2_X1 D1709 ( .Y(D1709_Y), .B(D5960_Y), .A(D5872_Y));
KC_NOR2_X1 D1708 ( .Y(D1708_Y), .B(D7629_Y), .A(D4416_Y));
KC_NOR2_X1 D1704 ( .Y(D1704_Y), .B(D7785_Y), .A(D7563_Y));
KC_NOR2_X1 D1697 ( .Y(D1697_Y), .B(D6433_Y), .A(D485_Q));
KC_NOR2_X1 D1696 ( .Y(D1696_Y), .B(D6465_Y), .A(D1745_Y));
KC_NOR2_X1 D1695 ( .Y(D1695_Y), .B(D4961_Y), .A(D6465_Y));
KC_NOR2_X1 D1690 ( .Y(D1690_Y), .B(D6783_Y), .A(D1932_Y));
KC_NOR2_X1 D1689 ( .Y(D1689_Y), .B(D6795_Y), .A(D6782_Y));
KC_NOR2_X1 D1688 ( .Y(D1688_Y), .B(D875_Y), .A(D6782_Y));
KC_NOR2_X1 D1682 ( .Y(D1682_Y), .B(D6943_Y), .A(D6935_Y));
KC_NOR2_X1 D1590 ( .Y(D1590_Y), .B(D4359_Y), .A(D6034_Y));
KC_NOR2_X1 D1581 ( .Y(D1581_Y), .B(D1584_Y), .A(D4444_Y));
KC_NOR2_X1 D1572 ( .Y(D1572_Y), .B(D1574_Y), .A(D4637_Q));
KC_NOR2_X1 D1568 ( .Y(D1568_Y), .B(D4922_Y), .A(D4941_Y));
KC_NOR2_X1 D1567 ( .Y(D1567_Y), .B(D1570_Y), .A(D4911_Y));
KC_NOR2_X1 D1563 ( .Y(D1563_Y), .B(D4869_Y), .A(D4960_Y));
KC_NOR2_X1 D1562 ( .Y(D1562_Y), .B(D4914_Y), .A(D4910_Y));
KC_NOR2_X1 D1555 ( .Y(D1555_Y), .B(D5372_Y), .A(D5259_Y));
KC_NOR2_X1 D1554 ( .Y(D1554_Y), .B(D875_Y), .A(D5259_Y));
KC_NOR2_X1 D54 ( .Y(D54_Y), .B(D7641_Y), .A(D53_Y));
KC_NOR2_X1 D53 ( .Y(D53_Y), .B(D4596_Y), .A(D307_Y));
KC_NOR2_X1 D1438 ( .Y(D1438_Y), .B(D2738_Y), .A(D2820_Y));
KC_NOR2_X1 D1437 ( .Y(D1437_Y), .B(D1434_Y), .A(D2818_Y));
KC_NOR2_X1 D1436 ( .Y(D1436_Y), .B(D2738_Y), .A(D2836_Y));
KC_NOR2_X1 D1435 ( .Y(D1435_Y), .B(D2765_Y), .A(D2820_Y));
KC_NOR2_X1 D1430 ( .Y(D1430_Y), .B(D3190_Q), .A(D3187_Q));
KC_NOR2_X1 D1422 ( .Y(D1422_Y), .B(D3237_Y), .A(D3283_Q));
KC_NOR2_X1 D1421 ( .Y(D1421_Y), .B(D1468_Y), .A(D1424_Y));
KC_NOR2_X1 D1419 ( .Y(D1419_Y), .B(D1417_Y), .A(D1519_Y));
KC_NOR2_X1 D1415 ( .Y(D1415_Y), .B(D3521_Y), .A(D5044_Y));
KC_NOR2_X1 D1407 ( .Y(D1407_Y), .B(D6260_Y), .A(D497_Y));
KC_NOR2_X1 D1343 ( .Y(D1343_Y), .B(D1341_Y), .A(D16542_Y));
KC_NOR2_X1 D1281 ( .Y(D1281_Y), .B(D1271_Y), .A(D1378_Q));
KC_NOR2_X1 D1274 ( .Y(D1274_Y), .B(D13775_Y), .A(D13810_Q));
KC_NOR2_X1 D1272 ( .Y(D1272_Y), .B(D15963_Y), .A(D15937_S));
KC_NOR2_X1 D1091 ( .Y(D1091_Y), .B(D13536_Y), .A(D12949_Y));
KC_NOR2_X1 D1084 ( .Y(D1084_Y), .B(D9742_Y), .A(D8422_Y));
KC_NOR2_X1 D1082 ( .Y(D1082_Y), .B(D1597_Y), .A(D5520_Y));
KC_NOR2_X1 D984 ( .Y(D984_Y), .B(D874_Y), .A(D14137_Y));
KC_NOR2_X1 D979 ( .Y(D979_Y), .B(D1107_Y), .A(D10905_Y));
KC_NOR2_X1 D973 ( .Y(D973_Y), .B(D5451_Y), .A(D5441_Y));
KC_NOR2_X1 D972 ( .Y(D972_Y), .B(D5452_Y), .A(D5442_Y));
KC_NOR2_X1 D962 ( .Y(D962_Y), .B(D13330_Y), .A(D14132_Y));
KC_NOR2_X1 D865 ( .Y(D865_Y), .B(D10856_Y), .A(D10321_Y));
KC_NOR2_X1 D854 ( .Y(D854_Y), .B(D8264_Y), .A(D1944_Q));
KC_NOR2_X1 D756 ( .Y(D756_Y), .B(D845_Y), .A(D845_Y));
KC_NOR2_X1 D755 ( .Y(D755_Y), .B(D14564_Y), .A(D15611_Y));
KC_NOR2_X1 D753 ( .Y(D753_Y), .B(D841_Y), .A(D13392_Y));
KC_NOR2_X1 D640 ( .Y(D640_Y), .B(D14653_Y), .A(D14046_Y));
KC_NOR2_X1 D625 ( .Y(D625_Y), .B(D739_Y), .A(D8242_Y));
KC_NOR2_X1 D572 ( .Y(D572_Y), .B(D15302_Y), .A(D15310_Y));
KC_NOR2_X1 D567 ( .Y(D567_Y), .B(D16090_Y), .A(D16088_Y));
KC_NOR2_X1 D566 ( .Y(D566_Y), .B(D15302_Y), .A(D15278_Y));
KC_NOR2_X1 D373 ( .Y(D373_Y), .B(D481_Y), .A(D7563_Y));
KC_NOR2_X1 D344 ( .Y(D344_Y), .B(D4631_Y), .A(D3142_Y));
KC_NOR2_X1 D343 ( .Y(D343_Y), .B(D102_Y), .A(D6177_Y));
KC_NOR2_X1 D288 ( .Y(D288_Y), .B(D6045_Y), .A(D7094_Y));
KC_NOR2_X1 D286 ( .Y(D286_Y), .B(D280_Y), .A(D5970_Y));
KC_NOR2_X1 D283 ( .Y(D283_Y), .B(D2127_Y), .A(D326_Q));
KC_NOR2_X1 D280 ( .Y(D280_Y), .B(D5974_Y), .A(D4415_Y));
KC_NOR2_X1 D277 ( .Y(D277_Y), .B(D5956_Y), .A(D8313_Q));
KC_NOR2_X1 D275 ( .Y(D275_Y), .B(D4149_Q), .A(D8313_Q));
KC_NOR2_X1 D249 ( .Y(D249_Y), .B(D5999_Y), .A(D4298_Y));
KC_NOR2_X1 D245 ( .Y(D245_Y), .B(D8866_Y), .A(D8896_Q));
KC_NOR2_X1 D205 ( .Y(D205_Y), .B(D5725_Y), .A(D208_Y));
KC_NOR2_X1 D201 ( .Y(D201_Y), .B(D5724_Y), .A(D5703_Y));
KC_NOR2_X1 D177 ( .Y(D177_Y), .B(D5673_Y), .A(D5668_Y));
KC_NOR2_X1 D174 ( .Y(D174_Y), .B(D7120_Y), .A(D7107_Y));
KC_NOR2_X1 D173 ( .Y(D173_Y), .B(D9922_Y), .A(D223_Y));
KC_NOR2_X1 D84 ( .Y(D84_Y), .B(D2591_Y), .A(D15271_Y));
KC_NOR2_X1 D77 ( .Y(D77_Y), .B(D12196_Y), .A(D7669_Y));
KC_NOR2_X1 D70 ( .Y(D70_Y), .B(D382_Y), .A(D9269_Y));
KC_NOR2_X1 D68 ( .Y(D68_Y), .B(D5036_Y), .A(D3426_Y));
KC_NOR2_X1 D65 ( .Y(D65_Y), .B(D8424_Y), .A(D8365_Y));
KC_NOR2_X1 D64 ( .Y(D64_Y), .B(D8497_Y), .A(D8422_Y));
KC_AOI22_X1 D16245 ( .A1(D15475_Y), .B0(D16289_Q), .B1(D15630_Y),     .Y(D16245_Y), .A0(D16270_Y));
KC_AOI22_X1 D16050 ( .A1(D16094_Y), .B0(D16059_Y), .B1(D16051_Y),     .Y(D16050_Y), .A0(D15335_Y));
KC_AOI22_X1 D15970 ( .A1(D13636_Y), .B0(D15998_Q), .B1(D1073_Y),     .Y(D15970_Y), .A0(D16010_Q));
KC_AOI22_X1 D15967 ( .A1(D13640_Y), .B0(D16013_Q), .B1(D2476_Y),     .Y(D15967_Y), .A0(D15994_Q));
KC_AOI22_X1 D15965 ( .A1(D13524_Y), .B0(D15999_Q), .B1(D14224_Y),     .Y(D15965_Y), .A0(D15992_Q));
KC_AOI22_X1 D15959 ( .A1(D13636_Y), .B0(D16012_Q), .B1(D1073_Y),     .Y(D15959_Y), .A0(D15991_Q));
KC_AOI22_X1 D15915 ( .A1(D14253_Y), .B0(D15999_Q), .B1(D936_Y),     .Y(D15915_Y), .A0(D1326_Q));
KC_AOI22_X1 D15914 ( .A1(D13629_Y), .B0(D1229_Q), .B1(D2476_Y),     .Y(D15914_Y), .A0(D15949_Q));
KC_AOI22_X1 D15911 ( .A1(D14253_Y), .B0(D15949_Q), .B1(D14254_Y),     .Y(D15911_Y), .A0(D16388_Q));
KC_AOI22_X1 D15907 ( .A1(D13640_Y), .B0(D16392_Q), .B1(D2476_Y),     .Y(D15907_Y), .A0(D1234_Q));
KC_AOI22_X1 D15906 ( .A1(D13525_Y), .B0(D16391_Q), .B1(D2475_Y),     .Y(D15906_Y), .A0(D2638_Q));
KC_AOI22_X1 D15905 ( .A1(D13525_Y), .B0(D15995_Q), .B1(D2475_Y),     .Y(D15905_Y), .A0(D15948_Q));
KC_AOI22_X1 D15903 ( .A1(D13525_Y), .B0(D15997_Q), .B1(D2475_Y),     .Y(D15903_Y), .A0(D1230_Q));
KC_AOI22_X1 D15902 ( .A1(D13524_Y), .B0(D16389_Q), .B1(D14224_Y),     .Y(D15902_Y), .A0(D1233_Q));
KC_AOI22_X1 D15890 ( .A1(D13634_Y), .B0(D1236_Q), .B1(D1071_Y),     .Y(D15890_Y), .A0(D16388_Q));
KC_AOI22_X1 D15886 ( .A1(D14175_Y), .B0(D15992_Q), .B1(D14174_Y),     .Y(D15886_Y), .A0(D15991_Q));
KC_AOI22_X1 D15885 ( .A1(D14175_Y), .B0(D15947_Q), .B1(D14174_Y),     .Y(D15885_Y), .A0(D16010_Q));
KC_AOI22_X1 D15880 ( .A1(D14172_Y), .B0(D1229_Q), .B1(D14252_Y),     .Y(D15880_Y), .A0(D15998_Q));
KC_AOI22_X1 D15879 ( .A1(D14257_Y), .B0(D1228_Q), .B1(D936_Y),     .Y(D15879_Y), .A0(D1236_Q));
KC_AOI22_X1 D15878 ( .A1(D13524_Y), .B0(D1228_Q), .B1(D14224_Y),     .Y(D15878_Y), .A0(D15947_Q));
KC_AOI22_X1 D15834 ( .A1(D14175_Y), .B0(D1233_Q), .B1(D14174_Y),     .Y(D15834_Y), .A0(D15869_Q));
KC_AOI22_X1 D15833 ( .A1(D14253_Y), .B0(D1234_Q), .B1(D14254_Y),     .Y(D15833_Y), .A0(D142_Q));
KC_AOI22_X1 D15832 ( .A1(D14172_Y), .B0(D16355_Q), .B1(D14252_Y),     .Y(D15832_Y), .A0(D15872_Q));
KC_AOI22_X1 D15830 ( .A1(D13634_Y), .B0(D16358_Q), .B1(D1071_Y),     .Y(D15830_Y), .A0(D16357_Q));
KC_AOI22_X1 D15828 ( .A1(D13636_Y), .B0(D15872_Q), .B1(D1073_Y),     .Y(D15828_Y), .A0(D15870_Q));
KC_AOI22_X1 D15827 ( .A1(D1071_Y), .B0(D1156_Q), .B1(D13634_Y),     .Y(D15827_Y), .A0(D16353_Q));
KC_AOI22_X1 D15825 ( .A1(D14253_Y), .B0(D16363_Q), .B1(D14254_Y),     .Y(D15825_Y), .A0(D1156_Q));
KC_AOI22_X1 D15824 ( .A1(D14224_Y), .B0(D144_Q), .B1(D13524_Y),     .Y(D15824_Y), .A0(D16359_Q));
KC_AOI22_X1 D15817 ( .A1(D14175_Y), .B0(D1148_Q), .B1(D14174_Y),     .Y(D15817_Y), .A0(D15870_Q));
KC_AOI22_X1 D15816 ( .A1(D14257_Y), .B0(D16369_Q), .B1(D936_Y),     .Y(D15816_Y), .A0(D16358_Q));
KC_AOI22_X1 D15815 ( .A1(D14253_Y), .B0(D1149_Q), .B1(D14254_Y),     .Y(D15815_Y), .A0(D16357_Q));
KC_AOI22_X1 D15814 ( .A1(D13525_Y), .B0(D16354_Q), .B1(D2475_Y),     .Y(D15814_Y), .A0(D15868_Q));
KC_AOI22_X1 D15812 ( .A1(D13524_Y), .B0(D16369_Q), .B1(D14224_Y),     .Y(D15812_Y), .A0(D1148_Q));
KC_AOI22_X1 D15811 ( .A1(D13636_Y), .B0(D16364_Q), .B1(D1073_Y),     .Y(D15811_Y), .A0(D15869_Q));
KC_AOI22_X1 D15809 ( .A1(D14172_Y), .B0(D16392_Q), .B1(D14252_Y),     .Y(D15809_Y), .A0(D16364_Q));
KC_AOI22_X1 D15808 ( .A1(D13629_Y), .B0(D16355_Q), .B1(D2476_Y),     .Y(D15808_Y), .A0(D1149_Q));
KC_AOI22_X1 D15744 ( .A1(D13525_Y), .B0(D1074_Q), .B1(D2475_Y),     .Y(D15744_Y), .A0(D15668_Q));
KC_AOI22_X1 D15743 ( .A1(D13524_Y), .B0(D925_Q), .B1(D14224_Y),     .Y(D15743_Y), .A0(D2639_Q));
KC_AOI22_X1 D15742 ( .A1(D14257_Y), .B0(D925_Q), .B1(D936_Y),     .Y(D15742_Y), .A0(D16340_Q));
KC_AOI22_X1 D15741 ( .A1(D13524_Y), .B0(D15797_Q), .B1(D14224_Y),     .Y(D15741_Y), .A0(D2640_Q));
KC_AOI22_X1 D15738 ( .A1(D13629_Y), .B0(D16319_Q), .B1(D2476_Y),     .Y(D15738_Y), .A0(D1053_Q));
KC_AOI22_X1 D15737 ( .A1(D14172_Y), .B0(D16319_Q), .B1(D14252_Y),     .Y(D15737_Y), .A0(D15711_Q));
KC_AOI22_X1 D15736 ( .A1(D14257_Y), .B0(D15797_Q), .B1(D936_Y),     .Y(D15736_Y), .A0(D1077_Q));
KC_AOI22_X1 D15733 ( .A1(D14175_Y), .B0(D2640_Q), .B1(D14174_Y),     .Y(D15733_Y), .A0(D924_Q));
KC_AOI22_X1 D15732 ( .A1(D14253_Y), .B0(D1053_Q), .B1(D14254_Y),     .Y(D15732_Y), .A0(D15796_Q));
KC_AOI22_X1 D15730 ( .A1(D13634_Y), .B0(D16340_Q), .B1(D1071_Y),     .Y(D15730_Y), .A0(D1070_Q));
KC_AOI22_X1 D15727 ( .A1(D13634_Y), .B0(D1077_Q), .B1(D1071_Y),     .Y(D15727_Y), .A0(D15796_Q));
KC_AOI22_X1 D15726 ( .A1(D14253_Y), .B0(D15795_Q), .B1(D14254_Y),     .Y(D15726_Y), .A0(D1070_Q));
KC_AOI22_X1 D15725 ( .A1(D14175_Y), .B0(D15792_Q), .B1(D14174_Y),     .Y(D15725_Y), .A0(D15793_Q));
KC_AOI22_X1 D15724 ( .A1(D13640_Y), .B0(D145_Q), .B1(D2476_Y),     .Y(D15724_Y), .A0(D15795_Q));
KC_AOI22_X1 D15723 ( .A1(D2475_Y), .B0(D15791_Q), .B1(D13525_Y),     .Y(D15723_Y), .A0(D16318_Q));
KC_AOI22_X1 D15721 ( .A1(D2476_Y), .B0(D1050_Q), .B1(D13629_Y),     .Y(D15721_Y), .A0(D16315_Q));
KC_AOI22_X1 D15719 ( .A1(D14172_Y), .B0(D16315_Q), .B1(D14252_Y),     .Y(D15719_Y), .A0(D16317_Q));
KC_AOI22_X1 D15718 ( .A1(D14257_Y), .B0(D16316_Q), .B1(D936_Y),     .Y(D15718_Y), .A0(D16362_Q));
KC_AOI22_X1 D15717 ( .A1(D14253_Y), .B0(D1050_Q), .B1(D14254_Y),     .Y(D15717_Y), .A0(D16346_Q));
KC_AOI22_X1 D15716 ( .A1(D14224_Y), .B0(D15792_Q), .B1(D13524_Y),     .Y(D15716_Y), .A0(D16316_Q));
KC_AOI22_X1 D15713 ( .A1(D1071_Y), .B0(D16346_Q), .B1(D13634_Y),     .Y(D15713_Y), .A0(D16362_Q));
KC_AOI22_X1 D15712 ( .A1(D14257_Y), .B0(D16359_Q), .B1(D936_Y),     .Y(D15712_Y), .A0(D16353_Q));
KC_AOI22_X1 D15708 ( .A1(D15479_Y), .B0(D2609_Y), .B1(D15706_Y),     .Y(D15708_Y), .A0(D15707_Y));
KC_AOI22_X1 D15702 ( .A1(D2609_Y), .B0(D15479_Y), .B1(D15703_Y),     .Y(D15702_Y), .A0(D15704_Y));
KC_AOI22_X1 D15646 ( .A1(D14841_Y), .B0(D2604_Y), .B1(D15627_Y),     .Y(D15646_Y), .A0(D15485_Y));
KC_AOI22_X1 D15645 ( .A1(D15479_Y), .B0(D2604_Y), .B1(D2610_Y),     .Y(D15645_Y), .A0(D15658_Y));
KC_AOI22_X1 D15644 ( .A1(D15480_Y), .B0(D15472_Y), .B1(D15657_Y),     .Y(D15644_Y), .A0(D14846_Y));
KC_AOI22_X1 D15643 ( .A1(D15626_Y), .B0(D2608_Y), .B1(D15647_Y),     .Y(D15643_Y), .A0(D15628_Y));
KC_AOI22_X1 D15642 ( .A1(D15615_Y), .B0(D15480_Y), .B1(D15492_Y),     .Y(D15642_Y), .A0(D15472_Y));
KC_AOI22_X1 D15641 ( .A1(D15488_Y), .B0(D15479_Y), .B1(D15626_Y),     .Y(D15641_Y), .A0(D2609_Y));
KC_AOI22_X1 D15640 ( .A1(D14847_Y), .B0(D15480_Y), .B1(D14867_Y),     .Y(D15640_Y), .A0(D15628_Y));
KC_AOI22_X1 D15639 ( .A1(D14853_Y), .B0(D2608_Y), .B1(D15637_Y),     .Y(D15639_Y), .A0(D15480_Y));
KC_AOI22_X1 D15633 ( .A1(D2583_Y), .B0(D14813_Y), .B1(D16166_Y),     .Y(D15633_Y), .A0(D15562_Y));
KC_AOI22_X1 D15632 ( .A1(D14386_Y), .B0(D14813_Y), .B1(D8888_Y),     .Y(D15632_Y), .A0(D15562_Y));
KC_AOI22_X1 D15631 ( .A1(D15627_Y), .B0(D14847_Y), .B1(D2606_Y),     .Y(D15631_Y), .A0(D15628_Y));
KC_AOI22_X1 D15624 ( .A1(D15656_Y), .B0(D15634_Y), .B1(D15655_Y),     .Y(D15624_Y), .A0(D14829_Y));
KC_AOI22_X1 D15623 ( .A1(D15651_Y), .B0(D8998_Y), .B1(D14840_Y),     .Y(D15623_Y), .A0(D14829_Y));
KC_AOI22_X1 D15622 ( .A1(D15082_Y), .B0(D14813_Y), .B1(D651_Y),     .Y(D15622_Y), .A0(D16461_Y));
KC_AOI22_X1 D15621 ( .A1(D2521_Y), .B0(D14813_Y), .B1(D2870_Y),     .Y(D15621_Y), .A0(D16461_Y));
KC_AOI22_X1 D15620 ( .A1(D14387_Y), .B0(D14813_Y), .B1(D9087_Y),     .Y(D15620_Y), .A0(D16461_Y));
KC_AOI22_X1 D15615 ( .A1(D14311_Y), .B0(D14813_Y), .B1(D9085_Y),     .Y(D15615_Y), .A0(D16461_Y));
KC_AOI22_X1 D15614 ( .A1(D15650_Y), .B0(D15634_Y), .B1(D15661_Y),     .Y(D15614_Y), .A0(D14829_Y));
KC_AOI22_X1 D15613 ( .A1(D15661_Y), .B0(D15634_Y), .B1(D15656_Y),     .Y(D15613_Y), .A0(D14829_Y));
KC_AOI22_X1 D15612 ( .A1(D15655_Y), .B0(D15634_Y), .B1(D15660_Y),     .Y(D15612_Y), .A0(D14829_Y));
KC_AOI22_X1 D15604 ( .A1(D15345_Y), .B0(D15348_Y), .B1(D15605_Y),     .Y(D15604_Y), .A0(D15606_Y));
KC_AOI22_X1 D15601 ( .A1(D15348_Y), .B0(D15345_Y), .B1(D15602_Y),     .Y(D15601_Y), .A0(D15603_Y));
KC_AOI22_X1 D15541 ( .A1(D15558_Y), .B0(D755_Y), .B1(D15557_Y),     .Y(D15541_Y), .A0(D14750_Y));
KC_AOI22_X1 D15536 ( .A1(D14749_Y), .B0(D15349_Y), .B1(D15525_Y),     .Y(D15536_Y), .A0(D15378_Y));
KC_AOI22_X1 D15535 ( .A1(D15348_Y), .B0(D15349_Y), .B1(D15526_Y),     .Y(D15535_Y), .A0(D15559_Y));
KC_AOI22_X1 D15527 ( .A1(D15800_Y), .B0(D15522_Y), .B1(D15438_Y),     .Y(D15527_Y), .A0(D15563_Y));
KC_AOI22_X1 D15521 ( .A1(D14396_Y), .B0(D15522_Y), .B1(D2871_Y),     .Y(D15521_Y), .A0(D15563_Y));
KC_AOI22_X1 D15520 ( .A1(D15800_Y), .B0(D15522_Y), .B1(D8889_Y),     .Y(D15520_Y), .A0(D15563_Y));
KC_AOI22_X1 D15519 ( .A1(D14181_Y), .B0(D15522_Y), .B1(D8886_Y),     .Y(D15519_Y), .A0(D15563_Y));
KC_AOI22_X1 D15518 ( .A1(D14314_Y), .B0(D15522_Y), .B1(D8902_Y),     .Y(D15518_Y), .A0(D15563_Y));
KC_AOI22_X1 D15515 ( .A1(D15426_Y), .B0(D755_Y), .B1(D15558_Y),     .Y(D15515_Y), .A0(D14750_Y));
KC_AOI22_X1 D15514 ( .A1(D15146_Y), .B0(D15522_Y), .B1(D9553_Y),     .Y(D15514_Y), .A0(D16461_Y));
KC_AOI22_X1 D15513 ( .A1(D15806_Y), .B0(D15522_Y), .B1(D8997_Y),     .Y(D15513_Y), .A0(D16461_Y));
KC_AOI22_X1 D15512 ( .A1(D15877_Y), .B0(D15522_Y), .B1(D6524_Y),     .Y(D15512_Y), .A0(D15563_Y));
KC_AOI22_X1 D15511 ( .A1(D15557_Y), .B0(D755_Y), .B1(D15556_Y),     .Y(D15511_Y), .A0(D14750_Y));
KC_AOI22_X1 D15510 ( .A1(D15556_Y), .B0(D755_Y), .B1(D15415_Y),     .Y(D15510_Y), .A0(D14750_Y));
KC_AOI22_X1 D15504 ( .A1(D16270_Y), .B0(D15969_Y), .B1(D15503_Y),     .Y(D15504_Y), .A0(D15505_Y));
KC_AOI22_X1 D15499 ( .A1(D15969_Y), .B0(D16270_Y), .B1(D15503_Y),     .Y(D15499_Y), .A0(D15500_Y));
KC_AOI22_X1 D15486 ( .A1(D15622_Y), .B0(D2616_Y), .B1(D15620_Y),     .Y(D15486_Y), .A0(D15485_Y));
KC_AOI22_X1 D15401 ( .A1(D14749_Y), .B0(D15349_Y), .B1(D15538_Y),     .Y(D15401_Y), .A0(D15365_Y));
KC_AOI22_X1 D15400 ( .A1(D15404_Y), .B0(D15359_Y), .B1(D771_Y),     .Y(D15400_Y), .A0(D15353_Y));
KC_AOI22_X1 D15399 ( .A1(D15528_Y), .B0(D15352_Y), .B1(D15517_Y),     .Y(D15399_Y), .A0(D15359_Y));
KC_AOI22_X1 D15398 ( .A1(D15359_Y), .B0(D15365_Y), .B1(D15551_Y),     .Y(D15398_Y), .A0(D15539_Y));
KC_AOI22_X1 D15393 ( .A1(D1188_Y), .B0(D2508_Y), .B1(D8888_Y),     .Y(D15393_Y), .A0(D13400_Y));
KC_AOI22_X1 D15381 ( .A1(D15055_Y), .B0(D2508_Y), .B1(D9085_Y),     .Y(D15381_Y), .A0(D13400_Y));
KC_AOI22_X1 D15370 ( .A1(D15512_Y), .B0(D15354_Y), .B1(D15514_Y),     .Y(D15370_Y), .A0(D15378_Y));
KC_AOI22_X1 D15368 ( .A1(D15521_Y), .B0(D15559_Y), .B1(D15354_Y),     .Y(D15368_Y), .A0(D15367_Y));
KC_AOI22_X1 D15358 ( .A1(D15518_Y), .B0(D15359_Y), .B1(D15384_Y),     .Y(D15358_Y), .A0(D15365_Y));
KC_AOI22_X1 D15356 ( .A1(D15346_Y), .B0(D15357_Y), .B1(D15376_Y),     .Y(D15356_Y), .A0(D15354_Y));
KC_AOI22_X1 D15347 ( .A1(D15523_Y), .B0(D15352_Y), .B1(D15355_Y),     .Y(D15347_Y), .A0(D15353_Y));
KC_AOI22_X1 D15343 ( .A1(D15346_Y), .B0(D15348_Y), .B1(D15523_Y),     .Y(D15343_Y), .A0(D15345_Y));
KC_AOI22_X1 D15342 ( .A1(D15525_Y), .B0(D15404_Y), .B1(D15364_Y),     .Y(D15342_Y), .A0(D15353_Y));
KC_AOI22_X1 D15222 ( .A1(D1072_Y), .B0(D16008_Q), .B1(D13710_Y),     .Y(D15222_Y), .A0(D1377_Q));
KC_AOI22_X1 D15221 ( .A1(D1072_Y), .B0(D1380_Q), .B1(D13710_Y),     .Y(D15221_Y), .A0(D15229_Q));
KC_AOI22_X1 D15181 ( .A1(D13636_Y), .B0(D15235_Q), .B1(D1073_Y),     .Y(D15181_Y), .A0(D15212_Q));
KC_AOI22_X1 D15179 ( .A1(D14176_Y), .B0(D1377_Q), .B1(D14259_Y),     .Y(D15179_Y), .A0(D16009_Q));
KC_AOI22_X1 D15178 ( .A1(D14257_Y), .B0(D15217_Q), .B1(D14254_Y),     .Y(D15178_Y), .A0(D1384_Q));
KC_AOI22_X1 D15177 ( .A1(D13640_Y), .B0(D15237_Q), .B1(D2476_Y),     .Y(D15177_Y), .A0(D15217_Q));
KC_AOI22_X1 D15175 ( .A1(D14256_Y), .B0(D1386_Q), .B1(D14172_Y),     .Y(D15175_Y), .A0(D15218_Q));
KC_AOI22_X1 D15174 ( .A1(D14256_Y), .B0(D15235_Q), .B1(D14172_Y),     .Y(D15174_Y), .A0(D15215_Q));
KC_AOI22_X1 D15173 ( .A1(D13635_Y), .B0(D15236_Q), .B1(D2477_Y),     .Y(D15173_Y), .A0(D15218_Q));
KC_AOI22_X1 D15169 ( .A1(D14176_Y), .B0(D15229_Q), .B1(D14259_Y),     .Y(D15169_Y), .A0(D15230_Q));
KC_AOI22_X1 D15168 ( .A1(D14176_Y), .B0(D1376_Q), .B1(D14259_Y),     .Y(D15168_Y), .A0(D15234_Q));
KC_AOI22_X1 D15167 ( .A1(D13635_Y), .B0(D16014_Q), .B1(D2477_Y),     .Y(D15167_Y), .A0(D15215_Q));
KC_AOI22_X1 D15163 ( .A1(D13634_Y), .B0(D15993_Q), .B1(D1071_Y),     .Y(D15163_Y), .A0(D1326_Q));
KC_AOI22_X1 D15162 ( .A1(D13634_Y), .B0(D1384_Q), .B1(D1071_Y),     .Y(D15162_Y), .A0(D15213_Q));
KC_AOI22_X1 D15160 ( .A1(D1072_Y), .B0(D15238_Q), .B1(D13710_Y),     .Y(D15160_Y), .A0(D1376_Q));
KC_AOI22_X1 D15109 ( .A1(D14256_Y), .B0(D16012_Q), .B1(D14172_Y),     .Y(D15109_Y), .A0(D1327_Q));
KC_AOI22_X1 D15108 ( .A1(D13635_Y), .B0(D16011_Q), .B1(D2477_Y),     .Y(D15108_Y), .A0(D1327_Q));
KC_AOI22_X1 D15104 ( .A1(D14255_Y), .B0(D15237_Q), .B1(D14252_Y),     .Y(D15104_Y), .A0(D15238_Q));
KC_AOI22_X1 D15103 ( .A1(D14440_Y), .B0(D15238_Q), .B1(D15107_Y),     .Y(D15103_Y), .A0(D14495_Q));
KC_AOI22_X1 D15097 ( .A1(D13526_Y), .B0(D16009_Q), .B1(D13510_Y),     .Y(D15097_Y), .A0(D15134_Q));
KC_AOI22_X1 D15093 ( .A1(D14173_Y), .B0(D1230_Q), .B1(D14171_Y),     .Y(D15093_Y), .A0(D15134_Q));
KC_AOI22_X1 D15090 ( .A1(D13635_Y), .B0(D16385_Q), .B1(D2477_Y),     .Y(D15090_Y), .A0(D15133_Q));
KC_AOI22_X1 D15088 ( .A1(D14256_Y), .B0(D15996_Q), .B1(D14255_Y),     .Y(D15088_Y), .A0(D15133_Q));
KC_AOI22_X1 D15087 ( .A1(D14255_Y), .B0(D16013_Q), .B1(D14252_Y),     .Y(D15087_Y), .A0(D16008_Q));
KC_AOI22_X1 D15086 ( .A1(D14258_Y), .B0(D15231_Q), .B1(D2519_Y),     .Y(D15086_Y), .A0(D15236_Q));
KC_AOI22_X1 D15085 ( .A1(D14258_Y), .B0(D15997_Q), .B1(D2519_Y),     .Y(D15085_Y), .A0(D16011_Q));
KC_AOI22_X1 D15045 ( .A1(D1072_Y), .B0(D15996_Q), .B1(D13710_Y),     .Y(D15045_Y), .A0(D2572_Q));
KC_AOI22_X1 D15044 ( .A1(D13526_Y), .B0(D1231_Q), .B1(D13510_Y),     .Y(D15044_Y), .A0(D1158_Q));
KC_AOI22_X1 D15043 ( .A1(D14256_Y), .B0(D16365_Q), .B1(D14255_Y),     .Y(D15043_Y), .A0(D1153_Q));
KC_AOI22_X1 D15040 ( .A1(D14256_Y), .B0(D15871_Q), .B1(D14255_Y),     .Y(D15040_Y), .A0(D15084_Q));
KC_AOI22_X1 D15036 ( .A1(D14256_Y), .B0(D14304_Q), .B1(D14255_Y),     .Y(D15036_Y), .A0(D1048_Q));
KC_AOI22_X1 D15035 ( .A1(D14171_Y), .B0(D14876_Q), .B1(D14144_Y),     .Y(D15035_Y), .A0(D2638_Q));
KC_AOI22_X1 D15034 ( .A1(D14171_Y), .B0(D14169_Q), .B1(D14144_Y),     .Y(D15034_Y), .A0(D15868_Q));
KC_AOI22_X1 D15033 ( .A1(D14171_Y), .B0(D14877_Q), .B1(D14144_Y),     .Y(D15033_Y), .A0(D15948_Q));
KC_AOI22_X1 D15030 ( .A1(D14173_Y), .B0(D16354_Q), .B1(D2519_Y),     .Y(D15030_Y), .A0(D1157_Q));
KC_AOI22_X1 D15029 ( .A1(D14258_Y), .B0(D2517_Q), .B1(D14145_Y),     .Y(D15029_Y), .A0(D16393_Q));
KC_AOI22_X1 D15028 ( .A1(D14258_Y), .B0(D14787_Q), .B1(D14145_Y),     .Y(D15028_Y), .A0(D16385_Q));
KC_AOI22_X1 D15027 ( .A1(D13526_Y), .B0(D1154_Q), .B1(D13510_Y),     .Y(D15027_Y), .A0(D1157_Q));
KC_AOI22_X1 D15026 ( .A1(D14258_Y), .B0(D14091_Q), .B1(D14145_Y),     .Y(D15026_Y), .A0(D16356_Q));
KC_AOI22_X1 D15023 ( .A1(D14176_Y), .B0(D1163_Q), .B1(D14259_Y),     .Y(D15023_Y), .A0(D1154_Q));
KC_AOI22_X1 D15021 ( .A1(D1072_Y), .B0(D15871_Q), .B1(D13710_Y),     .Y(D15021_Y), .A0(D1163_Q));
KC_AOI22_X1 D15020 ( .A1(D13635_Y), .B0(D16356_Q), .B1(D2477_Y),     .Y(D15020_Y), .A0(D15084_Q));
KC_AOI22_X1 D15017 ( .A1(D14173_Y), .B0(D16391_Q), .B1(D2519_Y),     .Y(D15017_Y), .A0(D1151_Q));
KC_AOI22_X1 D15016 ( .A1(D13635_Y), .B0(D16393_Q), .B1(D2477_Y),     .Y(D15016_Y), .A0(D1153_Q));
KC_AOI22_X1 D15015 ( .A1(D14173_Y), .B0(D15995_Q), .B1(D2519_Y),     .Y(D15015_Y), .A0(D1158_Q));
KC_AOI22_X1 D15013 ( .A1(D13526_Y), .B0(D2678_Q), .B1(D13510_Y),     .Y(D15013_Y), .A0(D1151_Q));
KC_AOI22_X1 D15011 ( .A1(D14176_Y), .B0(D14300_Q), .B1(D14259_Y),     .Y(D15011_Y), .A0(D2678_Q));
KC_AOI22_X1 D15010 ( .A1(D1072_Y), .B0(D16365_Q), .B1(D13710_Y),     .Y(D15010_Y), .A0(D14300_Q));
KC_AOI22_X1 D15007 ( .A1(D16365_Q), .B0(D14997_Q), .B1(D15009_Y),     .Y(D15007_Y), .A0(D15008_Y));
KC_AOI22_X1 D14957 ( .A1(D14175_Y), .B0(D2639_Q), .B1(D14174_Y),     .Y(D14957_Y), .A0(D14903_Q));
KC_AOI22_X1 D14956 ( .A1(D14173_Y), .B0(D1074_Q), .B1(D2519_Y),     .Y(D14956_Y), .A0(D14875_Q));
KC_AOI22_X1 D14955 ( .A1(D14173_Y), .B0(D16318_Q), .B1(D2519_Y),     .Y(D14955_Y), .A0(D14873_Q));
KC_AOI22_X1 D14953 ( .A1(D13636_Y), .B0(D14874_Q), .B1(D1073_Y),     .Y(D14953_Y), .A0(D14903_Q));
KC_AOI22_X1 D14951 ( .A1(D14176_Y), .B0(D1052_Q), .B1(D14259_Y),     .Y(D14951_Y), .A0(D14870_Q));
KC_AOI22_X1 D14950 ( .A1(D13635_Y), .B0(D2641_Q), .B1(D2477_Y),     .Y(D14950_Y), .A0(D14266_Q));
KC_AOI22_X1 D14949 ( .A1(D1072_Y), .B0(D1054_Q), .B1(D13710_Y),     .Y(D14949_Y), .A0(D1065_Q));
KC_AOI22_X1 D14948 ( .A1(D14256_Y), .B0(D1054_Q), .B1(D14255_Y),     .Y(D14948_Y), .A0(D14266_Q));
KC_AOI22_X1 D14944 ( .A1(D1072_Y), .B0(D14997_Q), .B1(D13710_Y),     .Y(D14944_Y), .A0(D1052_Q));
KC_AOI22_X1 D14943 ( .A1(D14256_Y), .B0(D14997_Q), .B1(D14255_Y),     .Y(D14943_Y), .A0(D14995_Q));
KC_AOI22_X1 D14942 ( .A1(D14172_Y), .B0(D145_Q), .B1(D14252_Y),     .Y(D14942_Y), .A0(D14874_Q));
KC_AOI22_X1 D14939 ( .A1(D13710_Y), .B0(D1051_Q), .B1(D1072_Y),     .Y(D14939_Y), .A0(D16314_Q));
KC_AOI22_X1 D14938 ( .A1(D13635_Y), .B0(D15669_Q), .B1(D2477_Y),     .Y(D14938_Y), .A0(D14995_Q));
KC_AOI22_X1 D14937 ( .A1(D14176_Y), .B0(D1051_Q), .B1(D14259_Y),     .Y(D14937_Y), .A0(D15794_Q));
KC_AOI22_X1 D14931 ( .A1(D14256_Y), .B0(D16314_Q), .B1(D14255_Y),     .Y(D14931_Y), .A0(D14996_Q));
KC_AOI22_X1 D14930 ( .A1(D2477_Y), .B0(D14996_Q), .B1(D13635_Y),     .Y(D14930_Y), .A0(D14872_Q));
KC_AOI22_X1 D14919 ( .A1(D14173_Y), .B0(D16361_Q), .B1(D2519_Y),     .Y(D14919_Y), .A0(D14263_Q));
KC_AOI22_X1 D14918 ( .A1(D13510_Y), .B0(D14263_Q), .B1(D13526_Y),     .Y(D14918_Y), .A0(D2516_Q));
KC_AOI22_X1 D14917 ( .A1(D14258_Y), .B0(D14118_Q), .B1(D14145_Y),     .Y(D14917_Y), .A0(D2679_Q));
KC_AOI22_X1 D14914 ( .A1(D14176_Y), .B0(D143_Q), .B1(D14259_Y),     .Y(D14914_Y), .A0(D2516_Q));
KC_AOI22_X1 D14913 ( .A1(D14171_Y), .B0(D14168_Q), .B1(D14144_Y),     .Y(D14913_Y), .A0(D15873_Q));
KC_AOI22_X1 D14910 ( .A1(D2573_Q), .B0(D2517_Q), .B1(D14912_Y),     .Y(D14910_Y), .A0(D14911_Y));
KC_AOI22_X1 D14845 ( .A1(D15000_Y), .B0(D14813_Y), .B1(D12139_Y),     .Y(D14845_Y), .A0(D15562_Y));
KC_AOI22_X1 D14841 ( .A1(D14392_Y), .B0(D14813_Y), .B1(D10205_Y),     .Y(D14841_Y), .A0(D15562_Y));
KC_AOI22_X1 D14839 ( .A1(D15000_Y), .B0(D14813_Y), .B1(D6111_Y),     .Y(D14839_Y), .A0(D15562_Y));
KC_AOI22_X1 D14838 ( .A1(D14146_Y), .B0(D14789_Q), .B1(D14147_Y),     .Y(D14838_Y), .A0(D14788_Q));
KC_AOI22_X1 D14834 ( .A1(D14258_Y), .B0(D14815_Q), .B1(D14145_Y),     .Y(D14834_Y), .A0(D14872_Q));
KC_AOI22_X1 D14833 ( .A1(D14171_Y), .B0(D14170_Q), .B1(D14144_Y),     .Y(D14833_Y), .A0(D14871_Q));
KC_AOI22_X1 D14832 ( .A1(D14171_Y), .B0(D14878_Q), .B1(D14144_Y),     .Y(D14832_Y), .A0(D15668_Q));
KC_AOI22_X1 D14831 ( .A1(D14171_Y), .B0(D2573_Q), .B1(D14144_Y),     .Y(D14831_Y), .A0(D15791_Q));
KC_AOI22_X1 D14825 ( .A1(D14146_Y), .B0(D14790_Q), .B1(D14147_Y),     .Y(D14825_Y), .A0(D820_Q));
KC_AOI22_X1 D14824 ( .A1(D14147_Y), .B0(D856_Q), .B1(D14146_Y),     .Y(D14824_Y), .A0(D14094_Q));
KC_AOI22_X1 D14823 ( .A1(D14147_Y), .B0(D818_Q), .B1(D14146_Y),     .Y(D14823_Y), .A0(D853_Q));
KC_AOI22_X1 D14822 ( .A1(D14146_Y), .B0(D815_Q), .B1(D14147_Y),     .Y(D14822_Y), .A0(D14808_Q));
KC_AOI22_X1 D14819 ( .A1(D14258_Y), .B0(D14117_Q), .B1(D14145_Y),     .Y(D14819_Y), .A0(D2641_Q));
KC_AOI22_X1 D14818 ( .A1(D14258_Y), .B0(D14814_Q), .B1(D14145_Y),     .Y(D14818_Y), .A0(D15669_Q));
KC_AOI22_X1 D14816 ( .A1(D13510_Y), .B0(D14873_Q), .B1(D13526_Y),     .Y(D14816_Y), .A0(D15794_Q));
KC_AOI22_X1 D14752 ( .A1(D15111_Y), .B0(D2508_Y), .B1(D12139_Y),     .Y(D14752_Y), .A0(D13400_Y));
KC_AOI22_X1 D14751 ( .A1(D14114_Y), .B0(D14113_Y), .B1(D14679_Y),     .Y(D14751_Y), .A0(D11228_Y));
KC_AOI22_X1 D14749 ( .A1(D14380_Y), .B0(D15522_Y), .B1(D15437_Y),     .Y(D14749_Y), .A0(D15563_Y));
KC_AOI22_X1 D14746 ( .A1(D2501_Y), .B0(D2508_Y), .B1(D16166_Y),     .Y(D14746_Y), .A0(D13400_Y));
KC_AOI22_X1 D14741 ( .A1(D15122_Y), .B0(D2508_Y), .B1(D2870_Y),     .Y(D14741_Y), .A0(D13400_Y));
KC_AOI22_X1 D14740 ( .A1(D14114_Y), .B0(D14113_Y), .B1(D15322_Y),     .Y(D14740_Y), .A0(D10797_Y));
KC_AOI22_X1 D14739 ( .A1(D14114_Y), .B0(D14113_Y), .B1(D508_Y),     .Y(D14739_Y), .A0(D10751_Y));
KC_AOI22_X1 D14738 ( .A1(D14114_Y), .B0(D14113_Y), .B1(D14515_Y),     .Y(D14738_Y), .A0(D12319_Y));
KC_AOI22_X1 D14737 ( .A1(D14976_Y), .B0(D2508_Y), .B1(D651_Y),     .Y(D14737_Y), .A0(D13400_Y));
KC_AOI22_X1 D14733 ( .A1(D14022_Y), .B0(D14679_Y), .B1(D14009_Y),     .Y(D14733_Y), .A0(D14790_Q));
KC_AOI22_X1 D14732 ( .A1(D14022_Y), .B0(D14515_Y), .B1(D14009_Y),     .Y(D14732_Y), .A0(D14789_Q));
KC_AOI22_X1 D14729 ( .A1(D14022_Y), .B0(D15322_Y), .B1(D14009_Y),     .Y(D14729_Y), .A0(D853_Q));
KC_AOI22_X1 D14724 ( .A1(D14138_Y), .B0(D14515_Y), .B1(D14130_Y),     .Y(D14724_Y), .A0(D14877_Q));
KC_AOI22_X1 D14723 ( .A1(D14010_Y), .B0(D14679_Y), .B1(D2496_Y),     .Y(D14723_Y), .A0(D2517_Q));
KC_AOI22_X1 D14722 ( .A1(D14010_Y), .B0(D15322_Y), .B1(D2496_Y),     .Y(D14722_Y), .A0(D14814_Q));
KC_AOI22_X1 D14721 ( .A1(D14010_Y), .B0(D508_Y), .B1(D2496_Y),     .Y(D14721_Y), .A0(D14815_Q));
KC_AOI22_X1 D14717 ( .A1(D14022_Y), .B0(D508_Y), .B1(D14009_Y),     .Y(D14717_Y), .A0(D815_Q));
KC_AOI22_X1 D14716 ( .A1(D14010_Y), .B0(D14515_Y), .B1(D2496_Y),     .Y(D14716_Y), .A0(D14787_Q));
KC_AOI22_X1 D14626 ( .A1(D14962_Y), .B0(D2508_Y), .B1(D6111_Y),     .Y(D14626_Y), .A0(D13400_Y));
KC_AOI22_X1 D14657 ( .A1(D14975_Y), .B0(D2508_Y), .B1(D8885_Y),     .Y(D14657_Y), .A0(D13400_Y));
KC_AOI22_X1 D14648 ( .A1(D14661_Y), .B0(D14662_Y), .B1(D14649_Y),     .Y(D14648_Y), .A0(D14650_Y));
KC_AOI22_X1 D14647 ( .A1(D15443_Y), .B0(D14656_Y), .B1(D15453_Y),     .Y(D14647_Y), .A0(D14656_Y));
KC_AOI22_X1 D14645 ( .A1(D14627_Y), .B0(D14655_Y), .B1(D14588_Y),     .Y(D14645_Y), .A0(D14742_Y));
KC_AOI22_X1 D14633 ( .A1(D15061_Y), .B0(D2508_Y), .B1(D8998_Y),     .Y(D14633_Y), .A0(D13400_Y));
KC_AOI22_X1 D14623 ( .A1(D14964_Y), .B0(D2508_Y), .B1(D16198_Y),     .Y(D14623_Y), .A0(D13400_Y));
KC_AOI22_X1 D14555 ( .A1(D14536_Y), .B0(D14529_Y), .B1(D14544_Y),     .Y(D14555_Y), .A0(D12278_Q));
KC_AOI22_X1 D14554 ( .A1(D14582_Y), .B0(D605_Q), .B1(D14536_Y),     .Y(D14554_Y), .A0(D2512_Y));
KC_AOI22_X1 D14551 ( .A1(D14536_Y), .B0(D14655_Y), .B1(D13912_Y),     .Y(D14551_Y), .A0(D12236_Q));
KC_AOI22_X1 D14550 ( .A1(D14581_Y), .B0(D14655_Y), .B1(D12218_Y),     .Y(D14550_Y), .A0(D2574_Q));
KC_AOI22_X1 D14538 ( .A1(D14736_Y), .B0(D14655_Y), .B1(D13911_Y),     .Y(D14538_Y), .A0(D12235_Q));
KC_AOI22_X1 D14537 ( .A1(D14736_Y), .B0(D14655_Y), .B1(D14590_Y),     .Y(D14537_Y), .A0(D12234_Q));
KC_AOI22_X1 D14533 ( .A1(D14736_Y), .B0(D14655_Y), .B1(D14592_Y),     .Y(D14533_Y), .A0(D12237_Q));
KC_AOI22_X1 D14482 ( .A1(D14487_Y), .B0(D1380_Q), .B1(D15161_Y),     .Y(D14482_Y), .A0(D14480_Y));
KC_AOI22_X1 D14450 ( .A1(D13636_Y), .B0(D14492_Q), .B1(D1073_Y),     .Y(D14450_Y), .A0(D14475_Q));
KC_AOI22_X1 D14449 ( .A1(D13634_Y), .B0(D14491_Q), .B1(D1071_Y),     .Y(D14449_Y), .A0(D13807_Q));
KC_AOI22_X1 D14448 ( .A1(D14464_Y), .B0(D15235_Q), .B1(D14453_Y),     .Y(D14448_Y), .A0(D14410_Y));
KC_AOI22_X1 D14447 ( .A1(D13636_Y), .B0(D1386_Q), .B1(D1073_Y),     .Y(D14447_Y), .A0(D1323_Q));
KC_AOI22_X1 D14442 ( .A1(D14460_Y), .B0(D14496_Q), .B1(D14417_Y),     .Y(D14442_Y), .A0(D14406_Y));
KC_AOI22_X1 D14434 ( .A1(D14256_Y), .B0(D14492_Q), .B1(D14172_Y),     .Y(D14434_Y), .A0(D13771_Q));
KC_AOI22_X1 D14433 ( .A1(D14370_Y), .B0(D16014_Q), .B1(D14438_Y),     .Y(D14433_Y), .A0(D14432_Y));
KC_AOI22_X1 D14429 ( .A1(D1072_Y), .B0(D1401_Q), .B1(D13710_Y),     .Y(D14429_Y), .A0(D13804_Q));
KC_AOI22_X1 D14428 ( .A1(D13634_Y), .B0(D14493_Q), .B1(D1071_Y),     .Y(D14428_Y), .A0(D15232_Q));
KC_AOI22_X1 D14426 ( .A1(D14257_Y), .B0(D15214_Q), .B1(D14254_Y),     .Y(D14426_Y), .A0(D14493_Q));
KC_AOI22_X1 D14425 ( .A1(D14253_Y), .B0(D14496_Q), .B1(D936_Y),     .Y(D14425_Y), .A0(D15232_Q));
KC_AOI22_X1 D14423 ( .A1(D14257_Y), .B0(D13816_Q), .B1(D14254_Y),     .Y(D14423_Y), .A0(D14491_Q));
KC_AOI22_X1 D14422 ( .A1(D14253_Y), .B0(D13808_Q), .B1(D936_Y),     .Y(D14422_Y), .A0(D1321_Q));
KC_AOI22_X1 D14421 ( .A1(D14176_Y), .B0(D14490_Q), .B1(D14259_Y),     .Y(D14421_Y), .A0(D1382_Q));
KC_AOI22_X1 D14420 ( .A1(D14257_Y), .B0(D13815_Q), .B1(D14254_Y),     .Y(D14420_Y), .A0(D14494_Q));
KC_AOI22_X1 D14416 ( .A1(D13524_Y), .B0(D14496_Q), .B1(D14224_Y),     .Y(D14416_Y), .A0(D15216_Q));
KC_AOI22_X1 D14411 ( .A1(D13524_Y), .B0(D13808_Q), .B1(D14224_Y),     .Y(D14411_Y), .A0(D13814_Q));
KC_AOI22_X1 D14409 ( .A1(D13640_Y), .B0(D1383_Q), .B1(D2476_Y),     .Y(D14409_Y), .A0(D15214_Q));
KC_AOI22_X1 D14402 ( .A1(D13634_Y), .B0(D14494_Q), .B1(D1071_Y),     .Y(D14402_Y), .A0(D1321_Q));
KC_AOI22_X1 D14401 ( .A1(D14463_Y), .B0(D14493_Q), .B1(D1268_Y),     .Y(D14401_Y), .A0(D14427_Y));
KC_AOI22_X1 D14398 ( .A1(D1072_Y), .B0(D14495_Q), .B1(D13710_Y),     .Y(D14398_Y), .A0(D14490_Q));
KC_AOI22_X1 D14357 ( .A1(D14255_Y), .B0(D13826_Q), .B1(D14252_Y),     .Y(D14357_Y), .A0(D14495_Q));
KC_AOI22_X1 D14347 ( .A1(D13526_Y), .B0(D15234_Q), .B1(D13510_Y),     .Y(D14347_Y), .A0(D2524_Q));
KC_AOI22_X1 D14346 ( .A1(D13526_Y), .B0(D15230_Q), .B1(D13510_Y),     .Y(D14346_Y), .A0(D2523_Q));
KC_AOI22_X1 D14345 ( .A1(D14362_Y), .B0(D15230_Q), .B1(D14350_Y),     .Y(D14345_Y), .A0(D14351_Y));
KC_AOI22_X1 D14339 ( .A1(D14173_Y), .B0(D13762_Q), .B1(D14171_Y),     .Y(D14339_Y), .A0(D13764_Q));
KC_AOI22_X1 D14337 ( .A1(D14173_Y), .B0(D14374_Q), .B1(D14171_Y),     .Y(D14337_Y), .A0(D2523_Q));
KC_AOI22_X1 D14333 ( .A1(D14173_Y), .B0(D13761_Q), .B1(D14171_Y),     .Y(D14333_Y), .A0(D14375_Q));
KC_AOI22_X1 D14332 ( .A1(D14364_Y), .B0(D1379_Q), .B1(D14335_Y),     .Y(D14332_Y), .A0(D1182_Y));
KC_AOI22_X1 D14331 ( .A1(D14173_Y), .B0(D1232_Q), .B1(D14171_Y),     .Y(D14331_Y), .A0(D2524_Q));
KC_AOI22_X1 D14330 ( .A1(D13525_Y), .B0(D1379_Q), .B1(D2475_Y),     .Y(D14330_Y), .A0(D14374_Q));
KC_AOI22_X1 D14326 ( .A1(D14175_Y), .B0(D13809_Q), .B1(D14174_Y),     .Y(D14326_Y), .A0(D13811_Q));
KC_AOI22_X1 D14325 ( .A1(D14175_Y), .B0(D13814_Q), .B1(D14174_Y),     .Y(D14325_Y), .A0(D14475_Q));
KC_AOI22_X1 D14323 ( .A1(D14176_Y), .B0(D13804_Q), .B1(D14259_Y),     .Y(D14323_Y), .A0(D13812_Q));
KC_AOI22_X1 D14321 ( .A1(D14258_Y), .B0(D1379_Q), .B1(D2519_Y),     .Y(D14321_Y), .A0(D16014_Q));
KC_AOI22_X1 D14320 ( .A1(D14253_Y), .B0(D13806_Q), .B1(D936_Y),     .Y(D14320_Y), .A0(D13807_Q));
KC_AOI22_X1 D14319 ( .A1(D14256_Y), .B0(D13827_Q), .B1(D14172_Y),     .Y(D14319_Y), .A0(D13760_Q));
KC_AOI22_X1 D14318 ( .A1(D14175_Y), .B0(D1325_Q), .B1(D14174_Y),     .Y(D14318_Y), .A0(D1323_Q));
KC_AOI22_X1 D14317 ( .A1(D14175_Y), .B0(D15216_Q), .B1(D14174_Y),     .Y(D14317_Y), .A0(D15212_Q));
KC_AOI22_X1 D14284 ( .A1(D14257_Y), .B0(D164_Q), .B1(D14254_Y),     .Y(D14284_Y), .A0(D14298_Q));
KC_AOI22_X1 D14283 ( .A1(D14175_Y), .B0(D13705_Q), .B1(D14174_Y),     .Y(D14283_Y), .A0(D1150_Q));
KC_AOI22_X1 D14280 ( .A1(D14256_Y), .B0(D14306_Q), .B1(D14172_Y),     .Y(D14280_Y), .A0(D13050_Q));
KC_AOI22_X1 D14279 ( .A1(D14255_Y), .B0(D14307_Q), .B1(D14252_Y),     .Y(D14279_Y), .A0(D14302_Q));
KC_AOI22_X1 D14278 ( .A1(D14253_Y), .B0(D14303_Q), .B1(D936_Y),     .Y(D14278_Y), .A0(D1147_Q));
KC_AOI22_X1 D14273 ( .A1(D14173_Y), .B0(D1159_Q), .B1(D14171_Y),     .Y(D14273_Y), .A0(D13765_Q));
KC_AOI22_X1 D14272 ( .A1(D14256_Y), .B0(D14316_Q), .B1(D14172_Y),     .Y(D14272_Y), .A0(D2468_Q));
KC_AOI22_X1 D14271 ( .A1(D14258_Y), .B0(D14297_Q), .B1(D2519_Y),     .Y(D14271_Y), .A0(D14299_Q));
KC_AOI22_X1 D14219 ( .A1(D14253_Y), .B0(D926_Q), .B1(D936_Y),     .Y(D14219_Y), .A0(D12994_Q));
KC_AOI22_X1 D14218 ( .A1(D14176_Y), .B0(D12993_Q), .B1(D14259_Y),     .Y(D14218_Y), .A0(D14166_Q));
KC_AOI22_X1 D14217 ( .A1(D14258_Y), .B0(D14167_Q), .B1(D2519_Y),     .Y(D14217_Y), .A0(D14239_Q));
KC_AOI22_X1 D14215 ( .A1(D14254_Y), .B0(D14243_Q), .B1(D14257_Y),     .Y(D14215_Y), .A0(D12995_Q));
KC_AOI22_X1 D14214 ( .A1(D14259_Y), .B0(D14264_Q), .B1(D14176_Y),     .Y(D14214_Y), .A0(D12997_Q));
KC_AOI22_X1 D14213 ( .A1(D14257_Y), .B0(D12992_Q), .B1(D14254_Y),     .Y(D14213_Y), .A0(D14246_Q));
KC_AOI22_X1 D14211 ( .A1(D14256_Y), .B0(D14242_Q), .B1(D14172_Y),     .Y(D14211_Y), .A0(D12991_Q));
KC_AOI22_X1 D14210 ( .A1(D14255_Y), .B0(D14236_Q), .B1(D14252_Y),     .Y(D14210_Y), .A0(D14244_Q));
KC_AOI22_X1 D14209 ( .A1(D14255_Y), .B0(D14196_Q), .B1(D14252_Y),     .Y(D14209_Y), .A0(D14241_Q));
KC_AOI22_X1 D14206 ( .A1(D14258_Y), .B0(D14245_Q), .B1(D2519_Y),     .Y(D14206_Y), .A0(D1066_Q));
KC_AOI22_X1 D14199 ( .A1(D14175_Y), .B0(D13711_Q), .B1(D14174_Y),     .Y(D14199_Y), .A0(D13703_Q));
KC_AOI22_X1 D14198 ( .A1(D14258_Y), .B0(D14240_Q), .B1(D2519_Y),     .Y(D14198_Y), .A0(D14237_Q));
KC_AOI22_X1 D14178 ( .A1(D14138_Y), .B0(D14517_Y), .B1(D14130_Y),     .Y(D14178_Y), .A0(D14169_Q));
KC_AOI22_X1 D14140 ( .A1(D14138_Y), .B0(D15329_Y), .B1(D14130_Y),     .Y(D14140_Y), .A0(D14168_Q));
KC_AOI22_X1 D14135 ( .A1(D14138_Y), .B0(D15323_Y), .B1(D14130_Y),     .Y(D14135_Y), .A0(D14170_Q));
KC_AOI22_X1 D14125 ( .A1(D14147_Y), .B0(D14093_Q), .B1(D14146_Y),     .Y(D14125_Y), .A0(D14092_Q));
KC_AOI22_X1 D14121 ( .A1(D14173_Y), .B0(D954_Q), .B1(D14171_Y),     .Y(D14121_Y), .A0(D928_Q));
KC_AOI22_X1 D14119 ( .A1(D14173_Y), .B0(D12921_Q), .B1(D14171_Y),     .Y(D14119_Y), .A0(D14165_Q));
KC_AOI22_X1 D14102 ( .A1(D14038_Y), .B0(D14034_Y), .B1(D14106_Y),     .Y(D14102_Y), .A0(D14107_Y));
KC_AOI22_X1 D14101 ( .A1(D14038_Y), .B0(D14034_Y), .B1(D14108_Y),     .Y(D14101_Y), .A0(D14103_Y));
KC_AOI22_X1 D14100 ( .A1(D14038_Y), .B0(D14034_Y), .B1(D14104_Y),     .Y(D14100_Y), .A0(D14105_Y));
KC_AOI22_X1 D14096 ( .A1(D12686_Q), .B0(D14033_Y), .B1(D13209_Q),     .Y(D14096_Y), .A0(D14077_Y));
KC_AOI22_X1 D14042 ( .A1(D12688_Q), .B0(D14033_Y), .B1(D13906_Y),     .Y(D14042_Y), .A0(D14077_Y));
KC_AOI22_X1 D14041 ( .A1(D14363_Y), .B0(D2508_Y), .B1(D13156_Y),     .Y(D14041_Y), .A0(D13400_Y));
KC_AOI22_X1 D14040 ( .A1(D12681_Q), .B0(D14033_Y), .B1(D13203_Q),     .Y(D14040_Y), .A0(D14077_Y));
KC_AOI22_X1 D14039 ( .A1(D2499_Y), .B0(D2508_Y), .B1(D10205_Y),     .Y(D14039_Y), .A0(D13400_Y));
KC_AOI22_X1 D14037 ( .A1(D14033_Y), .B0(D13279_Q), .B1(D14077_Y),     .Y(D14037_Y), .A0(D13976_Y));
KC_AOI22_X1 D14036 ( .A1(D12682_Q), .B0(D14033_Y), .B1(D12689_Q),     .Y(D14036_Y), .A0(D14077_Y));
KC_AOI22_X1 D14035 ( .A1(D12684_Q), .B0(D14033_Y), .B1(D13210_Q),     .Y(D14035_Y), .A0(D14077_Y));
KC_AOI22_X1 D14032 ( .A1(D13200_Q), .B0(D14033_Y), .B1(D2511_Y),     .Y(D14032_Y), .A0(D14077_Y));
KC_AOI22_X1 D14031 ( .A1(D14114_Y), .B0(D14113_Y), .B1(D15329_Y),     .Y(D14031_Y), .A0(D10291_Y));
KC_AOI22_X1 D14028 ( .A1(D14114_Y), .B0(D14113_Y), .B1(D14517_Y),     .Y(D14028_Y), .A0(D12320_Y));
KC_AOI22_X1 D14027 ( .A1(D14114_Y), .B0(D15323_Y), .B1(D14113_Y),     .Y(D14027_Y), .A0(D10794_Y));
KC_AOI22_X1 D14015 ( .A1(D14022_Y), .B0(D14517_Y), .B1(D14009_Y),     .Y(D14015_Y), .A0(D14094_Q));
KC_AOI22_X1 D14014 ( .A1(D14022_Y), .B0(D15329_Y), .B1(D14009_Y),     .Y(D14014_Y), .A0(D14109_Q));
KC_AOI22_X1 D14013 ( .A1(D14010_Y), .B0(D14517_Y), .B1(D2496_Y),     .Y(D14013_Y), .A0(D14091_Q));
KC_AOI22_X1 D14012 ( .A1(D14010_Y), .B0(D15323_Y), .B1(D2496_Y),     .Y(D14012_Y), .A0(D14117_Q));
KC_AOI22_X1 D14007 ( .A1(D14022_Y), .B0(D15323_Y), .B1(D14009_Y),     .Y(D14007_Y), .A0(D14092_Q));
KC_AOI22_X1 D13999 ( .A1(D13998_Q), .B0(D2461_Y), .B1(D13993_Q),     .Y(D13999_Y), .A0(D2462_Y));
KC_AOI22_X1 D13961 ( .A1(D13989_Q), .B0(D2509_Y), .B1(D6975_Y),     .Y(D13961_Y), .A0(D2462_Y));
KC_AOI22_X1 D13960 ( .A1(D13279_Q), .B0(D2461_Y), .B1(D696_Q),     .Y(D13960_Y), .A0(D2462_Y));
KC_AOI22_X1 D13959 ( .A1(D14365_Y), .B0(D2508_Y), .B1(D8887_Y),     .Y(D13959_Y), .A0(D13400_Y));
KC_AOI22_X1 D13954 ( .A1(D16125_Y), .B0(D13902_Y), .B1(D16200_Y),     .Y(D13954_Y), .A0(D13184_Y));
KC_AOI22_X1 D13949 ( .A1(D13272_Q), .B0(D2461_Y), .B1(D695_Q),     .Y(D13949_Y), .A0(D2462_Y));
KC_AOI22_X1 D13944 ( .A1(D13271_Q), .B0(D13281_Y), .B1(D13977_Y),     .Y(D13944_Y), .A0(D13254_Y));
KC_AOI22_X1 D13942 ( .A1(D13990_Q), .B0(D13281_Y), .B1(D13994_Q),     .Y(D13942_Y), .A0(D13254_Y));
KC_AOI22_X1 D13927 ( .A1(D14287_Y), .B0(D2508_Y), .B1(D9087_Y),     .Y(D13927_Y), .A0(D13400_Y));
KC_AOI22_X1 D13926 ( .A1(D13929_Y), .B0(D13930_Y), .B1(D13937_Y),     .Y(D13926_Y), .A0(D14044_Y));
KC_AOI22_X1 D13901 ( .A1(D13909_Q), .B0(D13955_Y), .B1(D14771_Y),     .Y(D13901_Y), .A0(D13904_Y));
KC_AOI22_X1 D13892 ( .A1(D13208_Q), .B0(D13281_Y), .B1(D2470_Y),     .Y(D13892_Y), .A0(D13254_Y));
KC_AOI22_X1 D13891 ( .A1(D13197_Q), .B0(D2461_Y), .B1(D2518_Q),     .Y(D13891_Y), .A0(D2462_Y));
KC_AOI22_X1 D13887 ( .A1(D12686_Q), .B0(D2461_Y), .B1(D13920_Q),     .Y(D13887_Y), .A0(D2462_Y));
KC_AOI22_X1 D13886 ( .A1(D13921_Q), .B0(D13955_Y), .B1(D14773_Y),     .Y(D13886_Y), .A0(D13904_Y));
KC_AOI22_X1 D13884 ( .A1(D12688_Q), .B0(D2461_Y), .B1(D13918_Q),     .Y(D13884_Y), .A0(D2462_Y));
KC_AOI22_X1 D13883 ( .A1(D12682_Q), .B0(D2461_Y), .B1(D13860_Q),     .Y(D13883_Y), .A0(D2462_Y));
KC_AOI22_X1 D13882 ( .A1(D13907_Q), .B0(D13955_Y), .B1(D14810_Y),     .Y(D13882_Y), .A0(D13904_Y));
KC_AOI22_X1 D13881 ( .A1(D12684_Q), .B0(D2461_Y), .B1(D619_Q),     .Y(D13881_Y), .A0(D2462_Y));
KC_AOI22_X1 D13877 ( .A1(D13195_Q), .B0(D2330_Y), .B1(D16080_Y),     .Y(D13877_Y), .A0(D13188_Y));
KC_AOI22_X1 D13876 ( .A1(D618_Q), .B0(D13955_Y), .B1(D14774_Y),     .Y(D13876_Y), .A0(D13904_Y));
KC_AOI22_X1 D13777 ( .A1(D13640_Y), .B0(D13810_Q), .B1(D2476_Y),     .Y(D13777_Y), .A0(D13816_Q));
KC_AOI22_X1 D13776 ( .A1(D13629_Y), .B0(D13826_Q), .B1(D2476_Y),     .Y(D13776_Y), .A0(D13815_Q));
KC_AOI22_X1 D13773 ( .A1(D13636_Y), .B0(D13827_Q), .B1(D1073_Y),     .Y(D13773_Y), .A0(D13811_Q));
KC_AOI22_X1 D13772 ( .A1(D13524_Y), .B0(D13806_Q), .B1(D14224_Y),     .Y(D13772_Y), .A0(D13809_Q));
KC_AOI22_X1 D13728 ( .A1(D13526_Y), .B0(D13812_Q), .B1(D13510_Y),     .Y(D13728_Y), .A0(D13764_Q));
KC_AOI22_X1 D13721 ( .A1(D13525_Y), .B0(D13759_Q), .B1(D2475_Y),     .Y(D13721_Y), .A0(D13761_Q));
KC_AOI22_X1 D13720 ( .A1(D13525_Y), .B0(D13813_Q), .B1(D2475_Y),     .Y(D13720_Y), .A0(D13762_Q));
KC_AOI22_X1 D13714 ( .A1(D13635_Y), .B0(D13805_Q), .B1(D2477_Y),     .Y(D13714_Y), .A0(D13760_Q));
KC_AOI22_X1 D13713 ( .A1(D13635_Y), .B0(D1375_Q), .B1(D2477_Y),     .Y(D13713_Y), .A0(D13771_Q));
KC_AOI22_X1 D13667 ( .A1(D13640_Y), .B0(D13770_Q), .B1(D2476_Y),     .Y(D13667_Y), .A0(D164_Q));
KC_AOI22_X1 D13661 ( .A1(D2332_Y), .B0(D14307_Q), .B1(D1091_Y),     .Y(D13661_Y), .A0(D12879_Y));
KC_AOI22_X1 D13660 ( .A1(D950_Y), .B0(D14303_Q), .B1(D2417_Y),     .Y(D13660_Y), .A0(D12879_Y));
KC_AOI22_X1 D13659 ( .A1(D949_Y), .B0(D14240_Q), .B1(D12939_Y),     .Y(D13659_Y), .A0(D12879_Y));
KC_AOI22_X1 D13648 ( .A1(D13636_Y), .B0(D14316_Q), .B1(D1073_Y),     .Y(D13648_Y), .A0(D1150_Q));
KC_AOI22_X1 D13647 ( .A1(D13524_Y), .B0(D2474_Q), .B1(D14224_Y),     .Y(D13647_Y), .A0(D13705_Q));
KC_AOI22_X1 D13643 ( .A1(D13635_Y), .B0(D14299_Q), .B1(D2477_Y),     .Y(D13643_Y), .A0(D2468_Q));
KC_AOI22_X1 D13642 ( .A1(D13525_Y), .B0(D14297_Q), .B1(D2475_Y),     .Y(D13642_Y), .A0(D1159_Q));
KC_AOI22_X1 D13551 ( .A1(D2371_Y), .B0(D12879_Y), .B1(D13027_Y),     .Y(D13551_Y), .A0(D13393_Y));
KC_AOI22_X1 D13577 ( .A1(D15774_Y), .B0(D13557_Y), .B1(D11276_Y),     .Y(D13577_Y), .A0(D14220_Y));
KC_AOI22_X1 D13576 ( .A1(D13558_Y), .B0(D13543_Y), .B1(D13601_Y),     .Y(D13576_Y), .A0(D12994_Q));
KC_AOI22_X1 D13575 ( .A1(D2401_Y), .B0(D12879_Y), .B1(D13699_Y),     .Y(D13575_Y), .A0(D13393_Y));
KC_AOI22_X1 D13565 ( .A1(D12950_Y), .B0(D12879_Y), .B1(D12970_Y),     .Y(D13565_Y), .A0(D13393_Y));
KC_AOI22_X1 D13463 ( .A1(D13459_Y), .B0(D2438_Y), .B1(D13503_Y),     .Y(D13463_Y), .A0(D13530_Q));
KC_AOI22_X1 D13453 ( .A1(D13457_Y), .B0(D13458_Y), .B1(D13498_Y),     .Y(D13453_Y), .A0(D14165_Q));
KC_AOI22_X1 D13440 ( .A1(D162_Y), .B0(D14305_Q), .B1(D13443_Y),     .Y(D13440_Y), .A0(D12879_Y));
KC_AOI22_X1 D13439 ( .A1(D13467_Y), .B0(D12879_Y), .B1(D13696_Y),     .Y(D13439_Y), .A0(D13393_Y));
KC_AOI22_X1 D13434 ( .A1(D12879_Y), .B0(D13393_Y), .B1(D13456_Y),     .Y(D13434_Y), .A0(D13512_Y));
KC_AOI22_X1 D13426 ( .A1(D13451_Y), .B0(D2435_Y), .B1(D13487_Y),     .Y(D13426_Y), .A0(D12921_Q));
KC_AOI22_X1 D13416 ( .A1(D13430_Y), .B0(D12879_Y), .B1(D13697_Y),     .Y(D13416_Y), .A0(D13393_Y));
KC_AOI22_X1 D13350 ( .A1(D12685_Q), .B0(D14033_Y), .B1(D13974_Y),     .Y(D13350_Y), .A0(D14077_Y));
KC_AOI22_X1 D13310 ( .A1(D13293_Y), .B0(D13378_Y), .B1(D13292_Y),     .Y(D13310_Y), .A0(D14019_Y));
KC_AOI22_X1 D13304 ( .A1(D13293_Y), .B0(D13292_Y), .B1(D13377_Y),     .Y(D13304_Y), .A0(D13318_Y));
KC_AOI22_X1 D13303 ( .A1(D2431_Y), .B0(D13378_Y), .B1(D13311_Y),     .Y(D13303_Y), .A0(D14019_Y));
KC_AOI22_X1 D13291 ( .A1(D2431_Y), .B0(D13377_Y), .B1(D13311_Y),     .Y(D13291_Y), .A0(D13318_Y));
KC_AOI22_X1 D13284 ( .A1(D12687_Q), .B0(D2461_Y), .B1(D13274_Q),     .Y(D13284_Y), .A0(D2462_Y));
KC_AOI22_X1 D13238 ( .A1(D13991_Q), .B0(D13281_Y), .B1(D693_Q),     .Y(D13238_Y), .A0(D13254_Y));
KC_AOI22_X1 D13237 ( .A1(D697_Q), .B0(D2461_Y), .B1(D13997_Q),     .Y(D13237_Y), .A0(D2462_Y));
KC_AOI22_X1 D13217 ( .A1(D692_Q), .B0(D13281_Y), .B1(D13216_Q),     .Y(D13217_Y), .A0(D13254_Y));
KC_AOI22_X1 D13182 ( .A1(D13200_Q), .B0(D2461_Y), .B1(D13201_Q),     .Y(D13182_Y), .A0(D2462_Y));
KC_AOI22_X1 D13181 ( .A1(D691_Q), .B0(D2461_Y), .B1(D13196_Q),     .Y(D13181_Y), .A0(D2462_Y));
KC_AOI22_X1 D13180 ( .A1(D13202_Q), .B0(D2461_Y), .B1(D13212_Q),     .Y(D13180_Y), .A0(D2462_Y));
KC_AOI22_X1 D13151 ( .A1(D11990_Y), .B0(D13148_Q), .B1(D12011_Y),     .Y(D13151_Y), .A0(D13143_Q));
KC_AOI22_X1 D13142 ( .A1(D13147_Q), .B0(D12010_Y), .B1(D13146_Q),     .Y(D13142_Y), .A0(D11438_Y));
KC_AOI22_X1 D13141 ( .A1(D1362_Q), .B0(D12010_Y), .B1(D1360_Q),     .Y(D13141_Y), .A0(D11438_Y));
KC_AOI22_X1 D13140 ( .A1(D11990_Y), .B0(D13146_Q), .B1(D12011_Y),     .Y(D13140_Y), .A0(D13147_Q));
KC_AOI22_X1 D13139 ( .A1(D13143_Q), .B0(D12010_Y), .B1(D13148_Q),     .Y(D13139_Y), .A0(D11438_Y));
KC_AOI22_X1 D13138 ( .A1(D11990_Y), .B0(D1359_Q), .B1(D12011_Y),     .Y(D13138_Y), .A0(D1361_Q));
KC_AOI22_X1 D13137 ( .A1(D11990_Y), .B0(D13802_Q), .B1(D12011_Y),     .Y(D13137_Y), .A0(D13820_Q));
KC_AOI22_X1 D13136 ( .A1(D11990_Y), .B0(D1360_Q), .B1(D12011_Y),     .Y(D13136_Y), .A0(D1362_Q));
KC_AOI22_X1 D13135 ( .A1(D13144_Q), .B0(D12010_Y), .B1(D13149_Q),     .Y(D13135_Y), .A0(D11438_Y));
KC_AOI22_X1 D13134 ( .A1(D11990_Y), .B0(D13149_Q), .B1(D12011_Y),     .Y(D13134_Y), .A0(D13144_Q));
KC_AOI22_X1 D13132 ( .A1(D12024_Y), .B0(D13120_Q), .B1(D12023_Y),     .Y(D13132_Y), .A0(D13116_Q));
KC_AOI22_X1 D13112 ( .A1(D12024_Y), .B0(D13118_Q), .B1(D12023_Y),     .Y(D13112_Y), .A0(D1306_Q));
KC_AOI22_X1 D13110 ( .A1(D2467_Q), .B0(D12025_Y), .B1(D2385_Q),     .Y(D13110_Y), .A0(D2301_Y));
KC_AOI22_X1 D13109 ( .A1(D1213_Q), .B0(D12025_Y), .B1(D13801_Q),     .Y(D13109_Y), .A0(D2301_Y));
KC_AOI22_X1 D13108 ( .A1(D12047_Y), .B0(D13801_Q), .B1(D12015_Y),     .Y(D13108_Y), .A0(D1213_Q));
KC_AOI22_X1 D13107 ( .A1(D130_Q), .B0(D12025_Y), .B1(D1305_Q),     .Y(D13107_Y), .A0(D2301_Y));
KC_AOI22_X1 D13106 ( .A1(D12047_Y), .B0(D1305_Q), .B1(D12015_Y),     .Y(D13106_Y), .A0(D130_Q));
KC_AOI22_X1 D13105 ( .A1(D12047_Y), .B0(D2385_Q), .B1(D12015_Y),     .Y(D13105_Y), .A0(D2467_Q));
KC_AOI22_X1 D13104 ( .A1(D12047_Y), .B0(D1307_Q), .B1(D12015_Y),     .Y(D13104_Y), .A0(D2384_Q));
KC_AOI22_X1 D13102 ( .A1(D1306_Q), .B0(D12051_Y), .B1(D13118_Q),     .Y(D13102_Y), .A0(D12050_Y));
KC_AOI22_X1 D13101 ( .A1(D13116_Q), .B0(D12051_Y), .B1(D13120_Q),     .Y(D13101_Y), .A0(D12050_Y));
KC_AOI22_X1 D13100 ( .A1(D1361_Q), .B0(D12010_Y), .B1(D1359_Q),     .Y(D13100_Y), .A0(D11438_Y));
KC_AOI22_X1 D13099 ( .A1(D13820_Q), .B0(D12010_Y), .B1(D13802_Q),     .Y(D13099_Y), .A0(D11438_Y));
KC_AOI22_X1 D13092 ( .A1(D13043_Q), .B0(D12051_Y), .B1(D13083_Q),     .Y(D13092_Y), .A0(D12050_Y));
KC_AOI22_X1 D13078 ( .A1(D13095_Q), .B0(D12012_Y), .B1(D13096_Q),     .Y(D13078_Y), .A0(D12052_Y));
KC_AOI22_X1 D13077 ( .A1(D12024_Y), .B0(D1217_Q), .B1(D12023_Y),     .Y(D13077_Y), .A0(D13080_Q));
KC_AOI22_X1 D13076 ( .A1(D12024_Y), .B0(D13083_Q), .B1(D12023_Y),     .Y(D13076_Y), .A0(D13043_Q));
KC_AOI22_X1 D13075 ( .A1(D13086_Q), .B0(D12012_Y), .B1(D13087_Q),     .Y(D13075_Y), .A0(D12052_Y));
KC_AOI22_X1 D13071 ( .A1(D12047_Y), .B0(D13799_Q), .B1(D12015_Y),     .Y(D13071_Y), .A0(D13756_Q));
KC_AOI22_X1 D13070 ( .A1(D13756_Q), .B0(D12025_Y), .B1(D13799_Q),     .Y(D13070_Y), .A0(D2301_Y));
KC_AOI22_X1 D13069 ( .A1(D13080_Q), .B0(D12051_Y), .B1(D1217_Q),     .Y(D13069_Y), .A0(D12050_Y));
KC_AOI22_X1 D13068 ( .A1(D12024_Y), .B0(D13081_Q), .B1(D12023_Y),     .Y(D13068_Y), .A0(D13088_Q));
KC_AOI22_X1 D13065 ( .A1(D16097_Q), .B0(D12051_Y), .B1(D1216_Q),     .Y(D13065_Y), .A0(D12050_Y));
KC_AOI22_X1 D13064 ( .A1(D13088_Q), .B0(D12051_Y), .B1(D13081_Q),     .Y(D13064_Y), .A0(D12050_Y));
KC_AOI22_X1 D13063 ( .A1(D12024_Y), .B0(D1216_Q), .B1(D12023_Y),     .Y(D13063_Y), .A0(D16097_Q));
KC_AOI22_X1 D13062 ( .A1(D12016_Y), .B0(D13045_Q), .B1(D12026_Y),     .Y(D13062_Y), .A0(D13044_Q));
KC_AOI22_X1 D13061 ( .A1(D12016_Y), .B0(D13087_Q), .B1(D12026_Y),     .Y(D13061_Y), .A0(D13086_Q));
KC_AOI22_X1 D13060 ( .A1(D12016_Y), .B0(D13096_Q), .B1(D12026_Y),     .Y(D13060_Y), .A0(D13095_Q));
KC_AOI22_X1 D13059 ( .A1(D13044_Q), .B0(D12012_Y), .B1(D13045_Q),     .Y(D13059_Y), .A0(D12052_Y));
KC_AOI22_X1 D13055 ( .A1(D13082_Q), .B0(D12012_Y), .B1(D1214_Q),     .Y(D13055_Y), .A0(D12052_Y));
KC_AOI22_X1 D13054 ( .A1(D12016_Y), .B0(D1214_Q), .B1(D12026_Y),     .Y(D13054_Y), .A0(D13082_Q));
KC_AOI22_X1 D13024 ( .A1(D13034_Q), .B0(D11991_Y), .B1(D13032_Q),     .Y(D13024_Y), .A0(D2277_Y));
KC_AOI22_X1 D13023 ( .A1(D11969_Y), .B0(D13035_Q), .B1(D11948_Y),     .Y(D13023_Y), .A0(D13041_Q));
KC_AOI22_X1 D13022 ( .A1(D11969_Y), .B0(D13038_Q), .B1(D11948_Y),     .Y(D13022_Y), .A0(D13040_Q));
KC_AOI22_X1 D13021 ( .A1(D11950_Y), .B0(D13039_Q), .B1(D11953_Y),     .Y(D13021_Y), .A0(D2388_Q));
KC_AOI22_X1 D13020 ( .A1(D2388_Q), .B0(D11952_Y), .B1(D13039_Q),     .Y(D13020_Y), .A0(D2272_Y));
KC_AOI22_X1 D13018 ( .A1(D12421_Y), .B0(D13663_Y), .B1(D2398_Y),     .Y(D13018_Y), .A0(D12879_Y));
KC_AOI22_X1 D13017 ( .A1(D13040_Q), .B0(D11991_Y), .B1(D13038_Q),     .Y(D13017_Y), .A0(D2277_Y));
KC_AOI22_X1 D13016 ( .A1(D12420_Y), .B0(D13662_Y), .B1(D2397_Y),     .Y(D13016_Y), .A0(D12879_Y));
KC_AOI22_X1 D13014 ( .A1(D13041_Q), .B0(D11991_Y), .B1(D13035_Q),     .Y(D13014_Y), .A0(D2277_Y));
KC_AOI22_X1 D13013 ( .A1(D11969_Y), .B0(D13031_Q), .B1(D11948_Y),     .Y(D13013_Y), .A0(D13033_Q));
KC_AOI22_X1 D13012 ( .A1(D13033_Q), .B0(D11991_Y), .B1(D13031_Q),     .Y(D13012_Y), .A0(D2277_Y));
KC_AOI22_X1 D12958 ( .A1(D11969_Y), .B0(D12986_Q), .B1(D11948_Y),     .Y(D12958_Y), .A0(D12985_Q));
KC_AOI22_X1 D12957 ( .A1(D11969_Y), .B0(D2389_Q), .B1(D11948_Y),     .Y(D12957_Y), .A0(D12987_Q));
KC_AOI22_X1 D12956 ( .A1(D13571_Y), .B0(D13567_Y), .B1(D12965_Y),     .Y(D12956_Y), .A0(D12996_Q));
KC_AOI22_X1 D12953 ( .A1(D13560_Y), .B0(D13548_Y), .B1(D12964_Y),     .Y(D12953_Y), .A0(D12993_Q));
KC_AOI22_X1 D12945 ( .A1(D11969_Y), .B0(D12984_Q), .B1(D11948_Y),     .Y(D12945_Y), .A0(D12983_Q));
KC_AOI22_X1 D12940 ( .A1(D11950_Y), .B0(D12982_Q), .B1(D11953_Y),     .Y(D12940_Y), .A0(D12980_Q));
KC_AOI22_X1 D12938 ( .A1(D11950_Y), .B0(D12978_Q), .B1(D11953_Y),     .Y(D12938_Y), .A0(D12979_Q));
KC_AOI22_X1 D12778 ( .A1(D12780_Y), .B0(D15474_Y), .B1(D12781_Y),     .Y(D12778_Y), .A0(D12804_Y));
KC_AOI22_X1 D12776 ( .A1(D12779_Y), .B0(D12788_Y), .B1(D12781_Y),     .Y(D12776_Y), .A0(D12804_Y));
KC_AOI22_X1 D12775 ( .A1(D12783_Y), .B0(D12787_Y), .B1(D12781_Y),     .Y(D12775_Y), .A0(D12804_Y));
KC_AOI22_X1 D12774 ( .A1(D12782_Y), .B0(D15491_Y), .B1(D12781_Y),     .Y(D12774_Y), .A0(D12804_Y));
KC_AOI22_X1 D12706 ( .A1(D13268_Q), .B0(D12739_Y), .B1(D12710_Y),     .Y(D12706_Y), .A0(D12298_Y));
KC_AOI22_X1 D12693 ( .A1(D12847_Y), .B0(D12254_Y), .B1(D12805_Y),     .Y(D12693_Y), .A0(D12712_Y));
KC_AOI22_X1 D12606 ( .A1(D11990_Y), .B0(D12610_Q), .B1(D12011_Y),     .Y(D12606_Y), .A0(D12607_Q));
KC_AOI22_X1 D12605 ( .A1(D13145_Q), .B0(D12010_Y), .B1(D1369_Q),     .Y(D12605_Y), .A0(D11438_Y));
KC_AOI22_X1 D12604 ( .A1(D1365_Q), .B0(D12010_Y), .B1(D1367_Q),     .Y(D12604_Y), .A0(D11438_Y));
KC_AOI22_X1 D12603 ( .A1(D11990_Y), .B0(D1367_Q), .B1(D12011_Y),     .Y(D12603_Y), .A0(D1365_Q));
KC_AOI22_X1 D12602 ( .A1(D12607_Q), .B0(D12010_Y), .B1(D12610_Q),     .Y(D12602_Y), .A0(D11438_Y));
KC_AOI22_X1 D12601 ( .A1(D12609_Q), .B0(D12010_Y), .B1(D12619_Q),     .Y(D12601_Y), .A0(D11438_Y));
KC_AOI22_X1 D12600 ( .A1(D11990_Y), .B0(D12619_Q), .B1(D12011_Y),     .Y(D12600_Y), .A0(D12609_Q));
KC_AOI22_X1 D12599 ( .A1(D12611_Q), .B0(D12010_Y), .B1(D12613_Q),     .Y(D12599_Y), .A0(D11438_Y));
KC_AOI22_X1 D12598 ( .A1(D11990_Y), .B0(D12613_Q), .B1(D12011_Y),     .Y(D12598_Y), .A0(D12611_Q));
KC_AOI22_X1 D12597 ( .A1(D12612_Q), .B0(D12010_Y), .B1(D12615_Q),     .Y(D12597_Y), .A0(D11438_Y));
KC_AOI22_X1 D12596 ( .A1(D11990_Y), .B0(D12615_Q), .B1(D12011_Y),     .Y(D12596_Y), .A0(D12612_Q));
KC_AOI22_X1 D12566 ( .A1(D12575_Q), .B0(D12012_Y), .B1(D12574_Q),     .Y(D12566_Y), .A0(D12052_Y));
KC_AOI22_X1 D12565 ( .A1(D12024_Y), .B0(D12579_Q), .B1(D12023_Y),     .Y(D12565_Y), .A0(D12583_Q));
KC_AOI22_X1 D12564 ( .A1(D12024_Y), .B0(D1311_Q), .B1(D12023_Y),     .Y(D12564_Y), .A0(D12577_Q));
KC_AOI22_X1 D12563 ( .A1(D13114_Q), .B0(D12012_Y), .B1(D13115_Q),     .Y(D12563_Y), .A0(D12052_Y));
KC_AOI22_X1 D12562 ( .A1(D12045_Q), .B0(D12025_Y), .B1(D2345_Q),     .Y(D12562_Y), .A0(D2301_Y));
KC_AOI22_X1 D12561 ( .A1(D12047_Y), .B0(D2345_Q), .B1(D12015_Y),     .Y(D12561_Y), .A0(D12045_Q));
KC_AOI22_X1 D12560 ( .A1(D12047_Y), .B0(D1310_Q), .B1(D12015_Y),     .Y(D12560_Y), .A0(D12581_Q));
KC_AOI22_X1 D12559 ( .A1(D12581_Q), .B0(D12025_Y), .B1(D1310_Q),     .Y(D12559_Y), .A0(D2301_Y));
KC_AOI22_X1 D12558 ( .A1(D2384_Q), .B0(D12025_Y), .B1(D1307_Q),     .Y(D12558_Y), .A0(D2301_Y));
KC_AOI22_X1 D12557 ( .A1(D12016_Y), .B0(D13115_Q), .B1(D12026_Y),     .Y(D12557_Y), .A0(D13114_Q));
KC_AOI22_X1 D12556 ( .A1(D12583_Q), .B0(D12051_Y), .B1(D12579_Q),     .Y(D12556_Y), .A0(D12050_Y));
KC_AOI22_X1 D12555 ( .A1(D12016_Y), .B0(D12574_Q), .B1(D12026_Y),     .Y(D12555_Y), .A0(D12575_Q));
KC_AOI22_X1 D12554 ( .A1(D12577_Q), .B0(D12051_Y), .B1(D1311_Q),     .Y(D12554_Y), .A0(D12050_Y));
KC_AOI22_X1 D12553 ( .A1(D12016_Y), .B0(D12576_Q), .B1(D12026_Y),     .Y(D12553_Y), .A0(D12584_Q));
KC_AOI22_X1 D12552 ( .A1(D12584_Q), .B0(D12012_Y), .B1(D12576_Q),     .Y(D12552_Y), .A0(D12052_Y));
KC_AOI22_X1 D12536 ( .A1(D12541_Q), .B0(D12012_Y), .B1(D1227_Q),     .Y(D12536_Y), .A0(D12052_Y));
KC_AOI22_X1 D12535 ( .A1(D12539_Q), .B0(D12012_Y), .B1(D12542_Q),     .Y(D12535_Y), .A0(D12052_Y));
KC_AOI22_X1 D12534 ( .A1(D12550_Q), .B0(D12012_Y), .B1(D12544_Q),     .Y(D12534_Y), .A0(D12052_Y));
KC_AOI22_X1 D12533 ( .A1(D12540_Q), .B0(D12051_Y), .B1(D2347_Q),     .Y(D12533_Y), .A0(D12050_Y));
KC_AOI22_X1 D12532 ( .A1(D12024_Y), .B0(D2347_Q), .B1(D12023_Y),     .Y(D12532_Y), .A0(D12540_Q));
KC_AOI22_X1 D12531 ( .A1(D12546_Q), .B0(D12051_Y), .B1(D2344_Q),     .Y(D12531_Y), .A0(D12050_Y));
KC_AOI22_X1 D12528 ( .A1(D12016_Y), .B0(D12543_Q), .B1(D12026_Y),     .Y(D12528_Y), .A0(D2348_Q));
KC_AOI22_X1 D12527 ( .A1(D12016_Y), .B0(D1227_Q), .B1(D12026_Y),     .Y(D12527_Y), .A0(D12541_Q));
KC_AOI22_X1 D12526 ( .A1(D12047_Y), .B0(D12507_Q), .B1(D12015_Y),     .Y(D12526_Y), .A0(D1142_Q));
KC_AOI22_X1 D12524 ( .A1(D2348_Q), .B0(D12012_Y), .B1(D12543_Q),     .Y(D12524_Y), .A0(D12052_Y));
KC_AOI22_X1 D12523 ( .A1(D12545_Q), .B0(D12051_Y), .B1(D1225_Q),     .Y(D12523_Y), .A0(D12050_Y));
KC_AOI22_X1 D12522 ( .A1(D12024_Y), .B0(D1225_Q), .B1(D12023_Y),     .Y(D12522_Y), .A0(D12545_Q));
KC_AOI22_X1 D12521 ( .A1(D12016_Y), .B0(D12542_Q), .B1(D12026_Y),     .Y(D12521_Y), .A0(D12539_Q));
KC_AOI22_X1 D12519 ( .A1(D1142_Q), .B0(D12025_Y), .B1(D12507_Q),     .Y(D12519_Y), .A0(D2301_Y));
KC_AOI22_X1 D12518 ( .A1(D12016_Y), .B0(D12544_Q), .B1(D12026_Y),     .Y(D12518_Y), .A0(D12550_Q));
KC_AOI22_X1 D12516 ( .A1(D12551_Q), .B0(D12051_Y), .B1(D2346_Q),     .Y(D12516_Y), .A0(D12050_Y));
KC_AOI22_X1 D12515 ( .A1(D12024_Y), .B0(D2346_Q), .B1(D12023_Y),     .Y(D12515_Y), .A0(D12551_Q));
KC_AOI22_X1 D12514 ( .A1(D12024_Y), .B0(D2344_Q), .B1(D12023_Y),     .Y(D12514_Y), .A0(D12546_Q));
KC_AOI22_X1 D12512 ( .A1(D2271_Y), .B0(D12496_Q), .B1(D2273_Y),     .Y(D12512_Y), .A0(D12506_Q));
KC_AOI22_X1 D12488 ( .A1(D12502_Q), .B0(D11929_Y), .B1(D1140_Q),     .Y(D12488_Y), .A0(D11930_Y));
KC_AOI22_X1 D12487 ( .A1(D11950_Y), .B0(D12458_Q), .B1(D11953_Y),     .Y(D12487_Y), .A0(D12452_Q));
KC_AOI22_X1 D12486 ( .A1(D11989_Y), .B0(D2349_Q), .B1(D11949_Y),     .Y(D12486_Y), .A0(D12505_Q));
KC_AOI22_X1 D12485 ( .A1(D12505_Q), .B0(D11951_Y), .B1(D2349_Q),     .Y(D12485_Y), .A0(D11981_Y));
KC_AOI22_X1 D12482 ( .A1(D11950_Y), .B0(D12454_Q), .B1(D11953_Y),     .Y(D12482_Y), .A0(D12455_Q));
KC_AOI22_X1 D12481 ( .A1(D2271_Y), .B0(D1136_Q), .B1(D2273_Y),     .Y(D12481_Y), .A0(D12497_Q));
KC_AOI22_X1 D12480 ( .A1(D12500_Q), .B0(D11951_Y), .B1(D12451_Q),     .Y(D12480_Y), .A0(D11981_Y));
KC_AOI22_X1 D12479 ( .A1(D11989_Y), .B0(D12451_Q), .B1(D11949_Y),     .Y(D12479_Y), .A0(D12500_Q));
KC_AOI22_X1 D12478 ( .A1(D12497_Q), .B0(D11929_Y), .B1(D1136_Q),     .Y(D12478_Y), .A0(D11930_Y));
KC_AOI22_X1 D12477 ( .A1(D2271_Y), .B0(D1140_Q), .B1(D2273_Y),     .Y(D12477_Y), .A0(D12502_Q));
KC_AOI22_X1 D12476 ( .A1(D12503_Q), .B0(D11929_Y), .B1(D12501_Q),     .Y(D12476_Y), .A0(D11930_Y));
KC_AOI22_X1 D12475 ( .A1(D12506_Q), .B0(D11929_Y), .B1(D12496_Q),     .Y(D12475_Y), .A0(D11930_Y));
KC_AOI22_X1 D12474 ( .A1(D2271_Y), .B0(D12501_Q), .B1(D2273_Y),     .Y(D12474_Y), .A0(D12503_Q));
KC_AOI22_X1 D12473 ( .A1(D11969_Y), .B0(D12495_Q), .B1(D11948_Y),     .Y(D12473_Y), .A0(D12494_Q));
KC_AOI22_X1 D12472 ( .A1(D12494_Q), .B0(D11991_Y), .B1(D12495_Q),     .Y(D12472_Y), .A0(D2277_Y));
KC_AOI22_X1 D12445 ( .A1(D11950_Y), .B0(D12461_Q), .B1(D11953_Y),     .Y(D12445_Y), .A0(D12462_Q));
KC_AOI22_X1 D12444 ( .A1(D11950_Y), .B0(D12466_Q), .B1(D11953_Y),     .Y(D12444_Y), .A0(D12465_Q));
KC_AOI22_X1 D12443 ( .A1(D12465_Q), .B0(D11952_Y), .B1(D12466_Q),     .Y(D12443_Y), .A0(D2272_Y));
KC_AOI22_X1 D12442 ( .A1(D12446_Y), .B0(D8340_Y), .B1(D12529_Y),     .Y(D12442_Y), .A0(D8348_Y));
KC_AOI22_X1 D12441 ( .A1(D12462_Q), .B0(D11952_Y), .B1(D12461_Q),     .Y(D12441_Y), .A0(D2272_Y));
KC_AOI22_X1 D12438 ( .A1(D11989_Y), .B0(D12463_Q), .B1(D11949_Y),     .Y(D12438_Y), .A0(D12464_Q));
KC_AOI22_X1 D12437 ( .A1(D12464_Q), .B0(D11951_Y), .B1(D12463_Q),     .Y(D12437_Y), .A0(D11981_Y));
KC_AOI22_X1 D12435 ( .A1(D12983_Q), .B0(D11991_Y), .B1(D12984_Q),     .Y(D12435_Y), .A0(D2277_Y));
KC_AOI22_X1 D12434 ( .A1(D2271_Y), .B0(D12459_Q), .B1(D2273_Y),     .Y(D12434_Y), .A0(D12460_Q));
KC_AOI22_X1 D12433 ( .A1(D12460_Q), .B0(D11929_Y), .B1(D12459_Q),     .Y(D12433_Y), .A0(D11930_Y));
KC_AOI22_X1 D12432 ( .A1(D12456_Q), .B0(D11951_Y), .B1(D12457_Q),     .Y(D12432_Y), .A0(D11981_Y));
KC_AOI22_X1 D12430 ( .A1(D11989_Y), .B0(D12457_Q), .B1(D11949_Y),     .Y(D12430_Y), .A0(D12456_Q));
KC_AOI22_X1 D12429 ( .A1(D12431_Y), .B0(D8340_Y), .B1(D13113_Y),     .Y(D12429_Y), .A0(D8348_Y));
KC_AOI22_X1 D12428 ( .A1(D12980_Q), .B0(D11952_Y), .B1(D12982_Q),     .Y(D12428_Y), .A0(D2272_Y));
KC_AOI22_X1 D12427 ( .A1(D12449_Q), .B0(D11951_Y), .B1(D12504_Q),     .Y(D12427_Y), .A0(D11981_Y));
KC_AOI22_X1 D12426 ( .A1(D11989_Y), .B0(D12504_Q), .B1(D11949_Y),     .Y(D12426_Y), .A0(D12449_Q));
KC_AOI22_X1 D12425 ( .A1(D12493_Y), .B0(D8340_Y), .B1(D13067_Y),     .Y(D12425_Y), .A0(D8348_Y));
KC_AOI22_X1 D12424 ( .A1(D12490_Y), .B0(D8340_Y), .B1(D13073_Y),     .Y(D12424_Y), .A0(D8348_Y));
KC_AOI22_X1 D12392 ( .A1(D12408_Q), .B0(D11952_Y), .B1(D12405_Q),     .Y(D12392_Y), .A0(D2272_Y));
KC_AOI22_X1 D12390 ( .A1(D12409_Q), .B0(D11929_Y), .B1(D12401_Q),     .Y(D12390_Y), .A0(D11930_Y));
KC_AOI22_X1 D12389 ( .A1(D11950_Y), .B0(D12404_Q), .B1(D11953_Y),     .Y(D12389_Y), .A0(D12403_Q));
KC_AOI22_X1 D12388 ( .A1(D12403_Q), .B0(D11952_Y), .B1(D12404_Q),     .Y(D12388_Y), .A0(D2272_Y));
KC_AOI22_X1 D12387 ( .A1(D12410_Q), .B0(D11951_Y), .B1(D12399_Q),     .Y(D12387_Y), .A0(D11981_Y));
KC_AOI22_X1 D12386 ( .A1(D12398_Q), .B0(D11951_Y), .B1(D12397_Q),     .Y(D12386_Y), .A0(D11981_Y));
KC_AOI22_X1 D12385 ( .A1(D11989_Y), .B0(D12406_Q), .B1(D11949_Y),     .Y(D12385_Y), .A0(D12407_Q));
KC_AOI22_X1 D12384 ( .A1(D2271_Y), .B0(D12401_Q), .B1(D2273_Y),     .Y(D12384_Y), .A0(D12409_Q));
KC_AOI22_X1 D12383 ( .A1(D11989_Y), .B0(D12397_Q), .B1(D11949_Y),     .Y(D12383_Y), .A0(D12398_Q));
KC_AOI22_X1 D12382 ( .A1(D11989_Y), .B0(D12399_Q), .B1(D11949_Y),     .Y(D12382_Y), .A0(D12410_Q));
KC_AOI22_X1 D12379 ( .A1(D12912_Q), .B0(D11991_Y), .B1(D12913_Q),     .Y(D12379_Y), .A0(D2277_Y));
KC_AOI22_X1 D12378 ( .A1(D12468_Q), .B0(D11929_Y), .B1(D12467_Q),     .Y(D12378_Y), .A0(D11930_Y));
KC_AOI22_X1 D12377 ( .A1(D2271_Y), .B0(D2352_Q), .B1(D2273_Y),     .Y(D12377_Y), .A0(D2351_Q));
KC_AOI22_X1 D12376 ( .A1(D11950_Y), .B0(D12405_Q), .B1(D11953_Y),     .Y(D12376_Y), .A0(D12408_Q));
KC_AOI22_X1 D12374 ( .A1(D12407_Q), .B0(D11951_Y), .B1(D12406_Q),     .Y(D12374_Y), .A0(D11981_Y));
KC_AOI22_X1 D12373 ( .A1(D12440_Y), .B0(D8340_Y), .B1(D12525_Y),     .Y(D12373_Y), .A0(D8348_Y));
KC_AOI22_X1 D12372 ( .A1(D12380_Y), .B0(D8340_Y), .B1(D12530_Y),     .Y(D12372_Y), .A0(D8348_Y));
KC_AOI22_X1 D12111 ( .A1(D12119_Q), .B0(D12117_Q), .B1(D12010_Y),     .Y(D12111_Y), .A0(D11438_Y));
KC_AOI22_X1 D12110 ( .A1(D12120_Q), .B0(D12010_Y), .B1(D12116_Q),     .Y(D12110_Y), .A0(D11438_Y));
KC_AOI22_X1 D12109 ( .A1(D11990_Y), .B0(D12122_Q), .B1(D12011_Y),     .Y(D12109_Y), .A0(D12121_Q));
KC_AOI22_X1 D12108 ( .A1(D12608_Q), .B0(D12010_Y), .B1(D12620_Q),     .Y(D12108_Y), .A0(D11438_Y));
KC_AOI22_X1 D12107 ( .A1(D11990_Y), .B0(D12116_Q), .B1(D12011_Y),     .Y(D12107_Y), .A0(D12120_Q));
KC_AOI22_X1 D12106 ( .A1(D11990_Y), .B0(D12117_Q), .B1(D12011_Y),     .Y(D12106_Y), .A0(D12119_Q));
KC_AOI22_X1 D12105 ( .A1(D11990_Y), .B0(D12620_Q), .B1(D12011_Y),     .Y(D12105_Y), .A0(D12608_Q));
KC_AOI22_X1 D12083 ( .A1(D12047_Y), .B0(D12087_Q), .B1(D12015_Y),     .Y(D12083_Y), .A0(D12093_Q));
KC_AOI22_X1 D12082 ( .A1(D12024_Y), .B0(D12090_Q), .B1(D12023_Y),     .Y(D12082_Y), .A0(D1316_Q));
KC_AOI22_X1 D12081 ( .A1(D12024_Y), .B0(D12096_Q), .B1(D12023_Y),     .Y(D12081_Y), .A0(D12095_Q));
KC_AOI22_X1 D12080 ( .A1(D12578_Q), .B0(D12051_Y), .B1(D12580_Q),     .Y(D12080_Y), .A0(D12050_Y));
KC_AOI22_X1 D12079 ( .A1(D12093_Q), .B0(D12025_Y), .B1(D12087_Q),     .Y(D12079_Y), .A0(D2301_Y));
KC_AOI22_X1 D12078 ( .A1(D12047_Y), .B0(D2289_Q), .B1(D12015_Y),     .Y(D12078_Y), .A0(D2291_Q));
KC_AOI22_X1 D12076 ( .A1(D2291_Q), .B0(D12025_Y), .B1(D2289_Q),     .Y(D12076_Y), .A0(D2301_Y));
KC_AOI22_X1 D12075 ( .A1(D12024_Y), .B0(D12580_Q), .B1(D12023_Y),     .Y(D12075_Y), .A0(D12578_Q));
KC_AOI22_X1 D12074 ( .A1(D11585_Q), .B0(D12025_Y), .B1(D12089_Q),     .Y(D12074_Y), .A0(D2301_Y));
KC_AOI22_X1 D12073 ( .A1(D12047_Y), .B0(D12089_Q), .B1(D12015_Y),     .Y(D12073_Y), .A0(D11585_Q));
KC_AOI22_X1 D12069 ( .A1(D1316_Q), .B0(D12051_Y), .B1(D12090_Q),     .Y(D12069_Y), .A0(D12050_Y));
KC_AOI22_X1 D12068 ( .A1(D12095_Q), .B0(D12051_Y), .B1(D12096_Q),     .Y(D12068_Y), .A0(D12050_Y));
KC_AOI22_X1 D12066 ( .A1(D12094_Q), .B0(D12012_Y), .B1(D12088_Q),     .Y(D12066_Y), .A0(D12052_Y));
KC_AOI22_X1 D12065 ( .A1(D12016_Y), .B0(D1317_Q), .B1(D12026_Y),     .Y(D12065_Y), .A0(D11584_Q));
KC_AOI22_X1 D12064 ( .A1(D12016_Y), .B0(D12088_Q), .B1(D12026_Y),     .Y(D12064_Y), .A0(D12094_Q));
KC_AOI22_X1 D12063 ( .A1(D12582_Q), .B0(D12012_Y), .B1(D12585_Q),     .Y(D12063_Y), .A0(D12052_Y));
KC_AOI22_X1 D12062 ( .A1(D12016_Y), .B0(D12585_Q), .B1(D12026_Y),     .Y(D12062_Y), .A0(D12582_Q));
KC_AOI22_X1 D12060 ( .A1(D12121_Q), .B0(D12010_Y), .B1(D12122_Q),     .Y(D12060_Y), .A0(D11438_Y));
KC_AOI22_X1 D12021 ( .A1(D2292_Q), .B0(D12025_Y), .B1(D12044_Q),     .Y(D12021_Y), .A0(D2301_Y));
KC_AOI22_X1 D12020 ( .A1(D12047_Y), .B0(D2290_Q), .B1(D12015_Y),     .Y(D12020_Y), .A0(D129_Q));
KC_AOI22_X1 D12019 ( .A1(D12052_Y), .B0(D12092_Q), .B1(D12012_Y),     .Y(D12019_Y), .A0(D2248_Q));
KC_AOI22_X1 D12014 ( .A1(D12047_Y), .B0(D1247_Q), .B1(D12015_Y),     .Y(D12014_Y), .A0(D12058_Q));
KC_AOI22_X1 D12009 ( .A1(D12058_Q), .B0(D12025_Y), .B1(D1247_Q),     .Y(D12009_Y), .A0(D2301_Y));
KC_AOI22_X1 D12008 ( .A1(D12047_Y), .B0(D12044_Q), .B1(D12015_Y),     .Y(D12008_Y), .A0(D2292_Q));
KC_AOI22_X1 D12007 ( .A1(D132_Q), .B0(D12025_Y), .B1(D1222_Q),     .Y(D12007_Y), .A0(D2301_Y));
KC_AOI22_X1 D12002 ( .A1(D12050_Y), .B0(D12046_Q), .B1(D12051_Y),     .Y(D12002_Y), .A0(D1312_Q));
KC_AOI22_X1 D12001 ( .A1(D12024_Y), .B0(D12046_Q), .B1(D12023_Y),     .Y(D12001_Y), .A0(D1312_Q));
KC_AOI22_X1 D11998 ( .A1(D2301_Y), .B0(D2290_Q), .B1(D12025_Y),     .Y(D11998_Y), .A0(D129_Q));
KC_AOI22_X1 D11997 ( .A1(D12016_Y), .B0(D12092_Q), .B1(D12026_Y),     .Y(D11997_Y), .A0(D2248_Q));
KC_AOI22_X1 D11944 ( .A1(D2271_Y), .B0(D1138_Q), .B1(D2273_Y),     .Y(D11944_Y), .A0(D1139_Q));
KC_AOI22_X1 D11943 ( .A1(D1139_Q), .B0(D11929_Y), .B1(D1138_Q),     .Y(D11943_Y), .A0(D11930_Y));
KC_AOI22_X1 D11939 ( .A1(D11975_Q), .B0(D11991_Y), .B1(D11971_Q),     .Y(D11939_Y), .A0(D2277_Y));
KC_AOI22_X1 D11938 ( .A1(D11969_Y), .B0(D11971_Q), .B1(D11948_Y),     .Y(D11938_Y), .A0(D11975_Q));
KC_AOI22_X1 D11937 ( .A1(D11972_Q), .B0(D11991_Y), .B1(D11973_Q),     .Y(D11937_Y), .A0(D2277_Y));
KC_AOI22_X1 D11936 ( .A1(D11969_Y), .B0(D11973_Q), .B1(D11948_Y),     .Y(D11936_Y), .A0(D11972_Q));
KC_AOI22_X1 D11935 ( .A1(D11969_Y), .B0(D1134_Q), .B1(D11948_Y),     .Y(D11935_Y), .A0(D1135_Q));
KC_AOI22_X1 D11934 ( .A1(D1135_Q), .B0(D11991_Y), .B1(D1134_Q),     .Y(D11934_Y), .A0(D2277_Y));
KC_AOI22_X1 D11902 ( .A1(D2294_Q), .B0(D11991_Y), .B1(D11864_Q),     .Y(D11902_Y), .A0(D2277_Y));
KC_AOI22_X1 D11901 ( .A1(D11969_Y), .B0(D11926_Q), .B1(D11948_Y),     .Y(D11901_Y), .A0(D11863_Q));
KC_AOI22_X1 D11899 ( .A1(D11950_Y), .B0(D1041_Q), .B1(D11953_Y),     .Y(D11899_Y), .A0(D1038_Q));
KC_AOI22_X1 D11898 ( .A1(D1038_Q), .B0(D11952_Y), .B1(D1041_Q),     .Y(D11898_Y), .A0(D2272_Y));
KC_AOI22_X1 D11897 ( .A1(D11989_Y), .B0(D11925_Q), .B1(D11949_Y),     .Y(D11897_Y), .A0(D11924_Q));
KC_AOI22_X1 D11896 ( .A1(D11924_Q), .B0(D11951_Y), .B1(D11925_Q),     .Y(D11896_Y), .A0(D11981_Y));
KC_AOI22_X1 D11895 ( .A1(D1034_Q), .B0(D11929_Y), .B1(D1035_Q),     .Y(D11895_Y), .A0(D11930_Y));
KC_AOI22_X1 D11894 ( .A1(D2271_Y), .B0(D1035_Q), .B1(D2273_Y),     .Y(D11894_Y), .A0(D1034_Q));
KC_AOI22_X1 D11892 ( .A1(D11918_Q), .B0(D11951_Y), .B1(D11920_Q),     .Y(D11892_Y), .A0(D11981_Y));
KC_AOI22_X1 D11891 ( .A1(D11917_Q), .B0(D11951_Y), .B1(D11919_Q),     .Y(D11891_Y), .A0(D11981_Y));
KC_AOI22_X1 D11890 ( .A1(D11989_Y), .B0(D11919_Q), .B1(D11949_Y),     .Y(D11890_Y), .A0(D11917_Q));
KC_AOI22_X1 D11889 ( .A1(D11989_Y), .B0(D11920_Q), .B1(D11949_Y),     .Y(D11889_Y), .A0(D11918_Q));
KC_AOI22_X1 D11886 ( .A1(D11950_Y), .B0(D1030_Q), .B1(D11953_Y),     .Y(D11886_Y), .A0(D11923_Q));
KC_AOI22_X1 D11885 ( .A1(D2271_Y), .B0(D11979_Q), .B1(D2273_Y),     .Y(D11885_Y), .A0(D11977_Q));
KC_AOI22_X1 D11884 ( .A1(D11922_Q), .B0(D11952_Y), .B1(D11921_Q),     .Y(D11884_Y), .A0(D2272_Y));
KC_AOI22_X1 D11883 ( .A1(D11923_Q), .B0(D11952_Y), .B1(D1030_Q),     .Y(D11883_Y), .A0(D2272_Y));
KC_AOI22_X1 D11882 ( .A1(D1026_Q), .B0(D11951_Y), .B1(D1027_Q),     .Y(D11882_Y), .A0(D11981_Y));
KC_AOI22_X1 D11881 ( .A1(D11989_Y), .B0(D1027_Q), .B1(D11949_Y),     .Y(D11881_Y), .A0(D1026_Q));
KC_AOI22_X1 D11880 ( .A1(D11950_Y), .B0(D11921_Q), .B1(D11953_Y),     .Y(D11880_Y), .A0(D11922_Q));
KC_AOI22_X1 D11879 ( .A1(D11977_Q), .B0(D11929_Y), .B1(D11979_Q),     .Y(D11879_Y), .A0(D11930_Y));
KC_AOI22_X1 D11841 ( .A1(D11860_Q), .B0(D11951_Y), .B1(D11870_Q),     .Y(D11841_Y), .A0(D11981_Y));
KC_AOI22_X1 D11840 ( .A1(D11981_Y), .B0(D11869_Q), .B1(D11951_Y),     .Y(D11840_Y), .A0(D11857_Q));
KC_AOI22_X1 D11839 ( .A1(D910_Q), .B0(D11951_Y), .B1(D12402_Q),     .Y(D11839_Y), .A0(D11981_Y));
KC_AOI22_X1 D11838 ( .A1(D11989_Y), .B0(D12402_Q), .B1(D11949_Y),     .Y(D11838_Y), .A0(D910_Q));
KC_AOI22_X1 D11836 ( .A1(D11989_Y), .B0(D11869_Q), .B1(D11949_Y),     .Y(D11836_Y), .A0(D11857_Q));
KC_AOI22_X1 D11835 ( .A1(D11989_Y), .B0(D11870_Q), .B1(D11949_Y),     .Y(D11835_Y), .A0(D11860_Q));
KC_AOI22_X1 D11833 ( .A1(D11856_Q), .B0(D11952_Y), .B1(D11868_Q),     .Y(D11833_Y), .A0(D2272_Y));
KC_AOI22_X1 D11832 ( .A1(D12569_Y), .B0(D8337_Y), .B1(D11760_Y),     .Y(D11832_Y), .A0(D8340_Y));
KC_AOI22_X1 D11831 ( .A1(D11862_Q), .B0(D11929_Y), .B1(D11858_Q),     .Y(D11831_Y), .A0(D11930_Y));
KC_AOI22_X1 D11830 ( .A1(D909_Q), .B0(D11952_Y), .B1(D919_Q),     .Y(D11830_Y), .A0(D2272_Y));
KC_AOI22_X1 D11829 ( .A1(D2272_Y), .B0(D11855_Q), .B1(D11952_Y),     .Y(D11829_Y), .A0(D11867_Q));
KC_AOI22_X1 D11828 ( .A1(D920_Q), .B0(D11929_Y), .B1(D12400_Q),     .Y(D11828_Y), .A0(D11930_Y));
KC_AOI22_X1 D11825 ( .A1(D2271_Y), .B0(D11871_Q), .B1(D2273_Y),     .Y(D11825_Y), .A0(D11861_Q));
KC_AOI22_X1 D11824 ( .A1(D11930_Y), .B0(D11871_Q), .B1(D11929_Y),     .Y(D11824_Y), .A0(D11861_Q));
KC_AOI22_X1 D11823 ( .A1(D11950_Y), .B0(D11855_Q), .B1(D11953_Y),     .Y(D11823_Y), .A0(D11867_Q));
KC_AOI22_X1 D11822 ( .A1(D2271_Y), .B0(D11858_Q), .B1(D2273_Y),     .Y(D11822_Y), .A0(D11862_Q));
KC_AOI22_X1 D11821 ( .A1(D11950_Y), .B0(D919_Q), .B1(D11953_Y),     .Y(D11821_Y), .A0(D909_Q));
KC_AOI22_X1 D11820 ( .A1(D11950_Y), .B0(D11868_Q), .B1(D11953_Y),     .Y(D11820_Y), .A0(D11856_Q));
KC_AOI22_X1 D11819 ( .A1(D2271_Y), .B0(D12400_Q), .B1(D2273_Y),     .Y(D11819_Y), .A0(D920_Q));
KC_AOI22_X1 D11818 ( .A1(D12067_Y), .B0(D8337_Y), .B1(D11771_Y),     .Y(D11818_Y), .A0(D8340_Y));
KC_AOI22_X1 D11817 ( .A1(D12003_Y), .B0(D8337_Y), .B1(D11761_Y),     .Y(D11817_Y), .A0(D8340_Y));
KC_AOI22_X1 D11816 ( .A1(D12077_Y), .B0(D8337_Y), .B1(D11744_Y),     .Y(D11816_Y), .A0(D8340_Y));
KC_AOI22_X1 D11814 ( .A1(D11969_Y), .B0(D11864_Q), .B1(D11948_Y),     .Y(D11814_Y), .A0(D2294_Q));
KC_AOI22_X1 D11813 ( .A1(D11969_Y), .B0(D2350_Q), .B1(D11948_Y),     .Y(D11813_Y), .A0(D2293_Q));
KC_AOI22_X1 D11812 ( .A1(D11969_Y), .B0(D915_Q), .B1(D11948_Y),     .Y(D11812_Y), .A0(D134_Q));
KC_AOI22_X1 D11811 ( .A1(D134_Q), .B0(D11991_Y), .B1(D915_Q),     .Y(D11811_Y), .A0(D2277_Y));
KC_AOI22_X1 D11774 ( .A1(D11802_Q), .B0(D10818_Y), .B1(D810_Q),     .Y(D11774_Y), .A0(D10765_Y));
KC_AOI22_X1 D11773 ( .A1(D10672_Y), .B0(D11719_Q), .B1(D10757_Y),     .Y(D11773_Y), .A0(D11804_Q));
KC_AOI22_X1 D11772 ( .A1(D10766_Y), .B0(D810_Q), .B1(D10727_Y),     .Y(D11772_Y), .A0(D11802_Q));
KC_AOI22_X1 D11769 ( .A1(D10804_Y), .B0(D11799_Q), .B1(D10663_Y),     .Y(D11769_Y), .A0(D11796_Q));
KC_AOI22_X1 D11768 ( .A1(D11796_Q), .B0(D10743_Y), .B1(D11799_Q),     .Y(D11768_Y), .A0(D10805_Y));
KC_AOI22_X1 D11766 ( .A1(D804_Q), .B0(D10818_Y), .B1(D807_Q),     .Y(D11766_Y), .A0(D10765_Y));
KC_AOI22_X1 D11765 ( .A1(D11798_Q), .B0(D10808_Y), .B1(D11801_Q),     .Y(D11765_Y), .A0(D10809_Y));
KC_AOI22_X1 D11764 ( .A1(D10766_Y), .B0(D807_Q), .B1(D10727_Y),     .Y(D11764_Y), .A0(D804_Q));
KC_AOI22_X1 D11763 ( .A1(D10749_Y), .B0(D11801_Q), .B1(D10750_Y),     .Y(D11763_Y), .A0(D11798_Q));
KC_AOI22_X1 D11759 ( .A1(D10672_Y), .B0(D802_Q), .B1(D10757_Y),     .Y(D11759_Y), .A0(D800_Q));
KC_AOI22_X1 D11758 ( .A1(D10749_Y), .B0(D798_Q), .B1(D10750_Y),     .Y(D11758_Y), .A0(D11793_Q));
KC_AOI22_X1 D11757 ( .A1(D11795_Q), .B0(D10742_Y), .B1(D799_Q),     .Y(D11757_Y), .A0(D10745_Y));
KC_AOI22_X1 D11756 ( .A1(D10672_Y), .B0(D799_Q), .B1(D10757_Y),     .Y(D11756_Y), .A0(D11795_Q));
KC_AOI22_X1 D11755 ( .A1(D10745_Y), .B0(D802_Q), .B1(D10742_Y),     .Y(D11755_Y), .A0(D800_Q));
KC_AOI22_X1 D11752 ( .A1(D11790_Q), .B0(D10743_Y), .B1(D2297_Q),     .Y(D11752_Y), .A0(D10805_Y));
KC_AOI22_X1 D11751 ( .A1(D10804_Y), .B0(D11788_Q), .B1(D10663_Y),     .Y(D11751_Y), .A0(D2296_Q));
KC_AOI22_X1 D11750 ( .A1(D11793_Q), .B0(D10808_Y), .B1(D798_Q),     .Y(D11750_Y), .A0(D10809_Y));
KC_AOI22_X1 D11749 ( .A1(D12337_Q), .B0(D10742_Y), .B1(D12336_Q),     .Y(D11749_Y), .A0(D10745_Y));
KC_AOI22_X1 D11748 ( .A1(D10749_Y), .B0(D11792_Q), .B1(D10750_Y),     .Y(D11748_Y), .A0(D11789_Q));
KC_AOI22_X1 D11747 ( .A1(D11791_Q), .B0(D10743_Y), .B1(D11794_Q),     .Y(D11747_Y), .A0(D10805_Y));
KC_AOI22_X1 D11746 ( .A1(D10805_Y), .B0(D11788_Q), .B1(D10743_Y),     .Y(D11746_Y), .A0(D2296_Q));
KC_AOI22_X1 D11745 ( .A1(D10804_Y), .B0(D11794_Q), .B1(D10663_Y),     .Y(D11745_Y), .A0(D11791_Q));
KC_AOI22_X1 D11743 ( .A1(D10672_Y), .B0(D12336_Q), .B1(D10757_Y),     .Y(D11743_Y), .A0(D12337_Q));
KC_AOI22_X1 D11742 ( .A1(D10804_Y), .B0(D2297_Q), .B1(D10663_Y),     .Y(D11742_Y), .A0(D11790_Q));
KC_AOI22_X1 D11741 ( .A1(D2295_Q), .B0(D10808_Y), .B1(D137_Q),     .Y(D11741_Y), .A0(D10809_Y));
KC_AOI22_X1 D11740 ( .A1(D10809_Y), .B0(D11792_Q), .B1(D10808_Y),     .Y(D11740_Y), .A0(D11789_Q));
KC_AOI22_X1 D11739 ( .A1(D10749_Y), .B0(D137_Q), .B1(D10750_Y),     .Y(D11739_Y), .A0(D2295_Q));
KC_AOI22_X1 D11736 ( .A1(D11683_Y), .B0(D136_Q), .B1(D11776_Y),     .Y(D11736_Y), .A0(D11255_Y));
KC_AOI22_X1 D11708 ( .A1(D10749_Y), .B0(D11723_Q), .B1(D10750_Y),     .Y(D11708_Y), .A0(D11724_Q));
KC_AOI22_X1 D11707 ( .A1(D10672_Y), .B0(D687_Q), .B1(D10757_Y),     .Y(D11707_Y), .A0(D11722_Q));
KC_AOI22_X1 D11706 ( .A1(D11725_Q), .B0(D10818_Y), .B1(D2288_Q),     .Y(D11706_Y), .A0(D10765_Y));
KC_AOI22_X1 D11705 ( .A1(D11722_Q), .B0(D10742_Y), .B1(D687_Q),     .Y(D11705_Y), .A0(D10745_Y));
KC_AOI22_X1 D11703 ( .A1(D11726_Q), .B0(D10808_Y), .B1(D690_Q),     .Y(D11703_Y), .A0(D10809_Y));
KC_AOI22_X1 D11702 ( .A1(D10749_Y), .B0(D690_Q), .B1(D10750_Y),     .Y(D11702_Y), .A0(D11726_Q));
KC_AOI22_X1 D11701 ( .A1(D10672_Y), .B0(D12306_Q), .B1(D10757_Y),     .Y(D11701_Y), .A0(D728_Q));
KC_AOI22_X1 D11698 ( .A1(D11724_Q), .B0(D10808_Y), .B1(D11723_Q),     .Y(D11698_Y), .A0(D10809_Y));
KC_AOI22_X1 D11696 ( .A1(D11735_Q), .B0(D10743_Y), .B1(D11734_Q),     .Y(D11696_Y), .A0(D10805_Y));
KC_AOI22_X1 D11695 ( .A1(D728_Q), .B0(D10742_Y), .B1(D12306_Q),     .Y(D11695_Y), .A0(D10745_Y));
KC_AOI22_X1 D11694 ( .A1(D10766_Y), .B0(D729_Q), .B1(D10727_Y),     .Y(D11694_Y), .A0(D11731_Q));
KC_AOI22_X1 D11693 ( .A1(D11731_Q), .B0(D10818_Y), .B1(D729_Q),     .Y(D11693_Y), .A0(D10765_Y));
KC_AOI22_X1 D11692 ( .A1(D10804_Y), .B0(D11734_Q), .B1(D10663_Y),     .Y(D11692_Y), .A0(D11735_Q));
KC_AOI22_X1 D11691 ( .A1(D11720_Q), .B0(D10743_Y), .B1(D11733_Q),     .Y(D11691_Y), .A0(D10805_Y));
KC_AOI22_X1 D11690 ( .A1(D10766_Y), .B0(D681_Q), .B1(D10727_Y),     .Y(D11690_Y), .A0(D678_Q));
KC_AOI22_X1 D11689 ( .A1(D10804_Y), .B0(D11733_Q), .B1(D10663_Y),     .Y(D11689_Y), .A0(D11720_Q));
KC_AOI22_X1 D11688 ( .A1(D11732_Q), .B0(D10742_Y), .B1(D12270_Q),     .Y(D11688_Y), .A0(D10745_Y));
KC_AOI22_X1 D11687 ( .A1(D10672_Y), .B0(D12270_Q), .B1(D10757_Y),     .Y(D11687_Y), .A0(D11732_Q));
KC_AOI22_X1 D11686 ( .A1(D11804_Q), .B0(D10742_Y), .B1(D11719_Q),     .Y(D11686_Y), .A0(D10745_Y));
KC_AOI22_X1 D11685 ( .A1(D11715_Q), .B0(D10808_Y), .B1(D684_Q),     .Y(D11685_Y), .A0(D10809_Y));
KC_AOI22_X1 D11684 ( .A1(D10749_Y), .B0(D684_Q), .B1(D10750_Y),     .Y(D11684_Y), .A0(D11715_Q));
KC_AOI22_X1 D11681 ( .A1(D10804_Y), .B0(D11718_Q), .B1(D10663_Y),     .Y(D11681_Y), .A0(D11803_Q));
KC_AOI22_X1 D11680 ( .A1(D11803_Q), .B0(D10743_Y), .B1(D11718_Q),     .Y(D11680_Y), .A0(D10805_Y));
KC_AOI22_X1 D11679 ( .A1(D678_Q), .B0(D10818_Y), .B1(D681_Q),     .Y(D11679_Y), .A0(D10765_Y));
KC_AOI22_X1 D11665 ( .A1(D11650_Y), .B0(D11671_Y), .B1(D11663_Y),     .Y(D11665_Y), .A0(D11663_Y));
KC_AOI22_X1 D11647 ( .A1(D10766_Y), .B0(D11662_Q), .B1(D10727_Y),     .Y(D11647_Y), .A0(D11659_Q));
KC_AOI22_X1 D11644 ( .A1(D10766_Y), .B0(D11656_Q), .B1(D10727_Y),     .Y(D11644_Y), .A0(D11661_Q));
KC_AOI22_X1 D11643 ( .A1(D11659_Q), .B0(D11662_Q), .B1(D10818_Y),     .Y(D11643_Y), .A0(D10765_Y));
KC_AOI22_X1 D11501 ( .A1(D12537_Y), .B0(D2249_Q), .B1(D11522_Y),     .Y(D11501_Y), .A0(D9725_Y));
KC_AOI22_X1 D11500 ( .A1(D12022_Y), .B0(D2251_Q), .B1(D11523_Y),     .Y(D11500_Y), .A0(D9725_Y));
KC_AOI22_X1 D11498 ( .A1(D12568_Y), .B0(D11543_Q), .B1(D11525_Y),     .Y(D11498_Y), .A0(D9725_Y));
KC_AOI22_X1 D11497 ( .A1(D12517_Y), .B0(D11537_Q), .B1(D11520_Y),     .Y(D11497_Y), .A0(D9725_Y));
KC_AOI22_X1 D11496 ( .A1(D12061_Y), .B0(D11539_Q), .B1(D11518_Y),     .Y(D11496_Y), .A0(D9725_Y));
KC_AOI22_X1 D11495 ( .A1(D12538_Y), .B0(D1219_Q), .B1(D11517_Y),     .Y(D11495_Y), .A0(D9725_Y));
KC_AOI22_X1 D11489 ( .A1(D1264_Y), .B0(D11538_Q), .B1(D11521_Y),     .Y(D11489_Y), .A0(D2032_Y));
KC_AOI22_X1 D11485 ( .A1(D12071_Y), .B0(D11542_Q), .B1(D11519_Y),     .Y(D11485_Y), .A0(D2032_Y));
KC_AOI22_X1 D11482 ( .A1(D13074_Y), .B0(D131_Q), .B1(D11514_Y),     .Y(D11482_Y), .A0(D2032_Y));
KC_AOI22_X1 D11480 ( .A1(D13057_Y), .B0(D1224_Q), .B1(D11516_Y),     .Y(D11480_Y), .A0(D9725_Y));
KC_AOI22_X1 D11434 ( .A1(D12489_Y), .B0(D2253_Q), .B1(D2234_Y),     .Y(D11434_Y), .A0(D11255_Y));
KC_AOI22_X1 D11433 ( .A1(D11947_Y), .B0(D11468_Q), .B1(D11441_Y),     .Y(D11433_Y), .A0(D8211_Y));
KC_AOI22_X1 D11429 ( .A1(D11440_Y), .B0(D11255_Y), .B1(D2269_Y),     .Y(D11429_Y), .A0(D11475_Q));
KC_AOI22_X1 D11427 ( .A1(D2184_Y), .B0(D11467_Q), .B1(D10903_Y),     .Y(D11427_Y), .A0(D11471_Q));
KC_AOI22_X1 D11423 ( .A1(D12484_Y), .B0(D11466_Q), .B1(D11442_Y),     .Y(D11423_Y), .A0(D11255_Y));
KC_AOI22_X1 D11422 ( .A1(D12436_Y), .B0(D11469_Q), .B1(D11439_Y),     .Y(D11422_Y), .A0(D11255_Y));
KC_AOI22_X1 D11371 ( .A1(D2254_Q), .B0(D2190_Y), .B1(D11401_Q),     .Y(D11371_Y), .A0(D2242_Y));
KC_AOI22_X1 D11370 ( .A1(D10990_Y), .B0(D11401_Q), .B1(D10912_Y),     .Y(D11370_Y), .A0(D2254_Q));
KC_AOI22_X1 D11368 ( .A1(D10990_Y), .B0(D11399_Q), .B1(D10912_Y),     .Y(D11368_Y), .A0(D11398_Q));
KC_AOI22_X1 D11367 ( .A1(D10990_Y), .B0(D11400_Q), .B1(D10912_Y),     .Y(D11367_Y), .A0(D1040_Q));
KC_AOI22_X1 D11362 ( .A1(D11398_Q), .B0(D2190_Y), .B1(D11399_Q),     .Y(D11362_Y), .A0(D2242_Y));
KC_AOI22_X1 D11361 ( .A1(D10990_Y), .B0(D11397_Q), .B1(D10912_Y),     .Y(D11361_Y), .A0(D11395_Q));
KC_AOI22_X1 D11360 ( .A1(D11394_Q), .B0(D11396_Q), .B1(D2190_Y),     .Y(D11360_Y), .A0(D2242_Y));
KC_AOI22_X1 D11359 ( .A1(D11395_Q), .B0(D2190_Y), .B1(D11397_Q),     .Y(D11359_Y), .A0(D2242_Y));
KC_AOI22_X1 D11356 ( .A1(D12491_Y), .B0(D11340_Q), .B1(D11378_Y),     .Y(D11356_Y), .A0(D11255_Y));
KC_AOI22_X1 D11355 ( .A1(D10990_Y), .B0(D11396_Q), .B1(D10912_Y),     .Y(D11355_Y), .A0(D11394_Q));
KC_AOI22_X1 D11351 ( .A1(D12492_Y), .B0(D11392_Q), .B1(D11376_Y),     .Y(D11351_Y), .A0(D11255_Y));
KC_AOI22_X1 D11301 ( .A1(D2276_Y), .B0(D11327_Q), .B1(D11307_Y),     .Y(D11301_Y), .A0(D11255_Y));
KC_AOI22_X1 D11298 ( .A1(D11837_Y), .B0(D11342_Q), .B1(D11311_Y),     .Y(D11298_Y), .A0(D11255_Y));
KC_AOI22_X1 D11291 ( .A1(D11878_Y), .B0(D11341_Q), .B1(D11306_Y),     .Y(D11291_Y), .A0(D11255_Y));
KC_AOI22_X1 D11290 ( .A1(D11309_Y), .B0(D11255_Y), .B1(D12375_Y),     .Y(D11290_Y), .A0(D11325_Q));
KC_AOI22_X1 D11289 ( .A1(D12423_Y), .B0(D11329_Q), .B1(D11304_Y),     .Y(D11289_Y), .A0(D11255_Y));
KC_AOI22_X1 D11284 ( .A1(D12439_Y), .B0(D11326_Q), .B1(D11312_Y),     .Y(D11284_Y), .A0(D11255_Y));
KC_AOI22_X1 D11283 ( .A1(D10990_Y), .B0(D11338_Q), .B1(D10912_Y),     .Y(D11283_Y), .A0(D11339_Q));
KC_AOI22_X1 D11282 ( .A1(D11339_Q), .B0(D2190_Y), .B1(D11338_Q),     .Y(D11282_Y), .A0(D2242_Y));
KC_AOI22_X1 D11281 ( .A1(D11335_Q), .B0(D2190_Y), .B1(D11337_Q),     .Y(D11281_Y), .A0(D2242_Y));
KC_AOI22_X1 D11280 ( .A1(D10990_Y), .B0(D11337_Q), .B1(D10912_Y),     .Y(D11280_Y), .A0(D11335_Q));
KC_AOI22_X1 D11227 ( .A1(D10766_Y), .B0(D11717_Q), .B1(D10727_Y),     .Y(D11227_Y), .A0(D11175_Q));
KC_AOI22_X1 D11226 ( .A1(D11266_Q), .B0(D10743_Y), .B1(D11274_Q),     .Y(D11226_Y), .A0(D10805_Y));
KC_AOI22_X1 D11225 ( .A1(D10672_Y), .B0(D677_Q), .B1(D10757_Y),     .Y(D11225_Y), .A0(D803_Q));
KC_AOI22_X1 D11224 ( .A1(D11267_Q), .B0(D10743_Y), .B1(D11275_Q),     .Y(D11224_Y), .A0(D10805_Y));
KC_AOI22_X1 D11223 ( .A1(D10804_Y), .B0(D11275_Q), .B1(D10663_Y),     .Y(D11223_Y), .A0(D11267_Q));
KC_AOI22_X1 D11221 ( .A1(D10749_Y), .B0(D11273_Q), .B1(D10750_Y),     .Y(D11221_Y), .A0(D11269_Q));
KC_AOI22_X1 D11220 ( .A1(D10804_Y), .B0(D806_Q), .B1(D10663_Y),     .Y(D11220_Y), .A0(D683_Q));
KC_AOI22_X1 D11219 ( .A1(D10749_Y), .B0(D11272_Q), .B1(D10750_Y),     .Y(D11219_Y), .A0(D11270_Q));
KC_AOI22_X1 D11216 ( .A1(D10749_Y), .B0(D809_Q), .B1(D10750_Y),     .Y(D11216_Y), .A0(D11268_Q));
KC_AOI22_X1 D11215 ( .A1(D11269_Q), .B0(D10808_Y), .B1(D11273_Q),     .Y(D11215_Y), .A0(D10809_Y));
KC_AOI22_X1 D11213 ( .A1(D11270_Q), .B0(D10808_Y), .B1(D11272_Q),     .Y(D11213_Y), .A0(D10809_Y));
KC_AOI22_X1 D11211 ( .A1(D11268_Q), .B0(D10808_Y), .B1(D809_Q),     .Y(D11211_Y), .A0(D10809_Y));
KC_AOI22_X1 D11208 ( .A1(D11699_Y), .B0(D11265_Q), .B1(D11237_Y),     .Y(D11208_Y), .A0(D11255_Y));
KC_AOI22_X1 D11207 ( .A1(D11697_Y), .B0(D11261_Q), .B1(D11239_Y),     .Y(D11207_Y), .A0(D11255_Y));
KC_AOI22_X1 D11206 ( .A1(D11222_Y), .B0(D11262_Q), .B1(D11238_Y),     .Y(D11206_Y), .A0(D8211_Y));
KC_AOI22_X1 D11203 ( .A1(D10675_Y), .B0(D11264_Q), .B1(D11234_Y),     .Y(D11203_Y), .A0(D8211_Y));
KC_AOI22_X1 D11198 ( .A1(D10754_Y), .B0(D11263_Q), .B1(D11235_Y),     .Y(D11198_Y), .A0(D8211_Y));
KC_AOI22_X1 D11195 ( .A1(D11218_Y), .B0(D2256_Q), .B1(D766_Y),     .Y(D11195_Y), .A0(D11255_Y));
KC_AOI22_X1 D11189 ( .A1(D11255_Y), .B0(D10790_Q), .B1(D11231_Y),     .Y(D11189_Y), .A0(D11762_Y));
KC_AOI22_X1 D11141 ( .A1(D11175_Q), .B0(D10818_Y), .B1(D11717_Q),     .Y(D11141_Y), .A0(D10765_Y));
KC_AOI22_X1 D11138 ( .A1(D10804_Y), .B0(D11274_Q), .B1(D10663_Y),     .Y(D11138_Y), .A0(D11266_Q));
KC_AOI22_X1 D11137 ( .A1(D10672_Y), .B0(D11178_Q), .B1(D10757_Y),     .Y(D11137_Y), .A0(D11176_Q));
KC_AOI22_X1 D11136 ( .A1(D11176_Q), .B0(D10742_Y), .B1(D11178_Q),     .Y(D11136_Y), .A0(D10745_Y));
KC_AOI22_X1 D11121 ( .A1(D10766_Y), .B0(D2247_Q), .B1(D10727_Y),     .Y(D11121_Y), .A0(D2245_Q));
KC_AOI22_X1 D11120 ( .A1(D2245_Q), .B0(D10818_Y), .B1(D2247_Q),     .Y(D11120_Y), .A0(D10765_Y));
KC_AOI22_X1 D11119 ( .A1(D10766_Y), .B0(D11125_Q), .B1(D10727_Y),     .Y(D11119_Y), .A0(D11126_Q));
KC_AOI22_X1 D11118 ( .A1(D11126_Q), .B0(D10818_Y), .B1(D11125_Q),     .Y(D11118_Y), .A0(D10765_Y));
KC_AOI22_X1 D11097 ( .A1(D9555_Y), .B0(D11110_Q), .B1(D10541_Y),     .Y(D11097_Y), .A0(D11109_Q));
KC_AOI22_X1 D11096 ( .A1(D2170_Y), .B0(D11082_Q), .B1(D10560_Y),     .Y(D11096_Y), .A0(D9265_Y));
KC_AOI22_X1 D11095 ( .A1(D11109_Q), .B0(D11013_Y), .B1(D11110_Q),     .Y(D11095_Y), .A0(D10985_Y));
KC_AOI22_X1 D11094 ( .A1(D9555_Y), .B0(D1366_Q), .B1(D10541_Y),     .Y(D11094_Y), .A0(D11104_Q));
KC_AOI22_X1 D11093 ( .A1(D11105_Q), .B0(D11013_Y), .B1(D11106_Q),     .Y(D11093_Y), .A0(D10985_Y));
KC_AOI22_X1 D11092 ( .A1(D9555_Y), .B0(D11106_Q), .B1(D10541_Y),     .Y(D11092_Y), .A0(D11105_Q));
KC_AOI22_X1 D11061 ( .A1(D10559_Y), .B0(D11075_Q), .B1(D10558_Y),     .Y(D11061_Y), .A0(D11073_Q));
KC_AOI22_X1 D11060 ( .A1(D9555_Y), .B0(D2215_Q), .B1(D10541_Y),     .Y(D11060_Y), .A0(D2216_Q));
KC_AOI22_X1 D11059 ( .A1(D10559_Y), .B0(D11084_Q), .B1(D10558_Y),     .Y(D11059_Y), .A0(D11076_Q));
KC_AOI22_X1 D11021 ( .A1(D5461_Y), .B0(D11030_Q), .B1(D10541_Y),     .Y(D11021_Y), .A0(D11035_Q));
KC_AOI22_X1 D11020 ( .A1(D11033_Q), .B0(D11013_Y), .B1(D11034_Q),     .Y(D11020_Y), .A0(D10985_Y));
KC_AOI22_X1 D11019 ( .A1(D11035_Q), .B0(D11030_Q), .B1(D11013_Y),     .Y(D11019_Y), .A0(D10985_Y));
KC_AOI22_X1 D11018 ( .A1(D11031_Q), .B0(D11013_Y), .B1(D2217_Q),     .Y(D11018_Y), .A0(D10985_Y));
KC_AOI22_X1 D11017 ( .A1(D5461_Y), .B0(D11026_Q), .B1(D10541_Y),     .Y(D11017_Y), .A0(D11056_Q));
KC_AOI22_X1 D11016 ( .A1(D11056_Q), .B0(D11013_Y), .B1(D11026_Q),     .Y(D11016_Y), .A0(D10985_Y));
KC_AOI22_X1 D11015 ( .A1(D12070_Y), .B0(D1218_Q), .B1(D11513_Y),     .Y(D11015_Y), .A0(D9725_Y));
KC_AOI22_X1 D10979 ( .A1(D2032_Y), .B0(D2250_Q), .B1(D11443_Y),     .Y(D10979_Y), .A0(D10978_Y));
KC_AOI22_X1 D10977 ( .A1(D11006_Y), .B0(D1133_Q), .B1(D10902_Y),     .Y(D10977_Y), .A0(D10993_Q));
KC_AOI22_X1 D10976 ( .A1(D10904_Y), .B0(D11470_Q), .B1(D979_Y),     .Y(D10976_Y), .A0(D1141_Q));
KC_AOI22_X1 D10974 ( .A1(D11006_Y), .B0(D10996_Q), .B1(D10902_Y),     .Y(D10974_Y), .A0(D11000_Q));
KC_AOI22_X1 D10973 ( .A1(D11000_Q), .B0(D2183_Y), .B1(D10996_Q),     .Y(D10973_Y), .A0(D11005_Y));
KC_AOI22_X1 D10970 ( .A1(D1141_Q), .B0(D10903_Y), .B1(D11470_Q),     .Y(D10970_Y), .A0(D2184_Y));
KC_AOI22_X1 D10969 ( .A1(D10999_Q), .B0(D2183_Y), .B1(D1137_Q),     .Y(D10969_Y), .A0(D11005_Y));
KC_AOI22_X1 D10968 ( .A1(D11005_Y), .B0(D1133_Q), .B1(D2183_Y),     .Y(D10968_Y), .A0(D10993_Q));
KC_AOI22_X1 D10934 ( .A1(D10889_Q), .B0(D2189_Y), .B1(D11330_Q),     .Y(D10934_Y), .A0(D10917_Y));
KC_AOI22_X1 D10933 ( .A1(D10880_Q), .B0(D2183_Y), .B1(D10888_Q),     .Y(D10933_Y), .A0(D11005_Y));
KC_AOI22_X1 D10932 ( .A1(D10890_Q), .B0(D10903_Y), .B1(D10882_Q),     .Y(D10932_Y), .A0(D2184_Y));
KC_AOI22_X1 D10931 ( .A1(D10951_Q), .B0(D2189_Y), .B1(D10954_Q),     .Y(D10931_Y), .A0(D10917_Y));
KC_AOI22_X1 D10930 ( .A1(D10886_Q), .B0(D2183_Y), .B1(D10887_Q),     .Y(D10930_Y), .A0(D11005_Y));
KC_AOI22_X1 D10928 ( .A1(D1040_Q), .B0(D2190_Y), .B1(D11400_Q),     .Y(D10928_Y), .A0(D2242_Y));
KC_AOI22_X1 D10927 ( .A1(D10950_Q), .B0(D2183_Y), .B1(D10942_Q),     .Y(D10927_Y), .A0(D11005_Y));
KC_AOI22_X1 D10925 ( .A1(D11006_Y), .B0(D10942_Q), .B1(D10902_Y),     .Y(D10925_Y), .A0(D10950_Q));
KC_AOI22_X1 D10924 ( .A1(D10990_Y), .B0(D10952_Q), .B1(D10912_Y),     .Y(D10924_Y), .A0(D10947_Q));
KC_AOI22_X1 D10923 ( .A1(D10947_Q), .B0(D2190_Y), .B1(D10952_Q),     .Y(D10923_Y), .A0(D2242_Y));
KC_AOI22_X1 D10922 ( .A1(D10948_Q), .B0(D2189_Y), .B1(D1029_Q),     .Y(D10922_Y), .A0(D10917_Y));
KC_AOI22_X1 D10921 ( .A1(D10955_Q), .B0(D10903_Y), .B1(D10944_Q),     .Y(D10921_Y), .A0(D2184_Y));
KC_AOI22_X1 D10920 ( .A1(D10904_Y), .B0(D10944_Q), .B1(D979_Y),     .Y(D10920_Y), .A0(D10955_Q));
KC_AOI22_X1 D10919 ( .A1(D1032_Q), .B0(D2189_Y), .B1(D10949_Q),     .Y(D10919_Y), .A0(D10917_Y));
KC_AOI22_X1 D10918 ( .A1(D10394_Y), .B0(D1029_Q), .B1(D10913_Y),     .Y(D10918_Y), .A0(D10948_Q));
KC_AOI22_X1 D10915 ( .A1(D10940_Q), .B0(D2189_Y), .B1(D1025_Q),     .Y(D10915_Y), .A0(D10917_Y));
KC_AOI22_X1 D10914 ( .A1(D10394_Y), .B0(D1025_Q), .B1(D10913_Y),     .Y(D10914_Y), .A0(D10940_Q));
KC_AOI22_X1 D10910 ( .A1(D10941_Q), .B0(D2189_Y), .B1(D10943_Q),     .Y(D10910_Y), .A0(D10917_Y));
KC_AOI22_X1 D10909 ( .A1(D10394_Y), .B0(D10943_Q), .B1(D10913_Y),     .Y(D10909_Y), .A0(D10941_Q));
KC_AOI22_X1 D10907 ( .A1(D11002_Q), .B0(D10903_Y), .B1(D10995_Q),     .Y(D10907_Y), .A0(D2184_Y));
KC_AOI22_X1 D10906 ( .A1(D10904_Y), .B0(D10995_Q), .B1(D979_Y),     .Y(D10906_Y), .A0(D11002_Q));
KC_AOI22_X1 D10900 ( .A1(D10904_Y), .B0(D2219_Q), .B1(D979_Y),     .Y(D10900_Y), .A0(D11001_Q));
KC_AOI22_X1 D10899 ( .A1(D11001_Q), .B0(D10903_Y), .B1(D2219_Q),     .Y(D10899_Y), .A0(D2184_Y));
KC_AOI22_X1 D10843 ( .A1(D10929_Y), .B0(D8348_Y), .B1(D11826_Y),     .Y(D10843_Y), .A0(D8345_Y));
KC_AOI22_X1 D10842 ( .A1(D10916_Y), .B0(D8348_Y), .B1(D11827_Y),     .Y(D10842_Y), .A0(D8345_Y));
KC_AOI22_X1 D10840 ( .A1(D11006_Y), .B0(D10887_Q), .B1(D10902_Y),     .Y(D10840_Y), .A0(D10886_Q));
KC_AOI22_X1 D10838 ( .A1(D2188_Y), .B0(D8348_Y), .B1(D11900_Y),     .Y(D10838_Y), .A0(D8345_Y));
KC_AOI22_X1 D10837 ( .A1(D10904_Y), .B0(D10891_Q), .B1(D979_Y),     .Y(D10837_Y), .A0(D10892_Q));
KC_AOI22_X1 D10836 ( .A1(D10904_Y), .B0(D10882_Q), .B1(D979_Y),     .Y(D10836_Y), .A0(D10890_Q));
KC_AOI22_X1 D10835 ( .A1(D10394_Y), .B0(D2255_Q), .B1(D10913_Y),     .Y(D10835_Y), .A0(D1043_Q));
KC_AOI22_X1 D10834 ( .A1(D10904_Y), .B0(D914_Q), .B1(D979_Y),     .Y(D10834_Y), .A0(D10884_Q));
KC_AOI22_X1 D10833 ( .A1(D11006_Y), .B0(D10888_Q), .B1(D10902_Y),     .Y(D10833_Y), .A0(D10880_Q));
KC_AOI22_X1 D10832 ( .A1(D11006_Y), .B0(D10883_Q), .B1(D10902_Y),     .Y(D10832_Y), .A0(D10881_Q));
KC_AOI22_X1 D10759 ( .A1(D11271_Q), .B0(D10743_Y), .B1(D808_Q),     .Y(D10759_Y), .A0(D10805_Y));
KC_AOI22_X1 D10758 ( .A1(D10749_Y), .B0(D805_Q), .B1(D10750_Y),     .Y(D10758_Y), .A0(D801_Q));
KC_AOI22_X1 D10755 ( .A1(D10710_Q), .B0(D10743_Y), .B1(D10802_Q),     .Y(D10755_Y), .A0(D10805_Y));
KC_AOI22_X1 D10752 ( .A1(D10801_Q), .B0(D10808_Y), .B1(D10800_Q),     .Y(D10752_Y), .A0(D10809_Y));
KC_AOI22_X1 D10738 ( .A1(D10692_Y), .B0(D10792_Q), .B1(D10773_Y),     .Y(D10738_Y), .A0(D8211_Y));
KC_AOI22_X1 D10737 ( .A1(D11214_Y), .B0(D10791_Q), .B1(D10772_Y),     .Y(D10737_Y), .A0(D8211_Y));
KC_AOI22_X1 D10736 ( .A1(D10760_Y), .B0(D10793_Q), .B1(D10774_Y),     .Y(D10736_Y), .A0(D8211_Y));
KC_AOI22_X1 D10733 ( .A1(D10680_Y), .B0(D10789_Q), .B1(D10769_Y),     .Y(D10733_Y), .A0(D8211_Y));
KC_AOI22_X1 D10703 ( .A1(D10724_Q), .B0(D10808_Y), .B1(D10721_Q),     .Y(D10703_Y), .A0(D10809_Y));
KC_AOI22_X1 D10702 ( .A1(D10749_Y), .B0(D10721_Q), .B1(D10750_Y),     .Y(D10702_Y), .A0(D10724_Q));
KC_AOI22_X1 D10700 ( .A1(D688_Q), .B0(D10742_Y), .B1(D10719_Q),     .Y(D10700_Y), .A0(D10745_Y));
KC_AOI22_X1 D10696 ( .A1(D10804_Y), .B0(D11180_Q), .B1(D10663_Y),     .Y(D10696_Y), .A0(D730_Q));
KC_AOI22_X1 D10695 ( .A1(D10749_Y), .B0(D689_Q), .B1(D10750_Y),     .Y(D10695_Y), .A0(D11182_Q));
KC_AOI22_X1 D10694 ( .A1(D10723_Q), .B0(D10808_Y), .B1(D10720_Q),     .Y(D10694_Y), .A0(D10809_Y));
KC_AOI22_X1 D10693 ( .A1(D10749_Y), .B0(D10720_Q), .B1(D10750_Y),     .Y(D10693_Y), .A0(D10723_Q));
KC_AOI22_X1 D10690 ( .A1(D10672_Y), .B0(D10722_Q), .B1(D10757_Y),     .Y(D10690_Y), .A0(D10234_Q));
KC_AOI22_X1 D10689 ( .A1(D10234_Q), .B0(D10742_Y), .B1(D10722_Q),     .Y(D10689_Y), .A0(D10745_Y));
KC_AOI22_X1 D10688 ( .A1(D10804_Y), .B0(D10716_Q), .B1(D10663_Y),     .Y(D10688_Y), .A0(D10714_Q));
KC_AOI22_X1 D10687 ( .A1(D730_Q), .B0(D10743_Y), .B1(D11180_Q),     .Y(D10687_Y), .A0(D10805_Y));
KC_AOI22_X1 D10686 ( .A1(D10714_Q), .B0(D10743_Y), .B1(D10716_Q),     .Y(D10686_Y), .A0(D10805_Y));
KC_AOI22_X1 D10685 ( .A1(D10672_Y), .B0(D686_Q), .B1(D10757_Y),     .Y(D10685_Y), .A0(D685_Q));
KC_AOI22_X1 D10684 ( .A1(D10804_Y), .B0(D10718_Q), .B1(D10663_Y),     .Y(D10684_Y), .A0(D10717_Q));
KC_AOI22_X1 D10683 ( .A1(D10717_Q), .B0(D10743_Y), .B1(D10718_Q),     .Y(D10683_Y), .A0(D10805_Y));
KC_AOI22_X1 D10682 ( .A1(D10672_Y), .B0(D11181_Q), .B1(D10757_Y),     .Y(D10682_Y), .A0(D11187_Q));
KC_AOI22_X1 D10679 ( .A1(D10713_Q), .B0(D10743_Y), .B1(D10708_Q),     .Y(D10679_Y), .A0(D10805_Y));
KC_AOI22_X1 D10678 ( .A1(D10804_Y), .B0(D10708_Q), .B1(D10663_Y),     .Y(D10678_Y), .A0(D10713_Q));
KC_AOI22_X1 D10677 ( .A1(D685_Q), .B0(D10742_Y), .B1(D686_Q),     .Y(D10677_Y), .A0(D10745_Y));
KC_AOI22_X1 D10674 ( .A1(D11187_Q), .B0(D10742_Y), .B1(D11181_Q),     .Y(D10674_Y), .A0(D10745_Y));
KC_AOI22_X1 D10673 ( .A1(D10709_Q), .B0(D10808_Y), .B1(D10712_Q),     .Y(D10673_Y), .A0(D10809_Y));
KC_AOI22_X1 D10671 ( .A1(D10749_Y), .B0(D10712_Q), .B1(D10750_Y),     .Y(D10671_Y), .A0(D10709_Q));
KC_AOI22_X1 D10670 ( .A1(D679_Q), .B0(D10742_Y), .B1(D10711_Q),     .Y(D10670_Y), .A0(D10745_Y));
KC_AOI22_X1 D10669 ( .A1(D10672_Y), .B0(D10711_Q), .B1(D10757_Y),     .Y(D10669_Y), .A0(D679_Q));
KC_AOI22_X1 D10668 ( .A1(D10672_Y), .B0(D11177_Q), .B1(D10757_Y),     .Y(D10668_Y), .A0(D682_Q));
KC_AOI22_X1 D10667 ( .A1(D10804_Y), .B0(D808_Q), .B1(D10663_Y),     .Y(D10667_Y), .A0(D11271_Q));
KC_AOI22_X1 D10666 ( .A1(D10672_Y), .B0(D10715_Q), .B1(D10757_Y),     .Y(D10666_Y), .A0(D680_Q));
KC_AOI22_X1 D10665 ( .A1(D680_Q), .B0(D10742_Y), .B1(D10715_Q),     .Y(D10665_Y), .A0(D10745_Y));
KC_AOI22_X1 D10662 ( .A1(D10804_Y), .B0(D10802_Q), .B1(D10663_Y),     .Y(D10662_Y), .A0(D10710_Q));
KC_AOI22_X1 D10661 ( .A1(D10749_Y), .B0(D10800_Q), .B1(D10750_Y),     .Y(D10661_Y), .A0(D10801_Q));
KC_AOI22_X1 D10640 ( .A1(D527_Q), .B0(D10818_Y), .B1(D10650_Q),     .Y(D10640_Y), .A0(D10765_Y));
KC_AOI22_X1 D10639 ( .A1(D127_Q), .B0(D10818_Y), .B1(D10184_Q),     .Y(D10639_Y), .A0(D10765_Y));
KC_AOI22_X1 D10638 ( .A1(D525_Q), .B0(D10818_Y), .B1(D2213_Q),     .Y(D10638_Y), .A0(D10765_Y));
KC_AOI22_X1 D10637 ( .A1(D10630_Q), .B0(D10818_Y), .B1(D10631_Q),     .Y(D10637_Y), .A0(D10765_Y));
KC_AOI22_X1 D10636 ( .A1(D10766_Y), .B0(D10650_Q), .B1(D10727_Y),     .Y(D10636_Y), .A0(D527_Q));
KC_AOI22_X1 D10635 ( .A1(D10185_Q), .B0(D10818_Y), .B1(D10183_Q),     .Y(D10635_Y), .A0(D10765_Y));
KC_AOI22_X1 D10609 ( .A1(D9555_Y), .B0(D1363_Q), .B1(D10541_Y),     .Y(D10609_Y), .A0(D10612_Q));
KC_AOI22_X1 D10608 ( .A1(D9555_Y), .B0(D10615_Q), .B1(D10541_Y),     .Y(D10608_Y), .A0(D10611_Q));
KC_AOI22_X1 D10607 ( .A1(D10612_Q), .B0(D11013_Y), .B1(D1363_Q),     .Y(D10607_Y), .A0(D10985_Y));
KC_AOI22_X1 D10606 ( .A1(D9555_Y), .B0(D10613_Q), .B1(D10541_Y),     .Y(D10606_Y), .A0(D10610_Q));
KC_AOI22_X1 D10605 ( .A1(D11104_Q), .B0(D11013_Y), .B1(D1366_Q),     .Y(D10605_Y), .A0(D10985_Y));
KC_AOI22_X1 D10604 ( .A1(D10611_Q), .B0(D11013_Y), .B1(D10615_Q),     .Y(D10604_Y), .A0(D10985_Y));
KC_AOI22_X1 D10589 ( .A1(D2170_Y), .B0(D11085_Q), .B1(D10560_Y),     .Y(D10589_Y), .A0(D11083_Q));
KC_AOI22_X1 D10588 ( .A1(D10559_Y), .B0(D10601_Q), .B1(D10558_Y),     .Y(D10588_Y), .A0(D10598_Q));
KC_AOI22_X1 D10587 ( .A1(D1144_Y), .B0(D1315_Q), .B1(D10535_Y),     .Y(D10587_Y), .A0(D10602_Q));
KC_AOI22_X1 D10586 ( .A1(D11074_Q), .B0(D11009_Y), .B1(D1309_Q),     .Y(D10586_Y), .A0(D11003_Y));
KC_AOI22_X1 D10582 ( .A1(D11078_Q), .B0(D11011_Y), .B1(D11077_Q),     .Y(D10582_Y), .A0(D11010_Y));
KC_AOI22_X1 D10581 ( .A1(D11079_Q), .B0(D11012_Y), .B1(D11080_Q),     .Y(D10581_Y), .A0(D11014_Y));
KC_AOI22_X1 D10580 ( .A1(D10559_Y), .B0(D11077_Q), .B1(D10558_Y),     .Y(D10580_Y), .A0(D11078_Q));
KC_AOI22_X1 D10578 ( .A1(D10598_Q), .B0(D11011_Y), .B1(D10601_Q),     .Y(D10578_Y), .A0(D11010_Y));
KC_AOI22_X1 D10577 ( .A1(D10602_Q), .B0(D11009_Y), .B1(D1315_Q),     .Y(D10577_Y), .A0(D11003_Y));
KC_AOI22_X1 D10576 ( .A1(D11076_Q), .B0(D11011_Y), .B1(D11084_Q),     .Y(D10576_Y), .A0(D11010_Y));
KC_AOI22_X1 D10575 ( .A1(D1144_Y), .B0(D1309_Q), .B1(D10535_Y),     .Y(D10575_Y), .A0(D11074_Q));
KC_AOI22_X1 D10574 ( .A1(D11083_Q), .B0(D11012_Y), .B1(D11085_Q),     .Y(D10574_Y), .A0(D11014_Y));
KC_AOI22_X1 D10573 ( .A1(D1144_Y), .B0(D10551_Q), .B1(D10535_Y),     .Y(D10573_Y), .A0(D10554_Q));
KC_AOI22_X1 D10572 ( .A1(D1144_Y), .B0(D10595_Q), .B1(D10535_Y),     .Y(D10572_Y), .A0(D9884_Q));
KC_AOI22_X1 D10571 ( .A1(D10599_Q), .B0(D11012_Y), .B1(D10597_Q),     .Y(D10571_Y), .A0(D11014_Y));
KC_AOI22_X1 D10570 ( .A1(D10603_Q), .B0(D11009_Y), .B1(D10600_Q),     .Y(D10570_Y), .A0(D11003_Y));
KC_AOI22_X1 D10567 ( .A1(D1144_Y), .B0(D10600_Q), .B1(D10535_Y),     .Y(D10567_Y), .A0(D10603_Q));
KC_AOI22_X1 D10566 ( .A1(D2170_Y), .B0(D10597_Q), .B1(D10560_Y),     .Y(D10566_Y), .A0(D10599_Q));
KC_AOI22_X1 D10564 ( .A1(D10594_Q), .B0(D11012_Y), .B1(D10596_Q),     .Y(D10564_Y), .A0(D11014_Y));
KC_AOI22_X1 D10561 ( .A1(D10552_Q), .B0(D11009_Y), .B1(D10555_Q),     .Y(D10561_Y), .A0(D11003_Y));
KC_AOI22_X1 D10540 ( .A1(D10553_Q), .B0(D11011_Y), .B1(D1221_Q),     .Y(D10540_Y), .A0(D11010_Y));
KC_AOI22_X1 D10539 ( .A1(D11010_Y), .B0(D1220_Q), .B1(D11011_Y),     .Y(D10539_Y), .A0(D1215_Q));
KC_AOI22_X1 D10538 ( .A1(D10559_Y), .B0(D11027_Q), .B1(D10558_Y),     .Y(D10538_Y), .A0(D1223_Q));
KC_AOI22_X1 D10537 ( .A1(D1223_Q), .B0(D11011_Y), .B1(D11027_Q),     .Y(D10537_Y), .A0(D11010_Y));
KC_AOI22_X1 D10534 ( .A1(D1144_Y), .B0(D10545_Q), .B1(D10535_Y),     .Y(D10534_Y), .A0(D10547_Q));
KC_AOI22_X1 D10533 ( .A1(D10559_Y), .B0(D1221_Q), .B1(D10558_Y),     .Y(D10533_Y), .A0(D10553_Q));
KC_AOI22_X1 D10532 ( .A1(D10559_Y), .B0(D1220_Q), .B1(D10558_Y),     .Y(D10532_Y), .A0(D1215_Q));
KC_AOI22_X1 D10529 ( .A1(D10550_Q), .B0(D11012_Y), .B1(D1226_Q),     .Y(D10529_Y), .A0(D11014_Y));
KC_AOI22_X1 D10528 ( .A1(D2170_Y), .B0(D1226_Q), .B1(D10560_Y),     .Y(D10528_Y), .A0(D10550_Q));
KC_AOI22_X1 D10527 ( .A1(D11003_Y), .B0(D10545_Q), .B1(D11009_Y),     .Y(D10527_Y), .A0(D10547_Q));
KC_AOI22_X1 D10526 ( .A1(D1144_Y), .B0(D10555_Q), .B1(D10535_Y),     .Y(D10526_Y), .A0(D10552_Q));
KC_AOI22_X1 D10525 ( .A1(D2170_Y), .B0(D2159_Q), .B1(D10560_Y),     .Y(D10525_Y), .A0(D10544_Q));
KC_AOI22_X1 D10524 ( .A1(D10549_Q), .B0(D11009_Y), .B1(D10548_Q),     .Y(D10524_Y), .A0(D11003_Y));
KC_AOI22_X1 D10523 ( .A1(D1144_Y), .B0(D10548_Q), .B1(D10535_Y),     .Y(D10523_Y), .A0(D10549_Q));
KC_AOI22_X1 D10469 ( .A1(D2170_Y), .B0(D10510_Q), .B1(D10560_Y),     .Y(D10469_Y), .A0(D10511_Q));
KC_AOI22_X1 D10468 ( .A1(D10511_Q), .B0(D11012_Y), .B1(D10510_Q),     .Y(D10468_Y), .A0(D11014_Y));
KC_AOI22_X1 D10461 ( .A1(D10546_Q), .B0(D11009_Y), .B1(D2156_Q),     .Y(D10461_Y), .A0(D11003_Y));
KC_AOI22_X1 D10390 ( .A1(D10422_Q), .B0(D10903_Y), .B1(D10424_Q),     .Y(D10390_Y), .A0(D2184_Y));
KC_AOI22_X1 D10445 ( .A1(D10426_Q), .B0(D10903_Y), .B1(D10425_Q),     .Y(D10445_Y), .A0(D2184_Y));
KC_AOI22_X1 D10444 ( .A1(D10990_Y), .B0(D10430_Q), .B1(D10912_Y),     .Y(D10444_Y), .A0(D10431_Q));
KC_AOI22_X1 D10443 ( .A1(D10394_Y), .B0(D10885_Q), .B1(D10913_Y),     .Y(D10443_Y), .A0(D913_Q));
KC_AOI22_X1 D10442 ( .A1(D10904_Y), .B0(D10428_Q), .B1(D979_Y),     .Y(D10442_Y), .A0(D10429_Q));
KC_AOI22_X1 D10441 ( .A1(D10904_Y), .B0(D10424_Q), .B1(D979_Y),     .Y(D10441_Y), .A0(D10422_Q));
KC_AOI22_X1 D10406 ( .A1(D133_Q), .B0(D2190_Y), .B1(D911_Q),     .Y(D10406_Y), .A0(D2242_Y));
KC_AOI22_X1 D10405 ( .A1(D10352_Q), .B0(D2190_Y), .B1(D917_Q),     .Y(D10405_Y), .A0(D2242_Y));
KC_AOI22_X1 D10404 ( .A1(D10990_Y), .B0(D911_Q), .B1(D10912_Y),     .Y(D10404_Y), .A0(D133_Q));
KC_AOI22_X1 D10403 ( .A1(D10427_Q), .B0(D2189_Y), .B1(D1037_Q),     .Y(D10403_Y), .A0(D10917_Y));
KC_AOI22_X1 D10401 ( .A1(D10394_Y), .B0(D1037_Q), .B1(D10913_Y),     .Y(D10401_Y), .A0(D10427_Q));
KC_AOI22_X1 D10398 ( .A1(D10394_Y), .B0(D10946_Q), .B1(D10913_Y),     .Y(D10398_Y), .A0(D1028_Q));
KC_AOI22_X1 D10397 ( .A1(D1028_Q), .B0(D2189_Y), .B1(D10946_Q),     .Y(D10397_Y), .A0(D10917_Y));
KC_AOI22_X1 D10396 ( .A1(D10394_Y), .B0(D10949_Q), .B1(D10913_Y),     .Y(D10396_Y), .A0(D1032_Q));
KC_AOI22_X1 D10395 ( .A1(D10904_Y), .B0(D10425_Q), .B1(D979_Y),     .Y(D10395_Y), .A0(D10426_Q));
KC_AOI22_X1 D10393 ( .A1(D2161_Q), .B0(D10903_Y), .B1(D10423_Q),     .Y(D10393_Y), .A0(D2184_Y));
KC_AOI22_X1 D10392 ( .A1(D10904_Y), .B0(D10423_Q), .B1(D979_Y),     .Y(D10392_Y), .A0(D2161_Q));
KC_AOI22_X1 D10387 ( .A1(D10990_Y), .B0(D10354_Q), .B1(D10912_Y),     .Y(D10387_Y), .A0(D10353_Q));
KC_AOI22_X1 D10386 ( .A1(D913_Q), .B0(D2189_Y), .B1(D10885_Q),     .Y(D10386_Y), .A0(D10917_Y));
KC_AOI22_X1 D10382 ( .A1(D11006_Y), .B0(D10417_Q), .B1(D10902_Y),     .Y(D10382_Y), .A0(D1013_Q));
KC_AOI22_X1 D10381 ( .A1(D9707_Q), .B0(D2183_Y), .B1(D10419_Q),     .Y(D10381_Y), .A0(D11005_Y));
KC_AOI22_X1 D10380 ( .A1(D11006_Y), .B0(D10419_Q), .B1(D10902_Y),     .Y(D10380_Y), .A0(D9707_Q));
KC_AOI22_X1 D10379 ( .A1(D10429_Q), .B0(D10903_Y), .B1(D10428_Q),     .Y(D10379_Y), .A0(D2184_Y));
KC_AOI22_X1 D10378 ( .A1(D1021_Q), .B0(D2183_Y), .B1(D10420_Q),     .Y(D10378_Y), .A0(D11005_Y));
KC_AOI22_X1 D10377 ( .A1(D11006_Y), .B0(D10418_Q), .B1(D10902_Y),     .Y(D10377_Y), .A0(D1016_Q));
KC_AOI22_X1 D10375 ( .A1(D1013_Q), .B0(D2183_Y), .B1(D10417_Q),     .Y(D10375_Y), .A0(D11005_Y));
KC_AOI22_X1 D10317 ( .A1(D10347_Q), .B0(D2190_Y), .B1(D10350_Q),     .Y(D10317_Y), .A0(D2242_Y));
KC_AOI22_X1 D10257 ( .A1(D1983_Y), .B0(D10201_Y), .B1(D9393_Y),     .Y(D10257_Y), .A0(D10302_Q));
KC_AOI22_X1 D10256 ( .A1(D1992_Y), .B0(D10681_Y), .B1(D9393_Y),     .Y(D10256_Y), .A0(D10294_Q));
KC_AOI22_X1 D10255 ( .A1(D1992_Y), .B0(D11228_Y), .B1(D9393_Y),     .Y(D10255_Y), .A0(D10296_Q));
KC_AOI22_X1 D10254 ( .A1(D1992_Y), .B0(D10291_Y), .B1(D9393_Y),     .Y(D10254_Y), .A0(D10303_Q));
KC_AOI22_X1 D10253 ( .A1(D1992_Y), .B0(D12319_Y), .B1(D9393_Y),     .Y(D10253_Y), .A0(D10302_Q));
KC_AOI22_X1 D10252 ( .A1(D1992_Y), .B0(D10794_Y), .B1(D9393_Y),     .Y(D10252_Y), .A0(D10300_Q));
KC_AOI22_X1 D10251 ( .A1(D1992_Y), .B0(D10797_Y), .B1(D9393_Y),     .Y(D10251_Y), .A0(D10299_Q));
KC_AOI22_X1 D10250 ( .A1(D1992_Y), .B0(D10751_Y), .B1(D9393_Y),     .Y(D10250_Y), .A0(D10301_Q));
KC_AOI22_X1 D10249 ( .A1(D1992_Y), .B0(D12320_Y), .B1(D9393_Y),     .Y(D10249_Y), .A0(D10311_Q));
KC_AOI22_X1 D10245 ( .A1(D1983_Y), .B0(D11276_Y), .B1(D9393_Y),     .Y(D10245_Y), .A0(D825_Q));
KC_AOI22_X1 D10230 ( .A1(D1983_Y), .B0(D10178_Y), .B1(D9393_Y),     .Y(D10230_Y), .A0(D10296_Q));
KC_AOI22_X1 D10199 ( .A1(D1983_Y), .B0(D11212_Y), .B1(D9393_Y),     .Y(D10199_Y), .A0(D10303_Q));
KC_AOI22_X1 D10198 ( .A1(D1983_Y), .B0(D11146_Y), .B1(D9393_Y),     .Y(D10198_Y), .A0(D10301_Q));
KC_AOI22_X1 D10135 ( .A1(D10136_Y), .B0(D11623_Y), .B1(D10137_Y),     .Y(D10135_Y), .A0(D12294_Y));
KC_AOI22_X1 D10036 ( .A1(D10032_Q), .B0(D8901_Y), .B1(D10047_Q),     .Y(D10036_Y), .A0(D8900_Y));
KC_AOI22_X1 D10019 ( .A1(D10051_Q), .B0(D8901_Y), .B1(D10009_Q),     .Y(D10019_Y), .A0(D9990_Y));
KC_AOI22_X1 D10018 ( .A1(D16790_Y), .B0(D2070_Y), .B1(D10033_Q),     .Y(D10018_Y), .A0(D7394_Y));
KC_AOI22_X1 D10016 ( .A1(D8237_Y), .B0(D2070_Y), .B1(D10051_Q),     .Y(D10016_Y), .A0(D7394_Y));
KC_AOI22_X1 D10015 ( .A1(D10033_Q), .B0(D8901_Y), .B1(D10032_Q),     .Y(D10015_Y), .A0(D8900_Y));
KC_AOI22_X1 D10014 ( .A1(D295_Y), .B0(D2070_Y), .B1(D10032_Q),     .Y(D10014_Y), .A0(D7394_Y));
KC_AOI22_X1 D10013 ( .A1(D10051_Q), .B0(D8901_Y), .B1(D10033_Q),     .Y(D10013_Y), .A0(D8900_Y));
KC_AOI22_X1 D10012 ( .A1(D7393_Y), .B0(D7313_Y), .B1(D10048_Q),     .Y(D10012_Y), .A0(D6248_Q));
KC_AOI22_X1 D10010 ( .A1(D10049_Q), .B0(D8901_Y), .B1(D10031_Q),     .Y(D10010_Y), .A0(D9990_Y));
KC_AOI22_X1 D10001 ( .A1(D230_Q), .B0(D8901_Y), .B1(D9984_Q),     .Y(D10001_Y), .A0(D8900_Y));
KC_AOI22_X1 D9997 ( .A1(D9099_Y), .B0(D2070_Y), .B1(D230_Q),     .Y(D9997_Y), .A0(D7393_Y));
KC_AOI22_X1 D9993 ( .A1(D10007_Q), .B0(D9990_Y), .B1(D2166_Q),     .Y(D9993_Y), .A0(D8900_Y));
KC_AOI22_X1 D9991 ( .A1(D9983_Q), .B0(D8901_Y), .B1(D10007_Q),     .Y(D9991_Y), .A0(D9990_Y));
KC_AOI22_X1 D9989 ( .A1(D10032_Q), .B0(D8901_Y), .B1(D2166_Q),     .Y(D9989_Y), .A0(D9990_Y));
KC_AOI22_X1 D9988 ( .A1(D10048_Q), .B0(D9990_Y), .B1(D10009_Q),     .Y(D9988_Y), .A0(D8900_Y));
KC_AOI22_X1 D9898 ( .A1(D9905_Q), .B0(D11013_Y), .B1(D9903_Q),     .Y(D9898_Y), .A0(D10985_Y));
KC_AOI22_X1 D9897 ( .A1(D9555_Y), .B0(D9903_Q), .B1(D10541_Y),     .Y(D9897_Y), .A0(D9905_Q));
KC_AOI22_X1 D9896 ( .A1(D1354_Q), .B0(D11013_Y), .B1(D1351_Q),     .Y(D9896_Y), .A0(D10985_Y));
KC_AOI22_X1 D9895 ( .A1(D9555_Y), .B0(D1351_Q), .B1(D10541_Y),     .Y(D9895_Y), .A0(D1354_Q));
KC_AOI22_X1 D9891 ( .A1(D10559_Y), .B0(D9880_Q), .B1(D10558_Y),     .Y(D9891_Y), .A0(D9883_Q));
KC_AOI22_X1 D9875 ( .A1(D1144_Y), .B0(D9886_Q), .B1(D10535_Y),     .Y(D9875_Y), .A0(D9888_Q));
KC_AOI22_X1 D9873 ( .A1(D1144_Y), .B0(D9887_Q), .B1(D10535_Y),     .Y(D9873_Y), .A0(D9885_Q));
KC_AOI22_X1 D9872 ( .A1(D9884_Q), .B0(D11009_Y), .B1(D10595_Q),     .Y(D9872_Y), .A0(D11003_Y));
KC_AOI22_X1 D9869 ( .A1(D8643_Q), .B0(D11009_Y), .B1(D8640_Q),     .Y(D9869_Y), .A0(D11003_Y));
KC_AOI22_X1 D9868 ( .A1(D9885_Q), .B0(D11009_Y), .B1(D9887_Q),     .Y(D9868_Y), .A0(D11003_Y));
KC_AOI22_X1 D9867 ( .A1(D9883_Q), .B0(D11011_Y), .B1(D9880_Q),     .Y(D9867_Y), .A0(D11010_Y));
KC_AOI22_X1 D9866 ( .A1(D9888_Q), .B0(D11009_Y), .B1(D9886_Q),     .Y(D9866_Y), .A0(D11003_Y));
KC_AOI22_X1 D9865 ( .A1(D9882_Q), .B0(D11011_Y), .B1(D9881_Q),     .Y(D9865_Y), .A0(D11010_Y));
KC_AOI22_X1 D9864 ( .A1(D10559_Y), .B0(D9881_Q), .B1(D10558_Y),     .Y(D9864_Y), .A0(D9882_Q));
KC_AOI22_X1 D9863 ( .A1(D10559_Y), .B0(D1297_Q), .B1(D10558_Y),     .Y(D9863_Y), .A0(D1290_Q));
KC_AOI22_X1 D9861 ( .A1(D8637_Q), .B0(D11011_Y), .B1(D1289_Q),     .Y(D9861_Y), .A0(D11010_Y));
KC_AOI22_X1 D9860 ( .A1(D2170_Y), .B0(D9879_Q), .B1(D10560_Y),     .Y(D9860_Y), .A0(D9878_Q));
KC_AOI22_X1 D9859 ( .A1(D9878_Q), .B0(D11012_Y), .B1(D9879_Q),     .Y(D9859_Y), .A0(D11014_Y));
KC_AOI22_X1 D9858 ( .A1(D2170_Y), .B0(D10596_Q), .B1(D10560_Y),     .Y(D9858_Y), .A0(D10594_Q));
KC_AOI22_X1 D9857 ( .A1(D9909_Q), .B0(D11012_Y), .B1(D8656_Q),     .Y(D9857_Y), .A0(D11014_Y));
KC_AOI22_X1 D9856 ( .A1(D10559_Y), .B0(D1289_Q), .B1(D10558_Y),     .Y(D9856_Y), .A0(D8637_Q));
KC_AOI22_X1 D9855 ( .A1(D10559_Y), .B0(D8632_Q), .B1(D10558_Y),     .Y(D9855_Y), .A0(D8635_Q));
KC_AOI22_X1 D9854 ( .A1(D2170_Y), .B0(D8656_Q), .B1(D10560_Y),     .Y(D9854_Y), .A0(D9909_Q));
KC_AOI22_X1 D9853 ( .A1(D9908_Q), .B0(D11012_Y), .B1(D9876_Q),     .Y(D9853_Y), .A0(D11014_Y));
KC_AOI22_X1 D9852 ( .A1(D10617_Q), .B0(D11012_Y), .B1(D9877_Q),     .Y(D9852_Y), .A0(D11014_Y));
KC_AOI22_X1 D9851 ( .A1(D2170_Y), .B0(D9877_Q), .B1(D10560_Y),     .Y(D9851_Y), .A0(D10617_Q));
KC_AOI22_X1 D9829 ( .A1(D5461_Y), .B0(D9838_Q), .B1(D10541_Y),     .Y(D9829_Y), .A0(D9836_Q));
KC_AOI22_X1 D9828 ( .A1(D1205_Q), .B0(D11013_Y), .B1(D1204_Q),     .Y(D9828_Y), .A0(D10985_Y));
KC_AOI22_X1 D9827 ( .A1(D5461_Y), .B0(D1204_Q), .B1(D10541_Y),     .Y(D9827_Y), .A0(D1205_Q));
KC_AOI22_X1 D9826 ( .A1(D5461_Y), .B0(D2078_Q), .B1(D10541_Y),     .Y(D9826_Y), .A0(D9842_Q));
KC_AOI22_X1 D9825 ( .A1(D9842_Q), .B0(D11013_Y), .B1(D2078_Q),     .Y(D9825_Y), .A0(D10985_Y));
KC_AOI22_X1 D9824 ( .A1(D9836_Q), .B0(D11013_Y), .B1(D9838_Q),     .Y(D9824_Y), .A0(D10985_Y));
KC_AOI22_X1 D9821 ( .A1(D8588_Q), .B0(D11012_Y), .B1(D122_Q),     .Y(D9821_Y), .A0(D11014_Y));
KC_AOI22_X1 D9819 ( .A1(D2170_Y), .B0(D122_Q), .B1(D10560_Y),     .Y(D9819_Y), .A0(D8588_Q));
KC_AOI22_X1 D9818 ( .A1(D8591_Q), .B0(D11009_Y), .B1(D8593_Q),     .Y(D9818_Y), .A0(D11003_Y));
KC_AOI22_X1 D9817 ( .A1(D1208_Q), .B0(D11009_Y), .B1(D1209_Q),     .Y(D9817_Y), .A0(D11003_Y));
KC_AOI22_X1 D9816 ( .A1(D1199_Q), .B0(D11012_Y), .B1(D1301_Q),     .Y(D9816_Y), .A0(D11014_Y));
KC_AOI22_X1 D9815 ( .A1(D9834_Q), .B0(D11012_Y), .B1(D2082_Q),     .Y(D9815_Y), .A0(D11014_Y));
KC_AOI22_X1 D9814 ( .A1(D9840_Q), .B0(D11009_Y), .B1(D9841_Q),     .Y(D9814_Y), .A0(D11003_Y));
KC_AOI22_X1 D9813 ( .A1(D2170_Y), .B0(D2082_Q), .B1(D10560_Y),     .Y(D9813_Y), .A0(D9834_Q));
KC_AOI22_X1 D9812 ( .A1(D2170_Y), .B0(D1301_Q), .B1(D10560_Y),     .Y(D9812_Y), .A0(D1199_Q));
KC_AOI22_X1 D9808 ( .A1(D1144_Y), .B0(D8593_Q), .B1(D10535_Y),     .Y(D9808_Y), .A0(D8591_Q));
KC_AOI22_X1 D9807 ( .A1(D1144_Y), .B0(D1209_Q), .B1(D10535_Y),     .Y(D9807_Y), .A0(D1208_Q));
KC_AOI22_X1 D9806 ( .A1(D10559_Y), .B0(D2084_Q), .B1(D10558_Y),     .Y(D9806_Y), .A0(D2085_Q));
KC_AOI22_X1 D9805 ( .A1(D2085_Q), .B0(D11011_Y), .B1(D2084_Q),     .Y(D9805_Y), .A0(D11010_Y));
KC_AOI22_X1 D9804 ( .A1(D1144_Y), .B0(D9841_Q), .B1(D10535_Y),     .Y(D9804_Y), .A0(D9840_Q));
KC_AOI22_X1 D9803 ( .A1(D10559_Y), .B0(D2083_Q), .B1(D10558_Y),     .Y(D9803_Y), .A0(D9892_Q));
KC_AOI22_X1 D9802 ( .A1(D1302_Q), .B0(D11011_Y), .B1(D1303_Q),     .Y(D9802_Y), .A0(D11010_Y));
KC_AOI22_X1 D9801 ( .A1(D10559_Y), .B0(D9890_Q), .B1(D10558_Y),     .Y(D9801_Y), .A0(D9889_Q));
KC_AOI22_X1 D9800 ( .A1(D9889_Q), .B0(D11011_Y), .B1(D9890_Q),     .Y(D9800_Y), .A0(D11010_Y));
KC_AOI22_X1 D9799 ( .A1(D9892_Q), .B0(D11011_Y), .B1(D2083_Q),     .Y(D9799_Y), .A0(D11010_Y));
KC_AOI22_X1 D9680 ( .A1(D10394_Y), .B0(D9611_Q), .B1(D10913_Y),     .Y(D9680_Y), .A0(D9606_Q));
KC_AOI22_X1 D9679 ( .A1(D9606_Q), .B0(D2189_Y), .B1(D9611_Q),     .Y(D9679_Y), .A0(D10917_Y));
KC_AOI22_X1 D9677 ( .A1(D10394_Y), .B0(D9613_Q), .B1(D10913_Y),     .Y(D9677_Y), .A0(D9612_Q));
KC_AOI22_X1 D9676 ( .A1(D10394_Y), .B0(D9614_Q), .B1(D10913_Y),     .Y(D9676_Y), .A0(D9608_Q));
KC_AOI22_X1 D9675 ( .A1(D9612_Q), .B0(D2189_Y), .B1(D9613_Q),     .Y(D9675_Y), .A0(D10917_Y));
KC_AOI22_X1 D9674 ( .A1(D9607_Q), .B0(D2189_Y), .B1(D9610_Q),     .Y(D9674_Y), .A0(D10917_Y));
KC_AOI22_X1 D9673 ( .A1(D10394_Y), .B0(D9610_Q), .B1(D10913_Y),     .Y(D9673_Y), .A0(D9607_Q));
KC_AOI22_X1 D9669 ( .A1(D10904_Y), .B0(D1020_Q), .B1(D979_Y),     .Y(D9669_Y), .A0(D1022_Q));
KC_AOI22_X1 D9665 ( .A1(D10904_Y), .B0(D9712_Q), .B1(D979_Y),     .Y(D9665_Y), .A0(D2080_Q));
KC_AOI22_X1 D9664 ( .A1(D10904_Y), .B0(D9714_Q), .B1(D979_Y),     .Y(D9664_Y), .A0(D9717_Q));
KC_AOI22_X1 D9663 ( .A1(D10904_Y), .B0(D9711_Q), .B1(D979_Y),     .Y(D9663_Y), .A0(D2081_Q));
KC_AOI22_X1 D9662 ( .A1(D1022_Q), .B0(D10903_Y), .B1(D1020_Q),     .Y(D9662_Y), .A0(D2184_Y));
KC_AOI22_X1 D9659 ( .A1(D2080_Q), .B0(D10903_Y), .B1(D9712_Q),     .Y(D9659_Y), .A0(D2184_Y));
KC_AOI22_X1 D9658 ( .A1(D9717_Q), .B0(D10903_Y), .B1(D9714_Q),     .Y(D9658_Y), .A0(D2184_Y));
KC_AOI22_X1 D9657 ( .A1(D2081_Q), .B0(D10903_Y), .B1(D9711_Q),     .Y(D9657_Y), .A0(D2184_Y));
KC_AOI22_X1 D9656 ( .A1(D11006_Y), .B0(D9706_Q), .B1(D10902_Y),     .Y(D9656_Y), .A0(D9703_Q));
KC_AOI22_X1 D9655 ( .A1(D9709_Q), .B0(D2183_Y), .B1(D9710_Q),     .Y(D9655_Y), .A0(D11005_Y));
KC_AOI22_X1 D9654 ( .A1(D1018_Q), .B0(D2183_Y), .B1(D1015_Q),     .Y(D9654_Y), .A0(D11005_Y));
KC_AOI22_X1 D9653 ( .A1(D11006_Y), .B0(D1015_Q), .B1(D10902_Y),     .Y(D9653_Y), .A0(D1018_Q));
KC_AOI22_X1 D9652 ( .A1(D11006_Y), .B0(D9710_Q), .B1(D10902_Y),     .Y(D9652_Y), .A0(D9709_Q));
KC_AOI22_X1 D9651 ( .A1(D9705_Q), .B0(D2183_Y), .B1(D9708_Q),     .Y(D9651_Y), .A0(D11005_Y));
KC_AOI22_X1 D9650 ( .A1(D11006_Y), .B0(D9708_Q), .B1(D10902_Y),     .Y(D9650_Y), .A0(D9705_Q));
KC_AOI22_X1 D9649 ( .A1(D9703_Q), .B0(D2183_Y), .B1(D9706_Q),     .Y(D9649_Y), .A0(D11005_Y));
KC_AOI22_X1 D9596 ( .A1(D904_Q), .B0(D2190_Y), .B1(D905_Q),     .Y(D9596_Y), .A0(D2242_Y));
KC_AOI22_X1 D9595 ( .A1(D10990_Y), .B0(D10350_Q), .B1(D10912_Y),     .Y(D9595_Y), .A0(D10347_Q));
KC_AOI22_X1 D9594 ( .A1(D9608_Q), .B0(D2189_Y), .B1(D9614_Q),     .Y(D9594_Y), .A0(D10917_Y));
KC_AOI22_X1 D9529 ( .A1(D1992_Y), .B0(D2119_Y), .B1(D9393_Y),     .Y(D9529_Y), .A0(D827_Q));
KC_AOI22_X1 D9388 ( .A1(D9518_Y), .B0(D8105_Y), .B1(D9550_Y),     .Y(D9388_Y), .A0(D8079_Y));
KC_AOI22_X1 D9307 ( .A1(D9301_Y), .B0(D9181_Y), .B1(D7896_Q),     .Y(D9307_Y), .A0(D7631_Y));
KC_AOI22_X1 D9305 ( .A1(D13097_Q), .B0(D9114_Y), .B1(D484_Q),     .Y(D9305_Y), .A0(D7631_Y));
KC_AOI22_X1 D9304 ( .A1(D9325_Q), .B0(D6077_Y), .B1(D9322_Q),     .Y(D9304_Y), .A0(D9114_Y));
KC_AOI22_X1 D9303 ( .A1(D9340_Y), .B0(D6077_Y), .B1(D9361_Q),     .Y(D9303_Y), .A0(D7631_Y));
KC_AOI22_X1 D9239 ( .A1(D7638_Y), .B0(D9181_Y), .B1(D7819_Y),     .Y(D9239_Y), .A0(D1918_Y));
KC_AOI22_X1 D9233 ( .A1(D154_Q), .B0(D9114_Y), .B1(D2094_Q),     .Y(D9233_Y), .A0(D9181_Y));
KC_AOI22_X1 D9232 ( .A1(D10164_Y), .B0(D7823_Y), .B1(D9181_Y),     .Y(D9232_Y), .A0(D7631_Y));
KC_AOI22_X1 D9189 ( .A1(D9159_Q), .B0(D9114_Y), .B1(D451_Q),     .Y(D9189_Y), .A0(D7499_Y));
KC_AOI22_X1 D9188 ( .A1(D419_Q), .B0(D9102_Y), .B1(D9215_Q),     .Y(D9188_Y), .A0(D5969_Y));
KC_AOI22_X1 D9185 ( .A1(D9218_Q), .B0(D9221_Q), .B1(D9102_Y),     .Y(D9185_Y), .A0(D5969_Y));
KC_AOI22_X1 D9184 ( .A1(D7638_Y), .B0(D6077_Y), .B1(D10143_Y),     .Y(D9184_Y), .A0(D7709_Y));
KC_AOI22_X1 D9183 ( .A1(D10109_Q), .B0(D6077_Y), .B1(D442_Q),     .Y(D9183_Y), .A0(D9102_Y));
KC_AOI22_X1 D9177 ( .A1(D9216_Q), .B0(D9114_Y), .B1(D449_Q),     .Y(D9177_Y), .A0(D7499_Y));
KC_AOI22_X1 D9173 ( .A1(D7638_Y), .B0(D6077_Y), .B1(D7477_Q),     .Y(D9173_Y), .A0(D7710_Y));
KC_AOI22_X1 D9170 ( .A1(D10108_Q), .B0(D6077_Y), .B1(D414_Q),     .Y(D9170_Y), .A0(D5969_Y));
KC_AOI22_X1 D9169 ( .A1(D9274_Q), .B0(D9102_Y), .B1(D9220_Q),     .Y(D9169_Y), .A0(D7499_Y));
KC_AOI22_X1 D9124 ( .A1(D9198_Y), .B0(D7494_Y), .B1(D9273_Q),     .Y(D9124_Y), .A0(D9068_Y));
KC_AOI22_X1 D9071 ( .A1(D40_Q), .B0(D7473_Y), .B1(D8063_Y),     .Y(D9071_Y), .A0(D9041_Y));
KC_AOI22_X1 D9063 ( .A1(D1864_Y), .B0(D308_Y), .B1(D8063_Y),     .Y(D9063_Y), .A0(D9160_Q));
KC_AOI22_X1 D9062 ( .A1(D7362_Y), .B0(D8071_Y), .B1(D350_Y),     .Y(D9062_Y), .A0(D9482_Y));
KC_AOI22_X1 D9060 ( .A1(D10061_Q), .B0(D7494_Y), .B1(D10062_Q),     .Y(D9060_Y), .A0(D9054_Y));
KC_AOI22_X1 D9051 ( .A1(D8069_Y), .B0(D9054_Y), .B1(D8952_Q),     .Y(D9051_Y), .A0(D7473_Y));
KC_AOI22_X1 D9049 ( .A1(D8062_Y), .B0(D7494_Y), .B1(D9280_Q),     .Y(D9049_Y), .A0(D7473_Y));
KC_AOI22_X1 D9048 ( .A1(D7957_Y), .B0(D7494_Y), .B1(D353_Q),     .Y(D9048_Y), .A0(D7473_Y));
KC_AOI22_X1 D9046 ( .A1(D615_Y), .B0(D7494_Y), .B1(D10059_Q),     .Y(D9046_Y), .A0(D7473_Y));
KC_AOI22_X1 D9044 ( .A1(D7481_Q), .B0(D9054_Y), .B1(D10060_Q),     .Y(D9044_Y), .A0(D9041_Y));
KC_AOI22_X1 D9043 ( .A1(D9021_Q), .B0(D7494_Y), .B1(D10058_Q),     .Y(D9043_Y), .A0(D9041_Y));
KC_AOI22_X1 D9038 ( .A1(D8066_Y), .B0(D308_Y), .B1(D8069_Y),     .Y(D9038_Y), .A0(D7473_Y));
KC_AOI22_X1 D9037 ( .A1(D8065_Y), .B0(D308_Y), .B1(D7957_Y),     .Y(D9037_Y), .A0(D7473_Y));
KC_AOI22_X1 D9036 ( .A1(D8953_Q), .B0(D7473_Y), .B1(D8064_Y),     .Y(D9036_Y), .A0(D9041_Y));
KC_AOI22_X1 D9035 ( .A1(D8070_Y), .B0(D7494_Y), .B1(D354_Q),     .Y(D9035_Y), .A0(D7473_Y));
KC_AOI22_X1 D9034 ( .A1(D6248_Q), .B0(D9054_Y), .B1(D2091_Q),     .Y(D9034_Y), .A0(D9041_Y));
KC_AOI22_X1 D9032 ( .A1(D9158_Y), .B0(D9041_Y), .B1(D9019_Q),     .Y(D9032_Y), .A0(D9068_Y));
KC_AOI22_X1 D9031 ( .A1(D9171_Y), .B0(D308_Y), .B1(D8064_Y),     .Y(D9031_Y), .A0(D9068_Y));
KC_AOI22_X1 D8983 ( .A1(D7315_Y), .B0(D8974_Y), .B1(D2665_Y),     .Y(D8983_Y), .A0(D7_Y));
KC_AOI22_X1 D8982 ( .A1(D8986_Y), .B0(D8895_Q), .B1(D7184_Y),     .Y(D8982_Y), .A0(D2095_Y));
KC_AOI22_X1 D8981 ( .A1(D8986_Y), .B0(D151_Q), .B1(D7184_Y),     .Y(D8981_Y), .A0(D9482_Y));
KC_AOI22_X1 D8979 ( .A1(D7315_Y), .B0(D8974_Y), .B1(D2075_Y),     .Y(D8979_Y), .A0(D305_Q));
KC_AOI22_X1 D8967 ( .A1(D8974_Y), .B0(D7430_Y), .B1(D8962_Y),     .Y(D8967_Y), .A0(D2861_Y));
KC_AOI22_X1 D8966 ( .A1(D8974_Y), .B0(D7430_Y), .B1(D9040_Y),     .Y(D8966_Y), .A0(D9005_Y));
KC_AOI22_X1 D8965 ( .A1(D8974_Y), .B0(D7430_Y), .B1(D52_Y),     .Y(D8965_Y), .A0(D2066_Y));
KC_AOI22_X1 D8961 ( .A1(D7362_Y), .B0(D9475_Y), .B1(D8986_Y),     .Y(D8961_Y), .A0(D9477_Y));
KC_AOI22_X1 D8960 ( .A1(D8917_Y), .B0(D7473_Y), .B1(D8061_Y),     .Y(D8960_Y), .A0(D9475_Y));
KC_AOI22_X1 D8959 ( .A1(D51_Y), .B0(D308_Y), .B1(D8068_Y), .Y(D8959_Y),     .A0(D9041_Y));
KC_AOI22_X1 D8926 ( .A1(D8900_Y), .B0(D273_Y), .B1(D8883_Y),     .Y(D8926_Y), .A0(D8954_Q));
KC_AOI22_X1 D8925 ( .A1(D8900_Y), .B0(D7_Y), .B1(D8883_Y), .Y(D8925_Y),     .A0(D273_Y));
KC_AOI22_X1 D8924 ( .A1(D8900_Y), .B0(D8954_Q), .B1(D8883_Y),     .Y(D8924_Y), .A0(D8824_Q));
KC_AOI22_X1 D8923 ( .A1(D9990_Y), .B0(D57_Y), .B1(D7456_Y),     .Y(D8923_Y), .A0(D273_Y));
KC_AOI22_X1 D8921 ( .A1(D2070_Y), .B0(D7394_Y), .B1(D8945_Y),     .Y(D8921_Y), .A0(D8897_Q));
KC_AOI22_X1 D8920 ( .A1(D7313_Y), .B0(D7394_Y), .B1(D8947_Y),     .Y(D8920_Y), .A0(D2090_Q));
KC_AOI22_X1 D8914 ( .A1(D9990_Y), .B0(D41_Y), .B1(D7456_Y),     .Y(D8914_Y), .A0(D7_Y));
KC_AOI22_X1 D8911 ( .A1(D9990_Y), .B0(D51_Y), .B1(D7456_Y),     .Y(D8911_Y), .A0(D272_Y));
KC_AOI22_X1 D8909 ( .A1(D9990_Y), .B0(D7613_Y), .B1(D7456_Y),     .Y(D8909_Y), .A0(D8954_Q));
KC_AOI22_X1 D8906 ( .A1(D7313_Y), .B0(D7393_Y), .B1(D334_Q),     .Y(D8906_Y), .A0(D273_Y));
KC_AOI22_X1 D8905 ( .A1(D7313_Y), .B0(D7393_Y), .B1(D9019_Q),     .Y(D8905_Y), .A0(D7_Y));
KC_AOI22_X1 D8879 ( .A1(D147_Q), .B0(D8901_Y), .B1(D8825_Q),     .Y(D8879_Y), .A0(D7345_Y));
KC_AOI22_X1 D8878 ( .A1(D9982_Q), .B0(D8901_Y), .B1(D231_Q),     .Y(D8878_Y), .A0(D7345_Y));
KC_AOI22_X1 D8873 ( .A1(D2070_Y), .B0(D7394_Y), .B1(D16794_Y),     .Y(D8873_Y), .A0(D8896_Q));
KC_AOI22_X1 D8872 ( .A1(D8883_Y), .B0(D8897_Q), .B1(D7345_Y),     .Y(D8872_Y), .A0(D8899_Q));
KC_AOI22_X1 D8867 ( .A1(D2070_Y), .B0(D7394_Y), .B1(D8892_Y),     .Y(D8867_Y), .A0(D8895_Q));
KC_AOI22_X1 D8863 ( .A1(D7345_Y), .B0(D2090_Q), .B1(D8883_Y),     .Y(D8863_Y), .A0(D8899_Q));
KC_AOI22_X1 D8858 ( .A1(D8899_Q), .B0(D8865_Y), .B1(D7430_Y),     .Y(D8858_Y), .A0(D9990_Y));
KC_AOI22_X1 D8857 ( .A1(D9990_Y), .B0(D7394_Y), .B1(D16793_Y),     .Y(D8857_Y), .A0(D8824_Q));
KC_AOI22_X1 D8856 ( .A1(D2070_Y), .B0(D7394_Y), .B1(D16792_Y),     .Y(D8856_Y), .A0(D305_Q));
KC_AOI22_X1 D8855 ( .A1(D9990_Y), .B0(D7394_Y), .B1(D1475_Y),     .Y(D8855_Y), .A0(D2090_Q));
KC_AOI22_X1 D8854 ( .A1(D9990_Y), .B0(D7394_Y), .B1(D8890_Y),     .Y(D8854_Y), .A0(D8897_Q));
KC_AOI22_X1 D8852 ( .A1(D2070_Y), .B0(D7394_Y), .B1(D16791_Y),     .Y(D8852_Y), .A0(D8898_Q));
KC_AOI22_X1 D8850 ( .A1(D8901_Y), .B0(D8955_Q), .B1(D8900_Y),     .Y(D8850_Y), .A0(D8896_Q));
KC_AOI22_X1 D8847 ( .A1(D2070_Y), .B0(D7394_Y), .B1(D8891_Y),     .Y(D8847_Y), .A0(D8955_Q));
KC_AOI22_X1 D8846 ( .A1(D8883_Y), .B0(D2090_Q), .B1(D8900_Y),     .Y(D8846_Y), .A0(D8824_Q));
KC_AOI22_X1 D8845 ( .A1(D8900_Y), .B0(D8897_Q), .B1(D8883_Y),     .Y(D8845_Y), .A0(D8898_Q));
KC_AOI22_X1 D8765 ( .A1(D8784_Y), .B0(D8763_Y), .B1(D8766_Y),     .Y(D8765_Y), .A0(D8746_Y));
KC_AOI22_X1 D8734 ( .A1(D8772_Y), .B0(D8812_Y), .B1(D8741_Y),     .Y(D8734_Y), .A0(D9480_Y));
KC_AOI22_X1 D8649 ( .A1(D2170_Y), .B0(D9876_Q), .B1(D10560_Y),     .Y(D8649_Y), .A0(D9908_Q));
KC_AOI22_X1 D8648 ( .A1(D6915_Y), .B0(D8658_Q), .B1(D6973_Y),     .Y(D8648_Y), .A0(D1353_Q));
KC_AOI22_X1 D8647 ( .A1(D6915_Y), .B0(D8657_Q), .B1(D6973_Y),     .Y(D8647_Y), .A0(D8651_Q));
KC_AOI22_X1 D8646 ( .A1(D6915_Y), .B0(D8655_Q), .B1(D6973_Y),     .Y(D8646_Y), .A0(D8650_Q));
KC_AOI22_X1 D8645 ( .A1(D8651_Q), .B0(D5542_Y), .B1(D8657_Q),     .Y(D8645_Y), .A0(D5543_Y));
KC_AOI22_X1 D8644 ( .A1(D8650_Q), .B0(D5542_Y), .B1(D8655_Q),     .Y(D8644_Y), .A0(D5543_Y));
KC_AOI22_X1 D8625 ( .A1(D7022_Y), .B0(D8344_Y), .B1(D10583_Y),     .Y(D8625_Y), .A0(D8346_Y));
KC_AOI22_X1 D8624 ( .A1(D7032_Y), .B0(D8344_Y), .B1(D10590_Y),     .Y(D8624_Y), .A0(D8346_Y));
KC_AOI22_X1 D8623 ( .A1(D1144_Y), .B0(D8639_Q), .B1(D10535_Y),     .Y(D8623_Y), .A0(D1296_Q));
KC_AOI22_X1 D8622 ( .A1(D1144_Y), .B0(D8640_Q), .B1(D10535_Y),     .Y(D8622_Y), .A0(D8643_Q));
KC_AOI22_X1 D8621 ( .A1(D7027_Y), .B0(D8344_Y), .B1(D10584_Y),     .Y(D8621_Y), .A0(D8346_Y));
KC_AOI22_X1 D8620 ( .A1(D1682_Y), .B0(D8641_Q), .B1(D6991_Y),     .Y(D8620_Y), .A0(D8634_Q));
KC_AOI22_X1 D8619 ( .A1(D5584_Y), .B0(D8344_Y), .B1(D9893_Y),     .Y(D8619_Y), .A0(D8346_Y));
KC_AOI22_X1 D8618 ( .A1(D8635_Q), .B0(D11011_Y), .B1(D8632_Q),     .Y(D8618_Y), .A0(D11010_Y));
KC_AOI22_X1 D8617 ( .A1(D1682_Y), .B0(D8638_Q), .B1(D6991_Y),     .Y(D8617_Y), .A0(D8636_Q));
KC_AOI22_X1 D8616 ( .A1(D8636_Q), .B0(D5497_Y), .B1(D8638_Q),     .Y(D8616_Y), .A0(D1082_Y));
KC_AOI22_X1 D8615 ( .A1(D5582_Y), .B0(D8344_Y), .B1(D9894_Y),     .Y(D8615_Y), .A0(D8346_Y));
KC_AOI22_X1 D8614 ( .A1(D5578_Y), .B0(D8344_Y), .B1(D9862_Y),     .Y(D8614_Y), .A0(D8346_Y));
KC_AOI22_X1 D8613 ( .A1(D8610_Y), .B0(D8344_Y), .B1(D10568_Y),     .Y(D8613_Y), .A0(D8346_Y));
KC_AOI22_X1 D8612 ( .A1(D1682_Y), .B0(D8633_Q), .B1(D6991_Y),     .Y(D8612_Y), .A0(D8630_Q));
KC_AOI22_X1 D8611 ( .A1(D8630_Q), .B0(D5497_Y), .B1(D8633_Q),     .Y(D8611_Y), .A0(D1082_Y));
KC_AOI22_X1 D8562 ( .A1(D5547_Y), .B0(D1927_Q), .B1(D7001_Y),     .Y(D8562_Y), .A0(D2032_Y));
KC_AOI22_X1 D8560 ( .A1(D12004_Y), .B0(D8594_Q), .B1(D1186_Y),     .Y(D8560_Y), .A0(D2032_Y));
KC_AOI22_X1 D8556 ( .A1(D5546_Y), .B0(D8344_Y), .B1(D9810_Y),     .Y(D8556_Y), .A0(D8346_Y));
KC_AOI22_X1 D8555 ( .A1(D6981_Y), .B0(D8344_Y), .B1(D9809_Y),     .Y(D8555_Y), .A0(D8346_Y));
KC_AOI22_X1 D8554 ( .A1(D1680_Y), .B0(D8344_Y), .B1(D10522_Y),     .Y(D8554_Y), .A0(D8346_Y));
KC_AOI22_X1 D8553 ( .A1(D8609_Y), .B0(D8344_Y), .B1(D9811_Y),     .Y(D8553_Y), .A0(D8346_Y));
KC_AOI22_X1 D8469 ( .A1(D8432_Y), .B0(D5496_Y), .B1(D2032_Y),     .Y(D8469_Y), .A0(D11390_Q));
KC_AOI22_X1 D8416 ( .A1(D5418_Y), .B0(D8345_Y), .B1(D10399_Y),     .Y(D8416_Y), .A0(D8278_Y));
KC_AOI22_X1 D8408 ( .A1(D5446_Y), .B0(D8345_Y), .B1(D9666_Y),     .Y(D8408_Y), .A0(D8278_Y));
KC_AOI22_X1 D8407 ( .A1(D3924_Y), .B0(D8345_Y), .B1(D9670_Y),     .Y(D8407_Y), .A0(D8278_Y));
KC_AOI22_X1 D8396 ( .A1(D3915_Y), .B0(D8345_Y), .B1(D9678_Y),     .Y(D8396_Y), .A0(D8278_Y));
KC_AOI22_X1 D8389 ( .A1(D5435_Y), .B0(D8345_Y), .B1(D10385_Y),     .Y(D8389_Y), .A0(D8278_Y));
KC_AOI22_X1 D8379 ( .A1(D5430_Y), .B0(D8345_Y), .B1(D9668_Y),     .Y(D8379_Y), .A0(D8278_Y));
KC_AOI22_X1 D8374 ( .A1(D3906_Y), .B0(D8345_Y), .B1(D10383_Y),     .Y(D8374_Y), .A0(D8278_Y));
KC_AOI22_X1 D8373 ( .A1(D1553_Y), .B0(D8345_Y), .B1(D10402_Y),     .Y(D8373_Y), .A0(D8278_Y));
KC_AOI22_X1 D8349 ( .A1(D1552_Y), .B0(D6744_Q), .B1(D91_Y),     .Y(D8349_Y), .A0(D6759_Y));
KC_AOI22_X1 D8347 ( .A1(D737_Y), .B0(D8345_Y), .B1(D10841_Y),     .Y(D8347_Y), .A0(D8278_Y));
KC_AOI22_X1 D8285 ( .A1(D5429_Y), .B0(D6826_Q), .B1(D8301_Y),     .Y(D8285_Y), .A0(D6759_Y));
KC_AOI22_X1 D8284 ( .A1(D8298_Y), .B0(D6759_Y), .B1(D5339_Y),     .Y(D8284_Y), .A0(D8463_Q));
KC_AOI22_X1 D8276 ( .A1(D3903_Y), .B0(D6829_Q), .B1(D8299_Y),     .Y(D8276_Y), .A0(D6759_Y));
KC_AOI22_X1 D8271 ( .A1(D5365_Y), .B0(D8345_Y), .B1(D10845_Y),     .Y(D8271_Y), .A0(D8278_Y));
KC_AOI22_X1 D8268 ( .A1(D3830_Y), .B0(D8345_Y), .B1(D10839_Y),     .Y(D8268_Y), .A0(D8278_Y));
KC_AOI22_X1 D8200 ( .A1(D11139_Y), .B0(D8339_Y), .B1(D6570_Y),     .Y(D8200_Y), .A0(D8337_Y));
KC_AOI22_X1 D8197 ( .A1(D740_Y), .B0(D796_Q), .B1(D8216_Y),     .Y(D8197_Y), .A0(D6759_Y));
KC_AOI22_X1 D8196 ( .A1(D3792_Y), .B0(D789_Q), .B1(D8218_Y),     .Y(D8196_Y), .A0(D8211_Y));
KC_AOI22_X1 D8195 ( .A1(D11682_Y), .B0(D8339_Y), .B1(D6624_Y),     .Y(D8195_Y), .A0(D8337_Y));
KC_AOI22_X1 D8189 ( .A1(D8199_Y), .B0(D8184_Y), .B1(D5288_Y),     .Y(D8189_Y), .A0(D8198_Y));
KC_AOI22_X1 D8188 ( .A1(D11217_Y), .B0(D8339_Y), .B1(D6619_Y),     .Y(D8188_Y), .A0(D8337_Y));
KC_AOI22_X1 D8180 ( .A1(D3829_Y), .B0(D8238_Q), .B1(D8214_Y),     .Y(D8180_Y), .A0(D6759_Y));
KC_AOI22_X1 D8176 ( .A1(D8199_Y), .B0(D8184_Y), .B1(D6709_Y),     .Y(D8176_Y), .A0(D8182_Y));
KC_AOI22_X1 D8173 ( .A1(D8199_Y), .B0(D8184_Y), .B1(D3776_Y),     .Y(D8173_Y), .A0(D8181_Y));
KC_AOI22_X1 D8168 ( .A1(D6759_Y), .B0(D785_Q), .B1(D8209_Y),     .Y(D8168_Y), .A0(D3776_Y));
KC_AOI22_X1 D8119 ( .A1(D5174_Y), .B0(D672_Q), .B1(D8127_Y),     .Y(D8119_Y), .A0(D8211_Y));
KC_AOI22_X1 D8118 ( .A1(D11709_Y), .B0(D8339_Y), .B1(D6634_Y),     .Y(D8118_Y), .A0(D8337_Y));
KC_AOI22_X1 D8113 ( .A1(D11704_Y), .B0(D8339_Y), .B1(D1557_Y),     .Y(D8113_Y), .A0(D8337_Y));
KC_AOI22_X1 D8112 ( .A1(D10698_Y), .B0(D8339_Y), .B1(D6576_Y),     .Y(D8112_Y), .A0(D8337_Y));
KC_AOI22_X1 D8104 ( .A1(D10697_Y), .B0(D8339_Y), .B1(D5155_Y),     .Y(D8104_Y), .A0(D8337_Y));
KC_AOI22_X1 D8103 ( .A1(D10200_Y), .B0(D8339_Y), .B1(D5171_Y),     .Y(D8103_Y), .A0(D8337_Y));
KC_AOI22_X1 D8100 ( .A1(D8135_Y), .B0(D8120_Y), .B1(D8835_Q),     .Y(D8100_Y), .A0(D7655_Y));
KC_AOI22_X1 D8097 ( .A1(D11140_Y), .B0(D8339_Y), .B1(D5173_Y),     .Y(D8097_Y), .A0(D8337_Y));
KC_AOI22_X1 D8096 ( .A1(D10691_Y), .B0(D8339_Y), .B1(D6584_Y),     .Y(D8096_Y), .A0(D8337_Y));
KC_AOI22_X1 D8080 ( .A1(D8148_Q), .B0(D8120_Y), .B1(D7475_Q),     .Y(D8080_Y), .A0(D8221_Y));
KC_AOI22_X1 D8075 ( .A1(D10756_Y), .B0(D8339_Y), .B1(D5166_Y),     .Y(D8075_Y), .A0(D8337_Y));
KC_AOI22_X1 D8074 ( .A1(D10676_Y), .B0(D8339_Y), .B1(D5159_Y),     .Y(D8074_Y), .A0(D8337_Y));
KC_AOI22_X1 D8012 ( .A1(D6585_Y), .B0(D8052_Q), .B1(D8026_Y),     .Y(D8012_Y), .A0(D8211_Y));
KC_AOI22_X1 D8010 ( .A1(D8211_Y), .B0(D8053_Q), .B1(D8024_Y),     .Y(D8010_Y), .A0(D5288_Y));
KC_AOI22_X1 D8004 ( .A1(D5180_Y), .B0(D669_Q), .B1(D8028_Y),     .Y(D8004_Y), .A0(D8211_Y));
KC_AOI22_X1 D7996 ( .A1(D8027_Y), .B0(D8211_Y), .B1(D5160_Y),     .Y(D7996_Y), .A0(D8055_Q));
KC_AOI22_X1 D7995 ( .A1(D8211_Y), .B0(D8054_Q), .B1(D8025_Y),     .Y(D7995_Y), .A0(D6580_Y));
KC_AOI22_X1 D7930 ( .A1(D7916_Y), .B0(D7963_Y), .B1(D7925_Y),     .Y(D7930_Y), .A0(D524_Q));
KC_AOI22_X1 D7906 ( .A1(D7916_Y), .B0(D727_Y), .B1(D7921_Y),     .Y(D7906_Y), .A0(D8466_Y));
KC_AOI22_X1 D7693 ( .A1(D7621_Y), .B0(D7733_Q), .B1(D2099_Y),     .Y(D7693_Y), .A0(D7499_Y));
KC_AOI22_X1 D7674 ( .A1(D7703_Y), .B0(D7740_Y), .B1(D7740_Y),     .Y(D7674_Y), .A0(D404_Y));
KC_AOI22_X1 D7619 ( .A1(D2099_Y), .B0(D9102_Y), .B1(D7621_Y),     .Y(D7619_Y), .A0(D7732_Q));
KC_AOI22_X1 D7568 ( .A1(D21_Y), .B0(D1870_Y), .B1(D6191_Y),     .Y(D7568_Y), .A0(D13287_Y));
KC_AOI22_X1 D7566 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D7595_Y),     .Y(D7566_Y), .A0(D724_Y));
KC_AOI22_X1 D7560 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D7599_Y),     .Y(D7560_Y), .A0(D13288_Y));
KC_AOI22_X1 D7552 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D7666_Y),     .Y(D7552_Y), .A0(D12764_Y));
KC_AOI22_X1 D7551 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D7592_Y),     .Y(D7551_Y), .A0(D12762_Y));
KC_AOI22_X1 D7546 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D358_Y),     .Y(D7546_Y), .A0(D725_Y));
KC_AOI22_X1 D7542 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D1949_Y),     .Y(D7542_Y), .A0(D13285_Y));
KC_AOI22_X1 D7540 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D1804_Y),     .Y(D7540_Y), .A0(D12761_Y));
KC_AOI22_X1 D7539 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D6188_Y),     .Y(D7539_Y), .A0(D12863_Y));
KC_AOI22_X1 D7498 ( .A1(D7503_Y), .B0(D6075_Y), .B1(D20_Y),     .Y(D7498_Y), .A0(D9147_Y));
KC_AOI22_X1 D7495 ( .A1(D1869_Y), .B0(D1870_Y), .B1(D7604_Y),     .Y(D7495_Y), .A0(D12763_Y));
KC_AOI22_X1 D7493 ( .A1(D1864_Y), .B0(D7494_Y), .B1(D7534_Q),     .Y(D7493_Y), .A0(D60_Q));
KC_AOI22_X1 D7492 ( .A1(D7362_Y), .B0(D7476_Q), .B1(D7494_Y),     .Y(D7492_Y), .A0(D9475_Y));
KC_AOI22_X1 D7420 ( .A1(D5966_Y), .B0(D9147_Y), .B1(D8908_Y),     .Y(D7420_Y), .A0(D6022_Y));
KC_AOI22_X1 D7346 ( .A1(D7538_Y), .B0(D7333_Y), .B1(D7500_Y),     .Y(D7346_Y), .A0(D7233_Y));
KC_AOI22_X1 D7339 ( .A1(D7390_Y), .B0(D1877_Y), .B1(D7410_Y),     .Y(D7339_Y), .A0(D7170_Y));
KC_AOI22_X1 D7332 ( .A1(D4444_Y), .B0(D7443_Y), .B1(D7333_Y),     .Y(D7332_Y), .A0(D247_Y));
KC_AOI22_X1 D7311 ( .A1(D4444_Y), .B0(D9479_Y), .B1(D7342_Y),     .Y(D7311_Y), .A0(D5863_Y));
KC_AOI22_X1 D7221 ( .A1(D2095_Y), .B0(D7234_Y), .B1(D7169_Y),     .Y(D7221_Y), .A0(D7193_Y));
KC_AOI22_X1 D7073 ( .A1(D6972_Y), .B0(D8654_Q), .B1(D6974_Y),     .Y(D7073_Y), .A0(D1350_Q));
KC_AOI22_X1 D7072 ( .A1(D7078_Q), .B0(D5509_Y), .B1(D7081_Q),     .Y(D7072_Y), .A0(D5540_Y));
KC_AOI22_X1 D7071 ( .A1(D1353_Q), .B0(D5542_Y), .B1(D8658_Q),     .Y(D7071_Y), .A0(D5543_Y));
KC_AOI22_X1 D7070 ( .A1(D7083_Q), .B0(D5509_Y), .B1(D8653_Q),     .Y(D7070_Y), .A0(D5540_Y));
KC_AOI22_X1 D7069 ( .A1(D7042_Q), .B0(D5498_Y), .B1(D7043_Q),     .Y(D7069_Y), .A0(D1596_Y));
KC_AOI22_X1 D7067 ( .A1(D6972_Y), .B0(D8653_Q), .B1(D6974_Y),     .Y(D7067_Y), .A0(D7083_Q));
KC_AOI22_X1 D7066 ( .A1(D7077_Q), .B0(D5509_Y), .B1(D8652_Q),     .Y(D7066_Y), .A0(D5540_Y));
KC_AOI22_X1 D7065 ( .A1(D1350_Q), .B0(D5509_Y), .B1(D8654_Q),     .Y(D7065_Y), .A0(D5540_Y));
KC_AOI22_X1 D7064 ( .A1(D1352_Q), .B0(D5498_Y), .B1(D7079_Q),     .Y(D7064_Y), .A0(D1596_Y));
KC_AOI22_X1 D7063 ( .A1(D6915_Y), .B0(D7056_Q), .B1(D6973_Y),     .Y(D7063_Y), .A0(D7054_Q));
KC_AOI22_X1 D7041 ( .A1(D7054_Q), .B0(D5542_Y), .B1(D7056_Q),     .Y(D7041_Y), .A0(D5543_Y));
KC_AOI22_X1 D7040 ( .A1(D1682_Y), .B0(D1933_Q), .B1(D6991_Y),     .Y(D7040_Y), .A0(D121_Q));
KC_AOI22_X1 D7038 ( .A1(D1298_Q), .B0(D5542_Y), .B1(D1300_Q),     .Y(D7038_Y), .A0(D5543_Y));
KC_AOI22_X1 D7037 ( .A1(D121_Q), .B0(D5497_Y), .B1(D1933_Q),     .Y(D7037_Y), .A0(D1082_Y));
KC_AOI22_X1 D7036 ( .A1(D6915_Y), .B0(D1300_Q), .B1(D6973_Y),     .Y(D7036_Y), .A0(D1298_Q));
KC_AOI22_X1 D7035 ( .A1(D5522_Y), .B0(D7051_Q), .B1(D6921_Y),     .Y(D7035_Y), .A0(D7047_Q));
KC_AOI22_X1 D7034 ( .A1(D6972_Y), .B0(D7048_Q), .B1(D6974_Y),     .Y(D7034_Y), .A0(D7046_Q));
KC_AOI22_X1 D7033 ( .A1(D1682_Y), .B0(D8642_Q), .B1(D6991_Y),     .Y(D7033_Y), .A0(D1295_Q));
KC_AOI22_X1 D7031 ( .A1(D7046_Q), .B0(D5509_Y), .B1(D7048_Q),     .Y(D7031_Y), .A0(D5540_Y));
KC_AOI22_X1 D7030 ( .A1(D1295_Q), .B0(D5497_Y), .B1(D8642_Q),     .Y(D7030_Y), .A0(D1082_Y));
KC_AOI22_X1 D7029 ( .A1(D7047_Q), .B0(D5498_Y), .B1(D7051_Q),     .Y(D7029_Y), .A0(D1596_Y));
KC_AOI22_X1 D7028 ( .A1(D6915_Y), .B0(D8631_Q), .B1(D6973_Y),     .Y(D7028_Y), .A0(D1356_Q));
KC_AOI22_X1 D7025 ( .A1(D1356_Q), .B0(D5542_Y), .B1(D8631_Q),     .Y(D7025_Y), .A0(D5543_Y));
KC_AOI22_X1 D7024 ( .A1(D7085_Q), .B0(D5498_Y), .B1(D7082_Q),     .Y(D7024_Y), .A0(D1596_Y));
KC_AOI22_X1 D7023 ( .A1(D6972_Y), .B0(D8652_Q), .B1(D6974_Y),     .Y(D7023_Y), .A0(D7077_Q));
KC_AOI22_X1 D7020 ( .A1(D6972_Y), .B0(D7081_Q), .B1(D6974_Y),     .Y(D7020_Y), .A0(D7078_Q));
KC_AOI22_X1 D7017 ( .A1(D7026_Y), .B0(D7008_Q), .B1(D6998_Y),     .Y(D7017_Y), .A0(D2032_Y));
KC_AOI22_X1 D6990 ( .A1(D6985_Y), .B0(D1774_Q), .B1(D7000_Y),     .Y(D6990_Y), .A0(D2032_Y));
KC_AOI22_X1 D6988 ( .A1(D1682_Y), .B0(D7007_Q), .B1(D6991_Y),     .Y(D6988_Y), .A0(D7006_Q));
KC_AOI22_X1 D6987 ( .A1(D2032_Y), .B0(D7005_Q), .B1(D6997_Y),     .Y(D6987_Y), .A0(D7068_Y));
KC_AOI22_X1 D6984 ( .A1(D6972_Y), .B0(D7004_Q), .B1(D6974_Y),     .Y(D6984_Y), .A0(D1211_Q));
KC_AOI22_X1 D6983 ( .A1(D7011_Q), .B0(D5497_Y), .B1(D7013_Q),     .Y(D6983_Y), .A0(D1082_Y));
KC_AOI22_X1 D6982 ( .A1(D6972_Y), .B0(D7012_Q), .B1(D6974_Y),     .Y(D6982_Y), .A0(D7014_Q));
KC_AOI22_X1 D6980 ( .A1(D6915_Y), .B0(D1784_Q), .B1(D6973_Y),     .Y(D6980_Y), .A0(D1783_Q));
KC_AOI22_X1 D6979 ( .A1(D1682_Y), .B0(D7013_Q), .B1(D6991_Y),     .Y(D6979_Y), .A0(D7011_Q));
KC_AOI22_X1 D6978 ( .A1(D7014_Q), .B0(D5509_Y), .B1(D7012_Q),     .Y(D6978_Y), .A0(D5540_Y));
KC_AOI22_X1 D6933 ( .A1(D2032_Y), .B0(D1126_Q), .B1(D6945_Y),     .Y(D6933_Y), .A0(D5501_Y));
KC_AOI22_X1 D6932 ( .A1(D1743_Y), .B0(D6930_Y), .B1(D5501_Y),     .Y(D6932_Y), .A0(D6928_Y));
KC_AOI22_X1 D6917 ( .A1(D6938_Y), .B0(D6919_Y), .B1(D7068_Y),     .Y(D6917_Y), .A0(D1683_Y));
KC_AOI22_X1 D6914 ( .A1(D2032_Y), .B0(D6970_Q), .B1(D6999_Y),     .Y(D6914_Y), .A0(D5599_Y));
KC_AOI22_X1 D6913 ( .A1(D6938_Y), .B0(D6919_Y), .B1(D5599_Y),     .Y(D6913_Y), .A0(D1684_Y));
KC_AOI22_X1 D6876 ( .A1(D6824_Q), .B0(D5440_Y), .B1(D6823_Q),     .Y(D6876_Y), .A0(D1628_Y));
KC_AOI22_X1 D6875 ( .A1(D976_Y), .B0(D903_Q), .B1(D993_Y), .Y(D6875_Y),     .A0(D6759_Y));
KC_AOI22_X1 D6874 ( .A1(D6818_Q), .B0(D6822_Q), .B1(D5440_Y),     .Y(D6874_Y), .A0(D1628_Y));
KC_AOI22_X1 D6870 ( .A1(D3916_Y), .B0(D1779_Q), .B1(D6884_Y),     .Y(D6870_Y), .A0(D6759_Y));
KC_AOI22_X1 D6865 ( .A1(D6853_Y), .B0(D6901_Q), .B1(D6869_Y),     .Y(D6865_Y), .A0(D6902_Q));
KC_AOI22_X1 D6858 ( .A1(D6897_Q), .B0(D972_Y), .B1(D6898_Q),     .Y(D6858_Y), .A0(D6862_Y));
KC_AOI22_X1 D6857 ( .A1(D6899_Q), .B0(D972_Y), .B1(D6895_Q),     .Y(D6857_Y), .A0(D6862_Y));
KC_AOI22_X1 D6852 ( .A1(D6853_Y), .B0(D6898_Q), .B1(D6869_Y),     .Y(D6852_Y), .A0(D6897_Q));
KC_AOI22_X1 D6851 ( .A1(D6862_Y), .B0(D6912_Q), .B1(D972_Y),     .Y(D6851_Y), .A0(D6911_Q));
KC_AOI22_X1 D6850 ( .A1(D6853_Y), .B0(D6895_Q), .B1(D6869_Y),     .Y(D6850_Y), .A0(D6899_Q));
KC_AOI22_X1 D6849 ( .A1(D6853_Y), .B0(D6912_Q), .B1(D6869_Y),     .Y(D6849_Y), .A0(D6911_Q));
KC_AOI22_X1 D6846 ( .A1(D6863_Y), .B0(D6896_Q), .B1(D6860_Y),     .Y(D6846_Y), .A0(D6893_Q));
KC_AOI22_X1 D6845 ( .A1(D5436_Y), .B0(D6896_Q), .B1(D973_Y),     .Y(D6845_Y), .A0(D6893_Q));
KC_AOI22_X1 D6844 ( .A1(D6878_Y), .B0(D1775_Q), .B1(D6861_Y),     .Y(D6844_Y), .A0(D1012_Q));
KC_AOI22_X1 D6841 ( .A1(D6863_Y), .B0(D6892_Q), .B1(D6860_Y),     .Y(D6841_Y), .A0(D1776_Q));
KC_AOI22_X1 D6840 ( .A1(D6966_Q), .B0(D973_Y), .B1(D6894_Q),     .Y(D6840_Y), .A0(D5436_Y));
KC_AOI22_X1 D6839 ( .A1(D1776_Q), .B0(D973_Y), .B1(D6892_Q),     .Y(D6839_Y), .A0(D5436_Y));
KC_AOI22_X1 D6838 ( .A1(D6878_Y), .B0(D6968_Q), .B1(D6861_Y),     .Y(D6838_Y), .A0(D6964_Q));
KC_AOI22_X1 D6837 ( .A1(D6878_Y), .B0(D5465_Q), .B1(D6861_Y),     .Y(D6837_Y), .A0(D117_Q));
KC_AOI22_X1 D6835 ( .A1(D6863_Y), .B0(D6894_Q), .B1(D6860_Y),     .Y(D6835_Y), .A0(D6966_Q));
KC_AOI22_X1 D6834 ( .A1(D6863_Y), .B0(D1777_Q), .B1(D6860_Y),     .Y(D6834_Y), .A0(D6969_Q));
KC_AOI22_X1 D6770 ( .A1(D6866_Y), .B0(D8339_Y), .B1(D6688_Y),     .Y(D6770_Y), .A0(D1920_Y));
KC_AOI22_X1 D6769 ( .A1(D6871_Y), .B0(D8339_Y), .B1(D6707_Y),     .Y(D6769_Y), .A0(D1920_Y));
KC_AOI22_X1 D6763 ( .A1(D5461_Y), .B0(D6822_Q), .B1(D6868_Y),     .Y(D6763_Y), .A0(D6818_Q));
KC_AOI22_X1 D6762 ( .A1(D6872_Y), .B0(D8339_Y), .B1(D6717_Y),     .Y(D6762_Y), .A0(D1920_Y));
KC_AOI22_X1 D6761 ( .A1(D6867_Y), .B0(D8339_Y), .B1(D6694_Y),     .Y(D6761_Y), .A0(D1920_Y));
KC_AOI22_X1 D6724 ( .A1(D6655_Q), .B0(D5266_Y), .B1(D6756_Q),     .Y(D6724_Y), .A0(D6695_Y));
KC_AOI22_X1 D6723 ( .A1(D6656_Q), .B0(D6760_Y), .B1(D6757_Q),     .Y(D6723_Y), .A0(D831_Y));
KC_AOI22_X1 D6722 ( .A1(D1689_Y), .B0(D6756_Q), .B1(D1688_Y),     .Y(D6722_Y), .A0(D6655_Q));
KC_AOI22_X1 D6721 ( .A1(D795_Q), .B0(D6689_Y), .B1(D6657_Q),     .Y(D6721_Y), .A0(D5322_Y));
KC_AOI22_X1 D6716 ( .A1(D5408_Y), .B0(D6657_Q), .B1(D1555_Y),     .Y(D6716_Y), .A0(D795_Q));
KC_AOI22_X1 D6715 ( .A1(D1801_Y), .B0(D6757_Q), .B1(D157_Y),     .Y(D6715_Y), .A0(D6656_Q));
KC_AOI22_X1 D6714 ( .A1(D1801_Y), .B0(D6752_Q), .B1(D157_Y),     .Y(D6714_Y), .A0(D6755_Q));
KC_AOI22_X1 D6712 ( .A1(D831_Y), .B0(D6752_Q), .B1(D6760_Y),     .Y(D6712_Y), .A0(D6755_Q));
KC_AOI22_X1 D6708 ( .A1(D5322_Y), .B0(D6753_Q), .B1(D6689_Y),     .Y(D6708_Y), .A0(D793_Q));
KC_AOI22_X1 D6706 ( .A1(D6759_Y), .B0(D6750_Q), .B1(D8213_Y),     .Y(D6706_Y), .A0(D6618_Y));
KC_AOI22_X1 D6705 ( .A1(D1689_Y), .B0(D6749_Q), .B1(D1688_Y),     .Y(D6705_Y), .A0(D6751_Q));
KC_AOI22_X1 D6704 ( .A1(D6695_Y), .B0(D6749_Q), .B1(D5266_Y),     .Y(D6704_Y), .A0(D6751_Q));
KC_AOI22_X1 D6703 ( .A1(D5408_Y), .B0(D6753_Q), .B1(D1555_Y),     .Y(D6703_Y), .A0(D793_Q));
KC_AOI22_X1 D6701 ( .A1(D6747_Q), .B0(D5266_Y), .B1(D6748_Q),     .Y(D6701_Y), .A0(D6695_Y));
KC_AOI22_X1 D6700 ( .A1(D1689_Y), .B0(D6748_Q), .B1(D1688_Y),     .Y(D6700_Y), .A0(D6747_Q));
KC_AOI22_X1 D6699 ( .A1(D8199_Y), .B0(D8184_Y), .B1(D6693_Y),     .Y(D6699_Y), .A0(D733_Y));
KC_AOI22_X1 D6697 ( .A1(D907_Q), .B0(D6689_Y), .B1(D1781_Q),     .Y(D6697_Y), .A0(D5322_Y));
KC_AOI22_X1 D6696 ( .A1(D6745_Q), .B0(D5266_Y), .B1(D6746_Q),     .Y(D6696_Y), .A0(D6695_Y));
KC_AOI22_X1 D6692 ( .A1(D6830_Q), .B0(D6689_Y), .B1(D6827_Q),     .Y(D6692_Y), .A0(D5322_Y));
KC_AOI22_X1 D6691 ( .A1(D1689_Y), .B0(D6746_Q), .B1(D1688_Y),     .Y(D6691_Y), .A0(D6745_Q));
KC_AOI22_X1 D6690 ( .A1(D1780_Q), .B0(D6760_Y), .B1(D6743_Q),     .Y(D6690_Y), .A0(D831_Y));
KC_AOI22_X1 D6687 ( .A1(D6828_Q), .B0(D6760_Y), .B1(D1782_Q),     .Y(D6687_Y), .A0(D831_Y));
KC_AOI22_X1 D6686 ( .A1(D5408_Y), .B0(D1781_Q), .B1(D1555_Y),     .Y(D6686_Y), .A0(D907_Q));
KC_AOI22_X1 D6685 ( .A1(D5408_Y), .B0(D6827_Q), .B1(D1555_Y),     .Y(D6685_Y), .A0(D6830_Q));
KC_AOI22_X1 D6684 ( .A1(D1801_Y), .B0(D1782_Q), .B1(D157_Y),     .Y(D6684_Y), .A0(D6828_Q));
KC_AOI22_X1 D6683 ( .A1(D1801_Y), .B0(D6743_Q), .B1(D157_Y),     .Y(D6683_Y), .A0(D1780_Q));
KC_AOI22_X1 D6641 ( .A1(D1689_Y), .B0(D6675_Q), .B1(D1688_Y),     .Y(D6641_Y), .A0(D6667_Q));
KC_AOI22_X1 D6640 ( .A1(D1689_Y), .B0(D673_Q), .B1(D1688_Y),     .Y(D6640_Y), .A0(D6666_Q));
KC_AOI22_X1 D6639 ( .A1(D6666_Q), .B0(D5266_Y), .B1(D673_Q),     .Y(D6639_Y), .A0(D6695_Y));
KC_AOI22_X1 D6638 ( .A1(D6667_Q), .B0(D5266_Y), .B1(D6675_Q),     .Y(D6638_Y), .A0(D6695_Y));
KC_AOI22_X1 D6636 ( .A1(D6663_Q), .B0(D6760_Y), .B1(D6662_Q),     .Y(D6636_Y), .A0(D831_Y));
KC_AOI22_X1 D6635 ( .A1(D1801_Y), .B0(D6662_Q), .B1(D157_Y),     .Y(D6635_Y), .A0(D6663_Q));
KC_AOI22_X1 D6632 ( .A1(D6672_Q), .B0(D5266_Y), .B1(D6673_Q),     .Y(D6632_Y), .A0(D6695_Y));
KC_AOI22_X1 D6631 ( .A1(D1689_Y), .B0(D6673_Q), .B1(D1688_Y),     .Y(D6631_Y), .A0(D6672_Q));
KC_AOI22_X1 D6630 ( .A1(D671_Q), .B0(D6689_Y), .B1(D6674_Q),     .Y(D6630_Y), .A0(D5322_Y));
KC_AOI22_X1 D6629 ( .A1(D6652_Q), .B0(D6760_Y), .B1(D6671_Q),     .Y(D6629_Y), .A0(D831_Y));
KC_AOI22_X1 D6628 ( .A1(D5408_Y), .B0(D6674_Q), .B1(D1555_Y),     .Y(D6628_Y), .A0(D671_Q));
KC_AOI22_X1 D6627 ( .A1(D1801_Y), .B0(D6671_Q), .B1(D157_Y),     .Y(D6627_Y), .A0(D6652_Q));
KC_AOI22_X1 D6626 ( .A1(D6668_Q), .B0(D6760_Y), .B1(D6669_Q),     .Y(D6626_Y), .A0(D831_Y));
KC_AOI22_X1 D6623 ( .A1(D670_Q), .B0(D6689_Y), .B1(D6670_Q),     .Y(D6623_Y), .A0(D5322_Y));
KC_AOI22_X1 D6622 ( .A1(D5408_Y), .B0(D6670_Q), .B1(D1555_Y),     .Y(D6622_Y), .A0(D670_Q));
KC_AOI22_X1 D6621 ( .A1(D6658_Q), .B0(D5266_Y), .B1(D6660_Q),     .Y(D6621_Y), .A0(D6695_Y));
KC_AOI22_X1 D6620 ( .A1(D1689_Y), .B0(D6660_Q), .B1(D1688_Y),     .Y(D6620_Y), .A0(D6658_Q));
KC_AOI22_X1 D6590 ( .A1(D1801_Y), .B0(D6608_Q), .B1(D157_Y),     .Y(D6590_Y), .A0(D6609_Q));
KC_AOI22_X1 D6588 ( .A1(D6611_Q), .B0(D6689_Y), .B1(D6612_Q),     .Y(D6588_Y), .A0(D5322_Y));
KC_AOI22_X1 D6587 ( .A1(D6609_Q), .B0(D6760_Y), .B1(D6608_Q),     .Y(D6587_Y), .A0(D831_Y));
KC_AOI22_X1 D6586 ( .A1(D591_Q), .B0(D6689_Y), .B1(D6596_Q),     .Y(D6586_Y), .A0(D5322_Y));
KC_AOI22_X1 D6583 ( .A1(D6607_Q), .B0(D6760_Y), .B1(D6599_Q),     .Y(D6583_Y), .A0(D831_Y));
KC_AOI22_X1 D6582 ( .A1(D1689_Y), .B0(D6610_Q), .B1(D1688_Y),     .Y(D6582_Y), .A0(D6597_Q));
KC_AOI22_X1 D6581 ( .A1(D6597_Q), .B0(D5266_Y), .B1(D6610_Q),     .Y(D6581_Y), .A0(D6695_Y));
KC_AOI22_X1 D6579 ( .A1(D6604_Q), .B0(D5266_Y), .B1(D6595_Q),     .Y(D6579_Y), .A0(D6695_Y));
KC_AOI22_X1 D6578 ( .A1(D5408_Y), .B0(D6603_Q), .B1(D1555_Y),     .Y(D6578_Y), .A0(D6601_Q));
KC_AOI22_X1 D6577 ( .A1(D6601_Q), .B0(D6689_Y), .B1(D6603_Q),     .Y(D6577_Y), .A0(D5322_Y));
KC_AOI22_X1 D6575 ( .A1(D1801_Y), .B0(D6594_Q), .B1(D157_Y),     .Y(D6575_Y), .A0(D6605_Q));
KC_AOI22_X1 D6574 ( .A1(D1689_Y), .B0(D6595_Q), .B1(D1688_Y),     .Y(D6574_Y), .A0(D6604_Q));
KC_AOI22_X1 D6573 ( .A1(D6605_Q), .B0(D6760_Y), .B1(D6594_Q),     .Y(D6573_Y), .A0(D831_Y));
KC_AOI22_X1 D6572 ( .A1(D6602_Q), .B0(D5266_Y), .B1(D6600_Q),     .Y(D6572_Y), .A0(D6695_Y));
KC_AOI22_X1 D6571 ( .A1(D1689_Y), .B0(D6600_Q), .B1(D1688_Y),     .Y(D6571_Y), .A0(D6602_Q));
KC_AOI22_X1 D6569 ( .A1(D6598_Q), .B0(D6689_Y), .B1(D6606_Q),     .Y(D6569_Y), .A0(D5322_Y));
KC_AOI22_X1 D6568 ( .A1(D1801_Y), .B0(D6599_Q), .B1(D157_Y),     .Y(D6568_Y), .A0(D6607_Q));
KC_AOI22_X1 D6289 ( .A1(D4823_Q), .B0(D1453_Y), .B1(D6382_Q),     .Y(D6289_Y), .A0(D3231_Y));
KC_AOI22_X1 D6223 ( .A1(D6278_Y), .B0(D6241_Y), .B1(D6249_Y),     .Y(D6223_Y), .A0(D6237_Y));
KC_AOI22_X1 D6094 ( .A1(D7662_Y), .B0(D13280_Q), .B1(D6093_Y),     .Y(D6094_Y), .A0(D266_Y));
KC_AOI22_X1 D6092 ( .A1(D7603_Y), .B0(D7512_Y), .B1(D1712_Y),     .Y(D6092_Y), .A0(D266_Y));
KC_AOI22_X1 D6004 ( .A1(D4454_Y), .B0(D7094_Y), .B1(D5950_Y),     .Y(D6004_Y), .A0(D7177_Y));
KC_AOI22_X1 D5842 ( .A1(D5906_Y), .B0(D9478_Y), .B1(D7307_Y),     .Y(D5842_Y), .A0(D5851_Y));
KC_AOI22_X1 D5832 ( .A1(D5902_Y), .B0(D6073_Q), .B1(D5829_Y),     .Y(D5832_Y), .A0(D235_Y));
KC_AOI22_X1 D5826 ( .A1(D254_Y), .B0(D5850_Y), .B1(D5935_Y),     .Y(D5826_Y), .A0(D7461_Y));
KC_AOI22_X1 D5770 ( .A1(D9476_Y), .B0(D5882_Y), .B1(D4130_Y),     .Y(D5770_Y), .A0(D7193_Y));
KC_AOI22_X1 D5765 ( .A1(D4165_Y), .B0(D7249_Y), .B1(D7264_Y),     .Y(D5765_Y), .A0(D5936_Y));
KC_AOI22_X1 D5764 ( .A1(D4133_Y), .B0(D7234_Y), .B1(D7264_Y),     .Y(D5764_Y), .A0(D5882_Y));
KC_AOI22_X1 D5757 ( .A1(D7282_Y), .B0(D4238_Y), .B1(D5789_Y),     .Y(D5757_Y), .A0(D199_Y));
KC_AOI22_X1 D5749 ( .A1(D5783_Y), .B0(D5722_Y), .B1(D5762_Y),     .Y(D5749_Y), .A0(D272_Y));
KC_AOI22_X1 D5740 ( .A1(D5816_Y), .B0(D5804_Y), .B1(D7270_Y),     .Y(D5740_Y), .A0(D4188_Y));
KC_AOI22_X1 D5739 ( .A1(D5887_Y), .B0(D4188_Y), .B1(D5901_Y),     .Y(D5739_Y), .A0(D5936_Y));
KC_AOI22_X1 D5733 ( .A1(D5936_Y), .B0(D5804_Y), .B1(D7285_Y),     .Y(D5733_Y), .A0(D1627_Y));
KC_AOI22_X1 D5732 ( .A1(D1617_Y), .B0(D5877_Y), .B1(D5684_Y),     .Y(D5732_Y), .A0(D5644_Y));
KC_AOI22_X1 D5718 ( .A1(D7240_Y), .B0(D3573_Y), .B1(D5730_Y),     .Y(D5718_Y), .A0(D7234_Y));
KC_AOI22_X1 D5715 ( .A1(D1590_Y), .B0(D5882_Y), .B1(D14_Y),     .Y(D5715_Y), .A0(D6039_Y));
KC_AOI22_X1 D5643 ( .A1(D7345_Y), .B0(D5645_Y), .B1(D4112_Y),     .Y(D5643_Y), .A0(D4131_Y));
KC_AOI22_X1 D5622 ( .A1(D5630_Q), .B0(D5509_Y), .B1(D5627_Q),     .Y(D5622_Y), .A0(D5540_Y));
KC_AOI22_X1 D5621 ( .A1(D6972_Y), .B0(D5627_Q), .B1(D6974_Y),     .Y(D5621_Y), .A0(D5630_Q));
KC_AOI22_X1 D5620 ( .A1(D4083_Q), .B0(D5498_Y), .B1(D4082_Q),     .Y(D5620_Y), .A0(D1596_Y));
KC_AOI22_X1 D5619 ( .A1(D5625_Q), .B0(D5509_Y), .B1(D5626_Q),     .Y(D5619_Y), .A0(D5540_Y));
KC_AOI22_X1 D5618 ( .A1(D6972_Y), .B0(D5626_Q), .B1(D6974_Y),     .Y(D5618_Y), .A0(D5625_Q));
KC_AOI22_X1 D5617 ( .A1(D5522_Y), .B0(D5624_Q), .B1(D6921_Y),     .Y(D5617_Y), .A0(D1348_Q));
KC_AOI22_X1 D5616 ( .A1(D1348_Q), .B0(D5498_Y), .B1(D5624_Q),     .Y(D5616_Y), .A0(D1596_Y));
KC_AOI22_X1 D5615 ( .A1(D6972_Y), .B0(D5603_Q), .B1(D6974_Y),     .Y(D5615_Y), .A0(D1288_Q));
KC_AOI22_X1 D5602 ( .A1(D1682_Y), .B0(D1499_Q), .B1(D6991_Y),     .Y(D5602_Y), .A0(D4050_Q));
KC_AOI22_X1 D5601 ( .A1(D4050_Q), .B0(D5497_Y), .B1(D1499_Q),     .Y(D5601_Y), .A0(D1082_Y));
KC_AOI22_X1 D5598 ( .A1(D1299_Q), .B0(D5498_Y), .B1(D5608_Q),     .Y(D5598_Y), .A0(D1596_Y));
KC_AOI22_X1 D5597 ( .A1(D6915_Y), .B0(D4049_Q), .B1(D6973_Y),     .Y(D5597_Y), .A0(D1500_Q));
KC_AOI22_X1 D5596 ( .A1(D1500_Q), .B0(D5542_Y), .B1(D4049_Q),     .Y(D5596_Y), .A0(D5543_Y));
KC_AOI22_X1 D5595 ( .A1(D4047_Q), .B0(D5498_Y), .B1(D4048_Q),     .Y(D5595_Y), .A0(D1596_Y));
KC_AOI22_X1 D5594 ( .A1(D5522_Y), .B0(D4048_Q), .B1(D6921_Y),     .Y(D5594_Y), .A0(D4047_Q));
KC_AOI22_X1 D5593 ( .A1(D1294_Q), .B0(D5497_Y), .B1(D1293_Q),     .Y(D5593_Y), .A0(D1082_Y));
KC_AOI22_X1 D5592 ( .A1(D1682_Y), .B0(D1293_Q), .B1(D6991_Y),     .Y(D5592_Y), .A0(D1294_Q));
KC_AOI22_X1 D5591 ( .A1(D5522_Y), .B0(D5608_Q), .B1(D6921_Y),     .Y(D5591_Y), .A0(D1299_Q));
KC_AOI22_X1 D5590 ( .A1(D1682_Y), .B0(D5607_Q), .B1(D6991_Y),     .Y(D5590_Y), .A0(D5606_Q));
KC_AOI22_X1 D5589 ( .A1(D5606_Q), .B0(D5497_Y), .B1(D5607_Q),     .Y(D5589_Y), .A0(D1082_Y));
KC_AOI22_X1 D5588 ( .A1(D1682_Y), .B0(D5604_Q), .B1(D6991_Y),     .Y(D5588_Y), .A0(D5605_Q));
KC_AOI22_X1 D5586 ( .A1(D1291_Q), .B0(D5542_Y), .B1(D4045_Q),     .Y(D5586_Y), .A0(D5543_Y));
KC_AOI22_X1 D5585 ( .A1(D5605_Q), .B0(D5497_Y), .B1(D5604_Q),     .Y(D5585_Y), .A0(D1082_Y));
KC_AOI22_X1 D5583 ( .A1(D6915_Y), .B0(D4045_Q), .B1(D6973_Y),     .Y(D5583_Y), .A0(D1291_Q));
KC_AOI22_X1 D5581 ( .A1(D6915_Y), .B0(D5631_Q), .B1(D6973_Y),     .Y(D5581_Y), .A0(D5632_Q));
KC_AOI22_X1 D5580 ( .A1(D1288_Q), .B0(D5509_Y), .B1(D5603_Q),     .Y(D5580_Y), .A0(D5540_Y));
KC_AOI22_X1 D5577 ( .A1(D6915_Y), .B0(D5629_Q), .B1(D6973_Y),     .Y(D5577_Y), .A0(D5633_Q));
KC_AOI22_X1 D5576 ( .A1(D5632_Q), .B0(D5542_Y), .B1(D5631_Q),     .Y(D5576_Y), .A0(D5543_Y));
KC_AOI22_X1 D5575 ( .A1(D5633_Q), .B0(D5542_Y), .B1(D5629_Q),     .Y(D5575_Y), .A0(D5543_Y));
KC_AOI22_X1 D5572 ( .A1(D5566_Q), .B0(D5497_Y), .B1(D5568_Q),     .Y(D5572_Y), .A0(D1082_Y));
KC_AOI22_X1 D5554 ( .A1(D5574_Q), .B0(D5497_Y), .B1(D1210_Q),     .Y(D5554_Y), .A0(D1082_Y));
KC_AOI22_X1 D5553 ( .A1(D1200_Q), .B0(D5497_Y), .B1(D1203_Q),     .Y(D5553_Y), .A0(D1082_Y));
KC_AOI22_X1 D5552 ( .A1(D1682_Y), .B0(D1210_Q), .B1(D6991_Y),     .Y(D5552_Y), .A0(D5574_Q));
KC_AOI22_X1 D5551 ( .A1(D1682_Y), .B0(D5560_Q), .B1(D6991_Y),     .Y(D5551_Y), .A0(D5561_Q));
KC_AOI22_X1 D5550 ( .A1(D1082_Y), .B0(D5560_Q), .B1(D5497_Y),     .Y(D5550_Y), .A0(D5561_Q));
KC_AOI22_X1 D5549 ( .A1(D1682_Y), .B0(D1203_Q), .B1(D6991_Y),     .Y(D5549_Y), .A0(D1200_Q));
KC_AOI22_X1 D5548 ( .A1(D6972_Y), .B0(D5569_Q), .B1(D6974_Y),     .Y(D5548_Y), .A0(D5567_Q));
KC_AOI22_X1 D5545 ( .A1(D5567_Q), .B0(D5509_Y), .B1(D5569_Q),     .Y(D5545_Y), .A0(D5540_Y));
KC_AOI22_X1 D5544 ( .A1(D1682_Y), .B0(D5568_Q), .B1(D6991_Y),     .Y(D5544_Y), .A0(D5566_Q));
KC_AOI22_X1 D5519 ( .A1(D5526_Q), .B0(D5348_Y), .B1(D5463_Q),     .Y(D5519_Y), .A0(D5407_Y));
KC_AOI22_X1 D5517 ( .A1(D5522_Y), .B0(D3972_Q), .B1(D6921_Y),     .Y(D5517_Y), .A0(D3961_Q));
KC_AOI22_X1 D5516 ( .A1(D6972_Y), .B0(D1125_Q), .B1(D6974_Y),     .Y(D5516_Y), .A0(D5528_Q));
KC_AOI22_X1 D5515 ( .A1(D5528_Q), .B0(D5509_Y), .B1(D1125_Q),     .Y(D5515_Y), .A0(D5540_Y));
KC_AOI22_X1 D5514 ( .A1(D6972_Y), .B0(D1132_Q), .B1(D6974_Y),     .Y(D5514_Y), .A0(D5525_Q));
KC_AOI22_X1 D5513 ( .A1(D5525_Q), .B0(D5509_Y), .B1(D1132_Q),     .Y(D5513_Y), .A0(D5540_Y));
KC_AOI22_X1 D5512 ( .A1(D5534_Q), .B0(D5509_Y), .B1(D1130_Q),     .Y(D5512_Y), .A0(D5540_Y));
KC_AOI22_X1 D5511 ( .A1(D6972_Y), .B0(D1130_Q), .B1(D6974_Y),     .Y(D5511_Y), .A0(D5534_Q));
KC_AOI22_X1 D5506 ( .A1(D6972_Y), .B0(D1122_Q), .B1(D6974_Y),     .Y(D5506_Y), .A0(D5531_Q));
KC_AOI22_X1 D5505 ( .A1(D3973_Q), .B0(D5498_Y), .B1(D5524_Q),     .Y(D5505_Y), .A0(D1596_Y));
KC_AOI22_X1 D5504 ( .A1(D3961_Q), .B0(D5498_Y), .B1(D3972_Q),     .Y(D5504_Y), .A0(D1596_Y));
KC_AOI22_X1 D5503 ( .A1(D5522_Y), .B0(D5524_Q), .B1(D6921_Y),     .Y(D5503_Y), .A0(D3973_Q));
KC_AOI22_X1 D5500 ( .A1(D1121_Q), .B0(D1202_Q), .B1(D5498_Y),     .Y(D5500_Y), .A0(D1596_Y));
KC_AOI22_X1 D5499 ( .A1(D5540_Y), .B0(D1122_Q), .B1(D5509_Y),     .Y(D5499_Y), .A0(D5531_Q));
KC_AOI22_X1 D5493 ( .A1(D7009_Q), .B0(D5542_Y), .B1(D1773_Q),     .Y(D5493_Y), .A0(D5543_Y));
KC_AOI22_X1 D5448 ( .A1(D1635_Q), .B0(D5348_Y), .B1(D5476_Q),     .Y(D5448_Y), .A0(D5407_Y));
KC_AOI22_X1 D5447 ( .A1(D118_Q), .B0(D5440_Y), .B1(D902_Q),     .Y(D5447_Y), .A0(D1628_Y));
KC_AOI22_X1 D5445 ( .A1(D5492_Q), .B0(D5345_Y), .B1(D5474_Q),     .Y(D5445_Y), .A0(D5346_Y));
KC_AOI22_X1 D5444 ( .A1(D5405_Y), .B0(D5476_Q), .B1(D5413_Y),     .Y(D5444_Y), .A0(D1635_Q));
KC_AOI22_X1 D5443 ( .A1(D5353_Y), .B0(D5474_Q), .B1(D5344_Y),     .Y(D5443_Y), .A0(D5492_Q));
KC_AOI22_X1 D5439 ( .A1(D5353_Y), .B0(D5468_Q), .B1(D5344_Y),     .Y(D5439_Y), .A0(D5470_Q));
KC_AOI22_X1 D5438 ( .A1(D5470_Q), .B0(D5345_Y), .B1(D5468_Q),     .Y(D5438_Y), .A0(D5346_Y));
KC_AOI22_X1 D5434 ( .A1(D5467_Q), .B0(D5345_Y), .B1(D5469_Q),     .Y(D5434_Y), .A0(D5346_Y));
KC_AOI22_X1 D5433 ( .A1(D5353_Y), .B0(D5469_Q), .B1(D5344_Y),     .Y(D5433_Y), .A0(D5467_Q));
KC_AOI22_X1 D5428 ( .A1(D5527_Q), .B0(D5348_Y), .B1(D5530_Q),     .Y(D5428_Y), .A0(D5407_Y));
KC_AOI22_X1 D5427 ( .A1(D5466_Q), .B0(D5345_Y), .B1(D5464_Q),     .Y(D5427_Y), .A0(D5346_Y));
KC_AOI22_X1 D5426 ( .A1(D5353_Y), .B0(D5464_Q), .B1(D5344_Y),     .Y(D5426_Y), .A0(D5466_Q));
KC_AOI22_X1 D5425 ( .A1(D6878_Y), .B0(D1129_Q), .B1(D6861_Y),     .Y(D5425_Y), .A0(D6967_Q));
KC_AOI22_X1 D5424 ( .A1(D117_Q), .B0(D5437_Y), .B1(D5465_Q),     .Y(D5424_Y), .A0(D5450_Y));
KC_AOI22_X1 D5423 ( .A1(D5356_Y), .B0(D1128_Q), .B1(D5354_Y),     .Y(D5423_Y), .A0(D3969_Q));
KC_AOI22_X1 D5422 ( .A1(D5529_Q), .B0(D5348_Y), .B1(D1634_Q),     .Y(D5422_Y), .A0(D5407_Y));
KC_AOI22_X1 D5421 ( .A1(D5405_Y), .B0(D5530_Q), .B1(D5413_Y),     .Y(D5421_Y), .A0(D5527_Q));
KC_AOI22_X1 D5367 ( .A1(D1637_Q), .B0(D5345_Y), .B1(D5402_Q),     .Y(D5367_Y), .A0(D5346_Y));
KC_AOI22_X1 D5364 ( .A1(D5353_Y), .B0(D5402_Q), .B1(D5344_Y),     .Y(D5364_Y), .A0(D1637_Q));
KC_AOI22_X1 D5363 ( .A1(D5405_Y), .B0(D1638_Q), .B1(D5413_Y),     .Y(D5363_Y), .A0(D906_Q));
KC_AOI22_X1 D5362 ( .A1(D906_Q), .B0(D5348_Y), .B1(D1638_Q),     .Y(D5362_Y), .A0(D5407_Y));
KC_AOI22_X1 D5352 ( .A1(D5356_Y), .B0(D5400_Q), .B1(D5354_Y),     .Y(D5352_Y), .A0(D5401_Q));
KC_AOI22_X1 D5351 ( .A1(D5401_Q), .B0(D5349_Y), .B1(D5400_Q),     .Y(D5351_Y), .A0(D5347_Y));
KC_AOI22_X1 D5343 ( .A1(D5405_Y), .B0(D5398_Q), .B1(D5413_Y),     .Y(D5343_Y), .A0(D5395_Q));
KC_AOI22_X1 D5338 ( .A1(D5395_Q), .B0(D5348_Y), .B1(D5398_Q),     .Y(D5338_Y), .A0(D5407_Y));
KC_AOI22_X1 D5337 ( .A1(D5353_Y), .B0(D5397_Q), .B1(D5344_Y),     .Y(D5337_Y), .A0(D5399_Q));
KC_AOI22_X1 D5336 ( .A1(D5399_Q), .B0(D5345_Y), .B1(D5397_Q),     .Y(D5336_Y), .A0(D5346_Y));
KC_AOI22_X1 D5335 ( .A1(D5356_Y), .B0(D5394_Q), .B1(D5354_Y),     .Y(D5335_Y), .A0(D5396_Q));
KC_AOI22_X1 D5334 ( .A1(D5495_Y), .B0(D8278_Y), .B1(D3769_Y),     .Y(D5334_Y), .A0(D8346_Y));
KC_AOI22_X1 D5333 ( .A1(D5507_Y), .B0(D8278_Y), .B1(D5276_Y),     .Y(D5333_Y), .A0(D8346_Y));
KC_AOI22_X1 D5332 ( .A1(D5494_Y), .B0(D8278_Y), .B1(D5277_Y),     .Y(D5332_Y), .A0(D8346_Y));
KC_AOI22_X1 D5292 ( .A1(D5405_Y), .B0(D5221_Q), .B1(D5413_Y),     .Y(D5292_Y), .A0(D5225_Q));
KC_AOI22_X1 D5291 ( .A1(D5230_Q), .B0(D5345_Y), .B1(D5226_Q),     .Y(D5291_Y), .A0(D5346_Y));
KC_AOI22_X1 D5290 ( .A1(D5319_Q), .B0(D5345_Y), .B1(D5320_Q),     .Y(D5290_Y), .A0(D5346_Y));
KC_AOI22_X1 D5289 ( .A1(D5229_Q), .B0(D5348_Y), .B1(D5222_Q),     .Y(D5289_Y), .A0(D5407_Y));
KC_AOI22_X1 D5287 ( .A1(D5392_Y), .B0(D5224_Q), .B1(D1554_Y),     .Y(D5287_Y), .A0(D5321_Q));
KC_AOI22_X1 D5286 ( .A1(D5353_Y), .B0(D5320_Q), .B1(D5344_Y),     .Y(D5286_Y), .A0(D5319_Q));
KC_AOI22_X1 D5285 ( .A1(D5346_Y), .B0(D5316_Q), .B1(D5345_Y),     .Y(D5285_Y), .A0(D5317_Q));
KC_AOI22_X1 D5284 ( .A1(D5315_Q), .B0(D5318_Q), .B1(D5265_Y),     .Y(D5284_Y), .A0(D5301_Y));
KC_AOI22_X1 D5283 ( .A1(D5407_Y), .B0(D5221_Q), .B1(D5348_Y),     .Y(D5283_Y), .A0(D5225_Q));
KC_AOI22_X1 D5282 ( .A1(D5353_Y), .B0(D5226_Q), .B1(D5344_Y),     .Y(D5282_Y), .A0(D5230_Q));
KC_AOI22_X1 D5281 ( .A1(D792_Q), .B0(D5349_Y), .B1(D5311_Q),     .Y(D5281_Y), .A0(D5347_Y));
KC_AOI22_X1 D5280 ( .A1(D5405_Y), .B0(D5222_Q), .B1(D5413_Y),     .Y(D5280_Y), .A0(D5229_Q));
KC_AOI22_X1 D5279 ( .A1(D5310_Q), .B0(D5349_Y), .B1(D5314_Q),     .Y(D5279_Y), .A0(D5347_Y));
KC_AOI22_X1 D5278 ( .A1(D5392_Y), .B0(D5318_Q), .B1(D1554_Y),     .Y(D5278_Y), .A0(D5315_Q));
KC_AOI22_X1 D5275 ( .A1(D5353_Y), .B0(D5316_Q), .B1(D5344_Y),     .Y(D5275_Y), .A0(D5317_Q));
KC_AOI22_X1 D5274 ( .A1(D5356_Y), .B0(D5314_Q), .B1(D5354_Y),     .Y(D5274_Y), .A0(D5310_Q));
KC_AOI22_X1 D5273 ( .A1(D5313_Q), .B0(D5265_Y), .B1(D5312_Q),     .Y(D5273_Y), .A0(D5301_Y));
KC_AOI22_X1 D5272 ( .A1(D5356_Y), .B0(D5306_Q), .B1(D5354_Y),     .Y(D5272_Y), .A0(D5309_Q));
KC_AOI22_X1 D5271 ( .A1(D5347_Y), .B0(D5306_Q), .B1(D5349_Y),     .Y(D5271_Y), .A0(D5309_Q));
KC_AOI22_X1 D5270 ( .A1(D5392_Y), .B0(D5312_Q), .B1(D1554_Y),     .Y(D5270_Y), .A0(D5313_Q));
KC_AOI22_X1 D5269 ( .A1(D5305_Q), .B0(D5349_Y), .B1(D5303_Q),     .Y(D5269_Y), .A0(D5347_Y));
KC_AOI22_X1 D5264 ( .A1(D5356_Y), .B0(D5303_Q), .B1(D5354_Y),     .Y(D5264_Y), .A0(D5305_Q));
KC_AOI22_X1 D5263 ( .A1(D786_Q), .B0(D5348_Y), .B1(D5304_Q),     .Y(D5263_Y), .A0(D5407_Y));
KC_AOI22_X1 D5262 ( .A1(D5308_Q), .B0(D5265_Y), .B1(D5307_Q),     .Y(D5262_Y), .A0(D5301_Y));
KC_AOI22_X1 D5261 ( .A1(D5392_Y), .B0(D5307_Q), .B1(D1554_Y),     .Y(D5261_Y), .A0(D5308_Q));
KC_AOI22_X1 D5257 ( .A1(D5302_Q), .B0(D5345_Y), .B1(D1636_Q),     .Y(D5257_Y), .A0(D5346_Y));
KC_AOI22_X1 D5256 ( .A1(D5405_Y), .B0(D5304_Q), .B1(D5413_Y),     .Y(D5256_Y), .A0(D786_Q));
KC_AOI22_X1 D5255 ( .A1(D5353_Y), .B0(D1636_Q), .B1(D5344_Y),     .Y(D5255_Y), .A0(D5302_Q));
KC_AOI22_X1 D5212 ( .A1(D5392_Y), .B0(D5237_Q), .B1(D1554_Y),     .Y(D5212_Y), .A0(D5236_Q));
KC_AOI22_X1 D5211 ( .A1(D5236_Q), .B0(D5265_Y), .B1(D5237_Q),     .Y(D5211_Y), .A0(D5301_Y));
KC_AOI22_X1 D5210 ( .A1(D5392_Y), .B0(D5232_Q), .B1(D1554_Y),     .Y(D5210_Y), .A0(D5228_Q));
KC_AOI22_X1 D5209 ( .A1(D5228_Q), .B0(D5265_Y), .B1(D5232_Q),     .Y(D5209_Y), .A0(D5301_Y));
KC_AOI22_X1 D5208 ( .A1(D5408_Y), .B0(D5238_Q), .B1(D1555_Y),     .Y(D5208_Y), .A0(D5239_Q));
KC_AOI22_X1 D5207 ( .A1(D5239_Q), .B0(D6689_Y), .B1(D5238_Q),     .Y(D5207_Y), .A0(D5322_Y));
KC_AOI22_X1 D5206 ( .A1(D5233_Q), .B0(D6760_Y), .B1(D675_Q),     .Y(D5206_Y), .A0(D831_Y));
KC_AOI22_X1 D5205 ( .A1(D5231_Q), .B0(D5265_Y), .B1(D5234_Q),     .Y(D5205_Y), .A0(D5301_Y));
KC_AOI22_X1 D5204 ( .A1(D5392_Y), .B0(D5234_Q), .B1(D1554_Y),     .Y(D5204_Y), .A0(D5231_Q));
KC_AOI22_X1 D5203 ( .A1(D5392_Y), .B0(D5227_Q), .B1(D1554_Y),     .Y(D5203_Y), .A0(D5223_Q));
KC_AOI22_X1 D5202 ( .A1(D5408_Y), .B0(D6659_Q), .B1(D1555_Y),     .Y(D5202_Y), .A0(D6661_Q));
KC_AOI22_X1 D5201 ( .A1(D5223_Q), .B0(D5265_Y), .B1(D5227_Q),     .Y(D5201_Y), .A0(D5301_Y));
KC_AOI22_X1 D5200 ( .A1(D5321_Q), .B0(D5265_Y), .B1(D5224_Q),     .Y(D5200_Y), .A0(D5301_Y));
KC_AOI22_X1 D5199 ( .A1(D5408_Y), .B0(D593_Q), .B1(D1555_Y),     .Y(D5199_Y), .A0(D5194_Q));
KC_AOI22_X1 D5179 ( .A1(D1801_Y), .B0(D5186_Q), .B1(D157_Y),     .Y(D5179_Y), .A0(D1643_Q));
KC_AOI22_X1 D5178 ( .A1(D590_Q), .B0(D6760_Y), .B1(D5185_Q),     .Y(D5178_Y), .A0(D831_Y));
KC_AOI22_X1 D5177 ( .A1(D1642_Q), .B0(D6760_Y), .B1(D5126_Q),     .Y(D5177_Y), .A0(D831_Y));
KC_AOI22_X1 D5176 ( .A1(D1643_Q), .B0(D6760_Y), .B1(D5186_Q),     .Y(D5176_Y), .A0(D831_Y));
KC_AOI22_X1 D5175 ( .A1(D5127_Q), .B0(D5266_Y), .B1(D1640_Q),     .Y(D5175_Y), .A0(D6695_Y));
KC_AOI22_X1 D5170 ( .A1(D1689_Y), .B0(D5196_Q), .B1(D1688_Y),     .Y(D5170_Y), .A0(D5198_Q));
KC_AOI22_X1 D5169 ( .A1(D596_Q), .B0(D6689_Y), .B1(D5197_Q),     .Y(D5169_Y), .A0(D5322_Y));
KC_AOI22_X1 D5168 ( .A1(D1689_Y), .B0(D1640_Q), .B1(D1688_Y),     .Y(D5168_Y), .A0(D5127_Q));
KC_AOI22_X1 D5167 ( .A1(D5198_Q), .B0(D5266_Y), .B1(D5196_Q),     .Y(D5167_Y), .A0(D6695_Y));
KC_AOI22_X1 D5165 ( .A1(D5408_Y), .B0(D5197_Q), .B1(D1555_Y),     .Y(D5165_Y), .A0(D596_Q));
KC_AOI22_X1 D5164 ( .A1(D5408_Y), .B0(D5195_Q), .B1(D1555_Y),     .Y(D5164_Y), .A0(D595_Q));
KC_AOI22_X1 D5163 ( .A1(D595_Q), .B0(D6689_Y), .B1(D5195_Q),     .Y(D5163_Y), .A0(D5322_Y));
KC_AOI22_X1 D5162 ( .A1(D1689_Y), .B0(D598_Q), .B1(D1688_Y),     .Y(D5162_Y), .A0(D597_Q));
KC_AOI22_X1 D5161 ( .A1(D597_Q), .B0(D5266_Y), .B1(D598_Q),     .Y(D5161_Y), .A0(D6695_Y));
KC_AOI22_X1 D5158 ( .A1(D5193_Q), .B0(D5266_Y), .B1(D5188_Q),     .Y(D5158_Y), .A0(D6695_Y));
KC_AOI22_X1 D5157 ( .A1(D5190_Q), .B0(D6760_Y), .B1(D5192_Q),     .Y(D5157_Y), .A0(D831_Y));
KC_AOI22_X1 D5156 ( .A1(D5189_Q), .B0(D5266_Y), .B1(D589_Q),     .Y(D5156_Y), .A0(D6695_Y));
KC_AOI22_X1 D5153 ( .A1(D1689_Y), .B0(D5188_Q), .B1(D1688_Y),     .Y(D5153_Y), .A0(D5193_Q));
KC_AOI22_X1 D5152 ( .A1(D5191_Q), .B0(D6760_Y), .B1(D594_Q),     .Y(D5152_Y), .A0(D831_Y));
KC_AOI22_X1 D5151 ( .A1(D1689_Y), .B0(D589_Q), .B1(D1688_Y),     .Y(D5151_Y), .A0(D5189_Q));
KC_AOI22_X1 D5150 ( .A1(D1801_Y), .B0(D5192_Q), .B1(D157_Y),     .Y(D5150_Y), .A0(D5190_Q));
KC_AOI22_X1 D5149 ( .A1(D1801_Y), .B0(D594_Q), .B1(D157_Y),     .Y(D5149_Y), .A0(D5191_Q));
KC_AOI22_X1 D5148 ( .A1(D1801_Y), .B0(D675_Q), .B1(D157_Y),     .Y(D5148_Y), .A0(D5233_Q));
KC_AOI22_X1 D5147 ( .A1(D5194_Q), .B0(D6689_Y), .B1(D593_Q),     .Y(D5147_Y), .A0(D5322_Y));
KC_AOI22_X1 D5146 ( .A1(D592_Q), .B0(D6689_Y), .B1(D5187_Q),     .Y(D5146_Y), .A0(D5322_Y));
KC_AOI22_X1 D5145 ( .A1(D5408_Y), .B0(D5187_Q), .B1(D1555_Y),     .Y(D5145_Y), .A0(D592_Q));
KC_AOI22_X1 D5144 ( .A1(D1801_Y), .B0(D5185_Q), .B1(D157_Y),     .Y(D5144_Y), .A0(D590_Q));
KC_AOI22_X1 D5143 ( .A1(D1801_Y), .B0(D5126_Q), .B1(D157_Y),     .Y(D5143_Y), .A0(D1642_Q));
KC_AOI22_X1 D5025 ( .A1(D3549_Y), .B0(D4887_Y), .B1(D5090_Y),     .Y(D5025_Y), .A0(D4907_Y));
KC_AOI22_X1 D5014 ( .A1(D5029_Y), .B0(D5022_Y), .B1(D1563_Y),     .Y(D5014_Y), .A0(D4900_Y));
KC_AOI22_X1 D4986 ( .A1(D5009_Y), .B0(D6449_Y), .B1(D4874_Y),     .Y(D4986_Y), .A0(D4877_Y));
KC_AOI22_X1 D4981 ( .A1(D5096_Y), .B0(D1900_Y), .B1(D5083_Y),     .Y(D4981_Y), .A0(D3633_Y));
KC_AOI22_X1 D4905 ( .A1(D4910_Y), .B0(D4942_Y), .B1(D4929_Y),     .Y(D4905_Y), .A0(D4908_Y));
KC_AOI22_X1 D4862 ( .A1(D4898_Y), .B0(D3410_Y), .B1(D3502_Y),     .Y(D4862_Y), .A0(D4874_Y));
KC_AOI22_X1 D4859 ( .A1(D1446_Y), .B0(D5036_Y), .B1(D3470_Y),     .Y(D4859_Y), .A0(D4900_Y));
KC_AOI22_X1 D4760 ( .A1(D4819_Q), .B0(D1453_Y), .B1(D6344_Q),     .Y(D4760_Y), .A0(D3231_Y));
KC_AOI22_X1 D4759 ( .A1(D3383_Q), .B0(D1453_Y), .B1(D6386_Q),     .Y(D4759_Y), .A0(D3231_Y));
KC_AOI22_X1 D4757 ( .A1(D4826_Q), .B0(D1453_Y), .B1(D1792_Q),     .Y(D4757_Y), .A0(D3231_Y));
KC_AOI22_X1 D4755 ( .A1(D4825_Q), .B0(D1453_Y), .B1(D1791_Q),     .Y(D4755_Y), .A0(D3231_Y));
KC_AOI22_X1 D4754 ( .A1(D1655_Q), .B0(D1453_Y), .B1(D6384_Q),     .Y(D4754_Y), .A0(D3231_Y));
KC_AOI22_X1 D4751 ( .A1(D3385_Q), .B0(D1453_Y), .B1(D452_Q),     .Y(D4751_Y), .A0(D3231_Y));
KC_AOI22_X1 D4570 ( .A1(D7787_Y), .B0(D1453_Y), .B1(D3127_Y),     .Y(D4570_Y), .A0(D4576_Y));
KC_AOI22_X1 D4423 ( .A1(D1593_Y), .B0(D4517_Y), .B1(D4481_Y),     .Y(D4423_Y), .A0(D4513_Y));
KC_AOI22_X1 D4344 ( .A1(D6007_Y), .B0(D249_Y), .B1(D7243_Y),     .Y(D4344_Y), .A0(D4361_Y));
KC_AOI22_X1 D4343 ( .A1(D4291_Y), .B0(D4301_Y), .B1(D4317_Y),     .Y(D4343_Y), .A0(D1629_Y));
KC_AOI22_X1 D4342 ( .A1(D4317_Y), .B0(D4291_Y), .B1(D4345_Y),     .Y(D4342_Y), .A0(D4361_Y));
KC_AOI22_X1 D4272 ( .A1(D4299_Y), .B0(D5936_Y), .B1(D7512_Y),     .Y(D4272_Y), .A0(D4380_Y));
KC_AOI22_X1 D4271 ( .A1(D4281_Y), .B0(D1583_Y), .B1(D4293_Y),     .Y(D4271_Y), .A0(D1629_Y));
KC_AOI22_X1 D4203 ( .A1(D4206_Y), .B0(D4244_Y), .B1(D4201_Y),     .Y(D4203_Y), .A0(D4240_Y));
KC_AOI22_X1 D4200 ( .A1(D5753_Y), .B0(D4132_Y), .B1(D4167_Y),     .Y(D4200_Y), .A0(D4149_Q));
KC_AOI22_X1 D4199 ( .A1(D4201_Y), .B0(D4239_Y), .B1(D4206_Y),     .Y(D4199_Y), .A0(D4241_Y));
KC_AOI22_X1 D4198 ( .A1(D4178_Y), .B0(D4243_Y), .B1(D5728_Y),     .Y(D4198_Y), .A0(D4122_Q));
KC_AOI22_X1 D4195 ( .A1(D4224_Y), .B0(D4158_Y), .B1(D7280_Y),     .Y(D4195_Y), .A0(D7225_Y));
KC_AOI22_X1 D4194 ( .A1(D7225_Y), .B0(D4158_Y), .B1(D7229_Y),     .Y(D4194_Y), .A0(D4136_Q));
KC_AOI22_X1 D4193 ( .A1(D4196_Y), .B0(D229_Q), .B1(D1615_Y),     .Y(D4193_Y), .A0(D8838_Y));
KC_AOI22_X1 D4192 ( .A1(D7293_Y), .B0(D7225_Y), .B1(D4168_Y),     .Y(D4192_Y), .A0(D4158_Y));
KC_AOI22_X1 D4191 ( .A1(D5881_Y), .B0(D4233_Y), .B1(D5730_Y),     .Y(D4191_Y), .A0(D4188_Y));
KC_AOI22_X1 D4190 ( .A1(D5753_Y), .B0(D4158_Y), .B1(D7282_Y),     .Y(D4190_Y), .A0(D4235_Q));
KC_AOI22_X1 D4189 ( .A1(D1613_Y), .B0(D199_Y), .B1(D7291_Y),     .Y(D4189_Y), .A0(D6039_Y));
KC_AOI22_X1 D4185 ( .A1(D4172_Y), .B0(D4237_Y), .B1(D260_Y),     .Y(D4185_Y), .A0(D232_Q));
KC_AOI22_X1 D4184 ( .A1(D7280_Y), .B0(D4245_Y), .B1(D5762_Y),     .Y(D4184_Y), .A0(D199_Y));
KC_AOI22_X1 D4183 ( .A1(D4196_Y), .B0(D4171_Y), .B1(D2090_Q),     .Y(D4183_Y), .A0(D4150_Y));
KC_AOI22_X1 D4182 ( .A1(D4133_Y), .B0(D4238_Y), .B1(D4174_Y),     .Y(D4182_Y), .A0(D5881_Y));
KC_AOI22_X1 D4181 ( .A1(D4356_Y), .B0(D4238_Y), .B1(D4370_Y),     .Y(D4181_Y), .A0(D4133_Y));
KC_AOI22_X1 D4180 ( .A1(D4250_Y), .B0(D4245_Y), .B1(D4159_Y),     .Y(D4180_Y), .A0(D4237_Y));
KC_AOI22_X1 D4179 ( .A1(D4133_Y), .B0(D4238_Y), .B1(D260_Y),     .Y(D4179_Y), .A0(D1590_Y));
KC_AOI22_X1 D4176 ( .A1(D4215_Y), .B0(D4188_Y), .B1(D4269_Y),     .Y(D4176_Y), .A0(D5863_Y));
KC_AOI22_X1 D4175 ( .A1(D4196_Y), .B0(D4237_Y), .B1(D4225_Y),     .Y(D4175_Y), .A0(D239_Q));
KC_AOI22_X1 D4164 ( .A1(D4130_Y), .B0(D4132_Y), .B1(D260_Y),     .Y(D4164_Y), .A0(D1590_Y));
KC_AOI22_X1 D4163 ( .A1(D4250_Y), .B0(D4241_Y), .B1(D4159_Y),     .Y(D4163_Y), .A0(D4239_Y));
KC_AOI22_X1 D4162 ( .A1(D4356_Y), .B0(D4132_Y), .B1(D4370_Y),     .Y(D4162_Y), .A0(D4130_Y));
KC_AOI22_X1 D4161 ( .A1(D4169_Y), .B0(D4188_Y), .B1(D4218_Y),     .Y(D4161_Y), .A0(D5863_Y));
KC_AOI22_X1 D4160 ( .A1(D4130_Y), .B0(D4132_Y), .B1(D4174_Y),     .Y(D4160_Y), .A0(D5881_Y));
KC_AOI22_X1 D4157 ( .A1(D4356_Y), .B0(D3572_Y), .B1(D4370_Y),     .Y(D4157_Y), .A0(D3573_Y));
KC_AOI22_X1 D4156 ( .A1(D4250_Y), .B0(D4244_Y), .B1(D4159_Y),     .Y(D4156_Y), .A0(D4240_Y));
KC_AOI22_X1 D4155 ( .A1(D4196_Y), .B0(D5693_Q), .B1(D1615_Y),     .Y(D4155_Y), .A0(D235_Y));
KC_AOI22_X1 D4154 ( .A1(D4129_Y), .B0(D4242_Y), .B1(D260_Y),     .Y(D4154_Y), .A0(D1590_Y));
KC_AOI22_X1 D4153 ( .A1(D4356_Y), .B0(D4242_Y), .B1(D4370_Y),     .Y(D4153_Y), .A0(D4129_Y));
KC_AOI22_X1 D4100 ( .A1(D4110_Y), .B0(D4099_Y), .B1(D4104_Y),     .Y(D4100_Y), .A0(D16135_Y));
KC_AOI22_X1 D4098 ( .A1(D7345_Y), .B0(D5645_Y), .B1(D4114_Y),     .Y(D4098_Y), .A0(D3573_Y));
KC_AOI22_X1 D4090 ( .A1(D4133_Y), .B0(D4233_Y), .B1(D236_Y),     .Y(D4090_Y), .A0(D7345_Y));
KC_AOI22_X1 D4089 ( .A1(D4130_Y), .B0(D4233_Y), .B1(D221_Y),     .Y(D4089_Y), .A0(D7345_Y));
KC_AOI22_X1 D4075 ( .A1(D5522_Y), .B0(D4082_Q), .B1(D6921_Y),     .Y(D4075_Y), .A0(D4083_Q));
KC_AOI22_X1 D4074 ( .A1(D4080_Q), .B0(D5498_Y), .B1(D4081_Q),     .Y(D4074_Y), .A0(D1596_Y));
KC_AOI22_X1 D3957 ( .A1(D5449_Y), .B0(D3974_Q), .B1(D5355_Y),     .Y(D3957_Y), .A0(D3963_Q));
KC_AOI22_X1 D3956 ( .A1(D3959_Q), .B0(D5340_Y), .B1(D3962_Q),     .Y(D3956_Y), .A0(D1628_Y));
KC_AOI22_X1 D3955 ( .A1(D3960_Q), .B0(D5340_Y), .B1(D3967_Q),     .Y(D3955_Y), .A0(D1628_Y));
KC_AOI22_X1 D3954 ( .A1(D3985_Q), .B0(D5340_Y), .B1(D3964_Q),     .Y(D3954_Y), .A0(D1628_Y));
KC_AOI22_X1 D3953 ( .A1(D5449_Y), .B0(D3964_Q), .B1(D5355_Y),     .Y(D3953_Y), .A0(D3985_Q));
KC_AOI22_X1 D3952 ( .A1(D5449_Y), .B0(D3962_Q), .B1(D5355_Y),     .Y(D3952_Y), .A0(D3959_Q));
KC_AOI22_X1 D3951 ( .A1(D1023_Q), .B0(D5345_Y), .B1(D1496_Q),     .Y(D3951_Y), .A0(D5346_Y));
KC_AOI22_X1 D3922 ( .A1(D5356_Y), .B0(D5491_Q), .B1(D5354_Y),     .Y(D3922_Y), .A0(D1019_Q));
KC_AOI22_X1 D3921 ( .A1(D3942_Q), .B0(D5349_Y), .B1(D1495_Q),     .Y(D3921_Y), .A0(D5347_Y));
KC_AOI22_X1 D3920 ( .A1(D3944_Q), .B0(D5340_Y), .B1(D3943_Q),     .Y(D3920_Y), .A0(D1628_Y));
KC_AOI22_X1 D3919 ( .A1(D5449_Y), .B0(D3943_Q), .B1(D5355_Y),     .Y(D3919_Y), .A0(D3944_Q));
KC_AOI22_X1 D3918 ( .A1(D5356_Y), .B0(D1495_Q), .B1(D5354_Y),     .Y(D3918_Y), .A0(D3942_Q));
KC_AOI22_X1 D3917 ( .A1(D3874_Q), .B0(D5348_Y), .B1(D3941_Q),     .Y(D3917_Y), .A0(D5407_Y));
KC_AOI22_X1 D3914 ( .A1(D5449_Y), .B0(D3938_Q), .B1(D5355_Y),     .Y(D3914_Y), .A0(D3935_Q));
KC_AOI22_X1 D3913 ( .A1(D3935_Q), .B0(D5340_Y), .B1(D3938_Q),     .Y(D3913_Y), .A0(D1628_Y));
KC_AOI22_X1 D3912 ( .A1(D5356_Y), .B0(D3936_Q), .B1(D5354_Y),     .Y(D3912_Y), .A0(D3934_Q));
KC_AOI22_X1 D3911 ( .A1(D3937_Q), .B0(D5348_Y), .B1(D3933_Q),     .Y(D3911_Y), .A0(D5407_Y));
KC_AOI22_X1 D3910 ( .A1(D5405_Y), .B0(D3933_Q), .B1(D5413_Y),     .Y(D3910_Y), .A0(D3937_Q));
KC_AOI22_X1 D3909 ( .A1(D1019_Q), .B0(D5349_Y), .B1(D5491_Q),     .Y(D3909_Y), .A0(D5347_Y));
KC_AOI22_X1 D3908 ( .A1(D5353_Y), .B0(D1496_Q), .B1(D5344_Y),     .Y(D3908_Y), .A0(D1023_Q));
KC_AOI22_X1 D3907 ( .A1(D5353_Y), .B0(D5472_Q), .B1(D5344_Y),     .Y(D3907_Y), .A0(D1017_Q));
KC_AOI22_X1 D3905 ( .A1(D1014_Q), .B0(D5345_Y), .B1(D5471_Q),     .Y(D3905_Y), .A0(D5346_Y));
KC_AOI22_X1 D3904 ( .A1(D5353_Y), .B0(D5471_Q), .B1(D5344_Y),     .Y(D3904_Y), .A0(D1014_Q));
KC_AOI22_X1 D3902 ( .A1(D3934_Q), .B0(D5349_Y), .B1(D3936_Q),     .Y(D3902_Y), .A0(D5347_Y));
KC_AOI22_X1 D3901 ( .A1(D1017_Q), .B0(D5345_Y), .B1(D5472_Q),     .Y(D3901_Y), .A0(D5346_Y));
KC_AOI22_X1 D3900 ( .A1(D5405_Y), .B0(D3929_Q), .B1(D5413_Y),     .Y(D3900_Y), .A0(D3925_Q));
KC_AOI22_X1 D3899 ( .A1(D5449_Y), .B0(D3931_Q), .B1(D5355_Y),     .Y(D3899_Y), .A0(D3927_Q));
KC_AOI22_X1 D3898 ( .A1(D3926_Q), .B0(D5349_Y), .B1(D3930_Q),     .Y(D3898_Y), .A0(D5347_Y));
KC_AOI22_X1 D3897 ( .A1(D5356_Y), .B0(D3930_Q), .B1(D5354_Y),     .Y(D3897_Y), .A0(D3926_Q));
KC_AOI22_X1 D3896 ( .A1(D3925_Q), .B0(D5348_Y), .B1(D3929_Q),     .Y(D3896_Y), .A0(D5407_Y));
KC_AOI22_X1 D3895 ( .A1(D3969_Q), .B0(D5349_Y), .B1(D1128_Q),     .Y(D3895_Y), .A0(D5347_Y));
KC_AOI22_X1 D3894 ( .A1(D3927_Q), .B0(D5340_Y), .B1(D3931_Q),     .Y(D3894_Y), .A0(D1628_Y));
KC_AOI22_X1 D3893 ( .A1(D1493_Q), .B0(D5349_Y), .B1(D1494_Q),     .Y(D3893_Y), .A0(D5347_Y));
KC_AOI22_X1 D3886 ( .A1(D5449_Y), .B0(D3879_Q), .B1(D5355_Y),     .Y(D3886_Y), .A0(D3880_Q));
KC_AOI22_X1 D3845 ( .A1(D3880_Q), .B0(D5340_Y), .B1(D3879_Q),     .Y(D3845_Y), .A0(D8267_Y));
KC_AOI22_X1 D3840 ( .A1(D3877_Q), .B0(D5340_Y), .B1(D3875_Q),     .Y(D3840_Y), .A0(D8267_Y));
KC_AOI22_X1 D3834 ( .A1(D5449_Y), .B0(D3875_Q), .B1(D5355_Y),     .Y(D3834_Y), .A0(D3877_Q));
KC_AOI22_X1 D3831 ( .A1(D5396_Q), .B0(D5349_Y), .B1(D5394_Q),     .Y(D3831_Y), .A0(D5347_Y));
KC_AOI22_X1 D3795 ( .A1(D665_Q), .B0(D5345_Y), .B1(D662_Q),     .Y(D3795_Y), .A0(D5346_Y));
KC_AOI22_X1 D3794 ( .A1(D3727_Q), .B0(D5348_Y), .B1(D667_Q),     .Y(D3794_Y), .A0(D5407_Y));
KC_AOI22_X1 D3793 ( .A1(D3818_Q), .B0(D5348_Y), .B1(D3726_Q),     .Y(D3793_Y), .A0(D5407_Y));
KC_AOI22_X1 D3791 ( .A1(D3819_Q), .B0(D5340_Y), .B1(D3816_Q),     .Y(D3791_Y), .A0(D8267_Y));
KC_AOI22_X1 D3790 ( .A1(D3817_Q), .B0(D5345_Y), .B1(D3725_Q),     .Y(D3790_Y), .A0(D5346_Y));
KC_AOI22_X1 D3789 ( .A1(D5353_Y), .B0(D3725_Q), .B1(D5344_Y),     .Y(D3789_Y), .A0(D3817_Q));
KC_AOI22_X1 D3788 ( .A1(D5353_Y), .B0(D662_Q), .B1(D5344_Y),     .Y(D3788_Y), .A0(D665_Q));
KC_AOI22_X1 D3787 ( .A1(D5405_Y), .B0(D667_Q), .B1(D5413_Y),     .Y(D3787_Y), .A0(D3727_Q));
KC_AOI22_X1 D3786 ( .A1(D5405_Y), .B0(D3726_Q), .B1(D5413_Y),     .Y(D3786_Y), .A0(D3818_Q));
KC_AOI22_X1 D3785 ( .A1(D5449_Y), .B0(D3741_Q), .B1(D5355_Y),     .Y(D3785_Y), .A0(D3740_Q));
KC_AOI22_X1 D3784 ( .A1(D5449_Y), .B0(D3816_Q), .B1(D5355_Y),     .Y(D3784_Y), .A0(D3819_Q));
KC_AOI22_X1 D3782 ( .A1(D3810_Q), .B0(D5349_Y), .B1(D790_Q),     .Y(D3782_Y), .A0(D5347_Y));
KC_AOI22_X1 D3781 ( .A1(D5449_Y), .B0(D3812_Q), .B1(D5355_Y),     .Y(D3781_Y), .A0(D3815_Q));
KC_AOI22_X1 D3780 ( .A1(D5356_Y), .B0(D790_Q), .B1(D5354_Y),     .Y(D3780_Y), .A0(D3810_Q));
KC_AOI22_X1 D3779 ( .A1(D5356_Y), .B0(D3813_Q), .B1(D5354_Y),     .Y(D3779_Y), .A0(D3811_Q));
KC_AOI22_X1 D3778 ( .A1(D3815_Q), .B0(D5340_Y), .B1(D3812_Q),     .Y(D3778_Y), .A0(D8267_Y));
KC_AOI22_X1 D3777 ( .A1(D3811_Q), .B0(D5349_Y), .B1(D3813_Q),     .Y(D3777_Y), .A0(D5347_Y));
KC_AOI22_X1 D3775 ( .A1(D5449_Y), .B0(D3804_Q), .B1(D5355_Y),     .Y(D3775_Y), .A0(D3807_Q));
KC_AOI22_X1 D3774 ( .A1(D3807_Q), .B0(D5340_Y), .B1(D3804_Q),     .Y(D3774_Y), .A0(D8267_Y));
KC_AOI22_X1 D3773 ( .A1(D3808_Q), .B0(D5348_Y), .B1(D3806_Q),     .Y(D3773_Y), .A0(D5407_Y));
KC_AOI22_X1 D3772 ( .A1(D5405_Y), .B0(D3806_Q), .B1(D5413_Y),     .Y(D3772_Y), .A0(D3808_Q));
KC_AOI22_X1 D3771 ( .A1(D3801_Q), .B0(D5348_Y), .B1(D3800_Q),     .Y(D3771_Y), .A0(D5407_Y));
KC_AOI22_X1 D3770 ( .A1(D3799_Q), .B0(D5349_Y), .B1(D3805_Q),     .Y(D3770_Y), .A0(D5347_Y));
KC_AOI22_X1 D3768 ( .A1(D3802_Q), .B0(D5340_Y), .B1(D1497_Q),     .Y(D3768_Y), .A0(D8267_Y));
KC_AOI22_X1 D3767 ( .A1(D5356_Y), .B0(D3805_Q), .B1(D5354_Y),     .Y(D3767_Y), .A0(D3799_Q));
KC_AOI22_X1 D3766 ( .A1(D5449_Y), .B0(D1497_Q), .B1(D5355_Y),     .Y(D3766_Y), .A0(D3802_Q));
KC_AOI22_X1 D3765 ( .A1(D5405_Y), .B0(D3800_Q), .B1(D5413_Y),     .Y(D3765_Y), .A0(D3801_Q));
KC_AOI22_X1 D3712 ( .A1(D3736_Q), .B0(D5265_Y), .B1(D3735_Q),     .Y(D3712_Y), .A0(D5301_Y));
KC_AOI22_X1 D3711 ( .A1(D5392_Y), .B0(D3735_Q), .B1(D1554_Y),     .Y(D3711_Y), .A0(D3736_Q));
KC_AOI22_X1 D3706 ( .A1(D5449_Y), .B0(D3734_Q), .B1(D5355_Y),     .Y(D3706_Y), .A0(D3739_Q));
KC_AOI22_X1 D3705 ( .A1(D3739_Q), .B0(D3734_Q), .B1(D5340_Y),     .Y(D3705_Y), .A0(D8267_Y));
KC_AOI22_X1 D3704 ( .A1(D5449_Y), .B0(D3743_Q), .B1(D5355_Y),     .Y(D3704_Y), .A0(D3742_Q));
KC_AOI22_X1 D3703 ( .A1(D3742_Q), .B0(D5340_Y), .B1(D3743_Q),     .Y(D3703_Y), .A0(D8267_Y));
KC_AOI22_X1 D3702 ( .A1(D3740_Q), .B0(D5340_Y), .B1(D3741_Q),     .Y(D3702_Y), .A0(D8267_Y));
KC_AOI22_X1 D3666 ( .A1(D3627_Q), .B0(D5265_Y), .B1(D1501_Q),     .Y(D3666_Y), .A0(D5301_Y));
KC_AOI22_X1 D3665 ( .A1(D1502_Q), .B0(D5265_Y), .B1(D3626_Q),     .Y(D3665_Y), .A0(D5301_Y));
KC_AOI22_X1 D3664 ( .A1(D3683_Q), .B0(D5265_Y), .B1(D3674_Q),     .Y(D3664_Y), .A0(D5301_Y));
KC_AOI22_X1 D3663 ( .A1(D5392_Y), .B0(D3626_Q), .B1(D1554_Y),     .Y(D3663_Y), .A0(D1502_Q));
KC_AOI22_X1 D3662 ( .A1(D5392_Y), .B0(D3674_Q), .B1(D1554_Y),     .Y(D3662_Y), .A0(D3683_Q));
KC_AOI22_X1 D3661 ( .A1(D5392_Y), .B0(D3684_Q), .B1(D1554_Y),     .Y(D3661_Y), .A0(D3685_Q));
KC_AOI22_X1 D3660 ( .A1(D3685_Q), .B0(D5265_Y), .B1(D3684_Q),     .Y(D3660_Y), .A0(D5301_Y));
KC_AOI22_X1 D3659 ( .A1(D5392_Y), .B0(D3678_Q), .B1(D1554_Y),     .Y(D3659_Y), .A0(D3672_Q));
KC_AOI22_X1 D3654 ( .A1(D5392_Y), .B0(D3679_Q), .B1(D1554_Y),     .Y(D3654_Y), .A0(D3680_Q));
KC_AOI22_X1 D3653 ( .A1(D3672_Q), .B0(D5265_Y), .B1(D3678_Q),     .Y(D3653_Y), .A0(D5301_Y));
KC_AOI22_X1 D3652 ( .A1(D3680_Q), .B0(D5265_Y), .B1(D3679_Q),     .Y(D3652_Y), .A0(D5301_Y));
KC_AOI22_X1 D3651 ( .A1(D3682_Q), .B0(D5265_Y), .B1(D3676_Q),     .Y(D3651_Y), .A0(D5301_Y));
KC_AOI22_X1 D3650 ( .A1(D5392_Y), .B0(D3676_Q), .B1(D1554_Y),     .Y(D3650_Y), .A0(D3682_Q));
KC_AOI22_X1 D3649 ( .A1(D5392_Y), .B0(D1501_Q), .B1(D1554_Y),     .Y(D3649_Y), .A0(D3627_Q));
KC_AOI22_X1 D3534 ( .A1(D3576_Q), .B0(D4960_Y), .B1(D3560_Y),     .Y(D3534_Y), .A0(D3459_Y));
KC_AOI22_X1 D3529 ( .A1(D3502_Y), .B0(D3540_Y), .B1(D3522_Y),     .Y(D3529_Y), .A0(D3067_Y));
KC_AOI22_X1 D3524 ( .A1(D3525_Y), .B0(D3419_Y), .B1(D3575_Q),     .Y(D3524_Y), .A0(D5012_Y));
KC_AOI22_X1 D3523 ( .A1(D5060_Y), .B0(D3531_Y), .B1(D4916_Y),     .Y(D3523_Y), .A0(D3388_Q));
KC_AOI22_X1 D3513 ( .A1(D3583_Y), .B0(D4887_Y), .B1(D473_Y),     .Y(D3513_Y), .A0(D3540_Y));
KC_AOI22_X1 D3512 ( .A1(D3421_Y), .B0(D5037_Y), .B1(D3502_Y),     .Y(D3512_Y), .A0(D5012_Y));
KC_AOI22_X1 D3511 ( .A1(D3531_Y), .B0(D3540_Y), .B1(D5012_Y),     .Y(D3511_Y), .A0(D3067_Y));
KC_AOI22_X1 D3505 ( .A1(D3559_Y), .B0(D6478_Y), .B1(D3507_Y),     .Y(D3505_Y), .A0(D3552_Y));
KC_AOI22_X1 D3485 ( .A1(D3449_Y), .B0(D3540_Y), .B1(D3419_Y),     .Y(D3485_Y), .A0(D1537_Y));
KC_AOI22_X1 D3444 ( .A1(D1466_Y), .B0(D4925_Y), .B1(D1452_Y),     .Y(D3444_Y), .A0(D3416_Y));
KC_AOI22_X1 D3441 ( .A1(D460_Y), .B0(D3421_Y), .B1(D437_Y),     .Y(D3441_Y), .A0(D4925_Y));
KC_AOI22_X1 D3433 ( .A1(D4885_Y), .B0(D4926_Y), .B1(D3468_Y),     .Y(D3433_Y), .A0(D3437_Y));
KC_AOI22_X1 D3418 ( .A1(D3509_Y), .B0(D3400_Y), .B1(D3475_Y),     .Y(D3418_Y), .A0(D4920_Y));
KC_AOI22_X1 D3417 ( .A1(D5022_Y), .B0(D4897_Y), .B1(D3487_Y),     .Y(D3417_Y), .A0(D446_Q));
KC_AOI22_X1 D3402 ( .A1(D3502_Y), .B0(D4902_Y), .B1(D3453_Y),     .Y(D3402_Y), .A0(D3459_Y));
KC_AOI22_X1 D3401 ( .A1(D5044_Y), .B0(D4960_Y), .B1(D3471_Y),     .Y(D3401_Y), .A0(D3416_Y));
KC_AOI22_X1 D3136 ( .A1(D3149_Y), .B0(D3250_Y), .B1(D3129_Y),     .Y(D3136_Y), .A0(D3349_Y));
KC_AOI22_X1 D3033 ( .A1(D3085_Y), .B0(D3068_Y), .B1(D3075_Y),     .Y(D3033_Y), .A0(D3074_Y));
KC_AOI22_X1 D2613 ( .A1(D15632_Y), .B0(D15658_Y), .B1(D2616_Y),     .Y(D2613_Y), .A0(D15484_Y));
KC_AOI22_X1 D2612 ( .A1(D15488_Y), .B0(D15489_Y), .B1(D15468_Y),     .Y(D2612_Y), .A0(D2616_Y));
KC_AOI22_X1 D2602 ( .A1(D13525_Y), .B0(D15670_Q), .B1(D2475_Y),     .Y(D2602_Y), .A0(D14871_Q));
KC_AOI22_X1 D2601 ( .A1(D2476_Y), .B0(D16363_Q), .B1(D13629_Y),     .Y(D2601_Y), .A0(D16360_Q));
KC_AOI22_X1 D2600 ( .A1(D14172_Y), .B0(D16360_Q), .B1(D14252_Y),     .Y(D2600_Y), .A0(D1155_Q));
KC_AOI22_X1 D2599 ( .A1(D14175_Y), .B0(D144_Q), .B1(D14174_Y),     .Y(D2599_Y), .A0(D15874_Q));
KC_AOI22_X1 D2598 ( .A1(D2475_Y), .B0(D15873_Q), .B1(D13525_Y),     .Y(D2598_Y), .A0(D16361_Q));
KC_AOI22_X1 D2597 ( .A1(D13634_Y), .B0(D16390_Q), .B1(D1071_Y),     .Y(D2597_Y), .A0(D142_Q));
KC_AOI22_X1 D2594 ( .A1(D14257_Y), .B0(D16389_Q), .B1(D936_Y),     .Y(D2594_Y), .A0(D16390_Q));
KC_AOI22_X1 D2542 ( .A1(D14138_Y), .B0(D15322_Y), .B1(D14130_Y),     .Y(D2542_Y), .A0(D14878_Q));
KC_AOI22_X1 D2541 ( .A1(D14138_Y), .B0(D508_Y), .B1(D14130_Y),     .Y(D2541_Y), .A0(D2573_Q));
KC_AOI22_X1 D2540 ( .A1(D14138_Y), .B0(D14679_Y), .B1(D14130_Y),     .Y(D2540_Y), .A0(D14876_Q));
KC_AOI22_X1 D2535 ( .A1(D14176_Y), .B0(D1065_Q), .B1(D14259_Y),     .Y(D2535_Y), .A0(D953_Q));
KC_AOI22_X1 D2534 ( .A1(D13526_Y), .B0(D953_Q), .B1(D13510_Y),     .Y(D2534_Y), .A0(D952_Q));
KC_AOI22_X1 D2533 ( .A1(D14173_Y), .B0(D15670_Q), .B1(D2519_Y),     .Y(D2533_Y), .A0(D952_Q));
KC_AOI22_X1 D2532 ( .A1(D13526_Y), .B0(D14870_Q), .B1(D13510_Y),     .Y(D2532_Y), .A0(D14875_Q));
KC_AOI22_X1 D2531 ( .A1(D13710_Y), .B0(D143_Q), .B1(D1072_Y),     .Y(D2531_Y), .A0(D14304_Q));
KC_AOI22_X1 D2530 ( .A1(D2477_Y), .B0(D1048_Q), .B1(D13635_Y),     .Y(D2530_Y), .A0(D2679_Q));
KC_AOI22_X1 D2527 ( .A1(D14176_Y), .B0(D2572_Q), .B1(D14259_Y),     .Y(D2527_Y), .A0(D1231_Q));
KC_AOI22_X1 D2497 ( .A1(D14010_Y), .B0(D15329_Y), .B1(D2496_Y),     .Y(D2497_Y), .A0(D14118_Q));
KC_AOI22_X1 D2495 ( .A1(D13293_Y), .B0(D13377_Y), .B1(D768_Y),     .Y(D2495_Y), .A0(D13317_Y));
KC_AOI22_X1 D2490 ( .A1(D14256_Y), .B0(D14164_Q), .B1(D14172_Y),     .Y(D2490_Y), .A0(D12996_Q));
KC_AOI22_X1 D2489 ( .A1(D14175_Y), .B0(D13530_Q), .B1(D14174_Y),     .Y(D2489_Y), .A0(D12918_Q));
KC_AOI22_X1 D2488 ( .A1(D14175_Y), .B0(D930_Q), .B1(D14174_Y),     .Y(D2488_Y), .A0(D12919_Q));
KC_AOI22_X1 D2485 ( .A1(D14173_Y), .B0(D13706_Q), .B1(D14171_Y),     .Y(D2485_Y), .A0(D14238_Q));
KC_AOI22_X1 D2484 ( .A1(D14176_Y), .B0(D13051_Q), .B1(D14259_Y),     .Y(D2484_Y), .A0(D14305_Q));
KC_AOI22_X1 D2483 ( .A1(D14257_Y), .B0(D1152_Q), .B1(D14254_Y),     .Y(D2483_Y), .A0(D2515_Q));
KC_AOI22_X1 D2482 ( .A1(D14255_Y), .B0(D13770_Q), .B1(D14252_Y),     .Y(D2482_Y), .A0(D14308_Q));
KC_AOI22_X1 D2481 ( .A1(D14176_Y), .B0(D1235_Q), .B1(D14259_Y),     .Y(D2481_Y), .A0(D14301_Q));
KC_AOI22_X1 D2480 ( .A1(D13526_Y), .B0(D1382_Q), .B1(D13510_Y),     .Y(D2480_Y), .A0(D14375_Q));
KC_AOI22_X1 D2479 ( .A1(D14255_Y), .B0(D13810_Q), .B1(D14252_Y),     .Y(D2479_Y), .A0(D1401_Q));
KC_AOI22_X1 D2437 ( .A1(D2431_Y), .B0(D13375_Y), .B1(D13377_Y),     .Y(D2437_Y), .A0(D13317_Y));
KC_AOI22_X1 D2424 ( .A1(D2427_Y), .B0(D13466_Y), .B1(D2447_Y),     .Y(D2424_Y), .A0(D12918_Q));
KC_AOI22_X1 D2415 ( .A1(D12422_Y), .B0(D2416_Y), .B1(D12933_Y),     .Y(D2415_Y), .A0(D12879_Y));
KC_AOI22_X1 D2412 ( .A1(D13526_Y), .B0(D14301_Q), .B1(D13510_Y),     .Y(D2412_Y), .A0(D13765_Q));
KC_AOI22_X1 D2404 ( .A1(D13229_Y), .B0(D13218_Y), .B1(D12685_Q),     .Y(D2404_Y), .A0(D13213_Q));
KC_AOI22_X1 D2369 ( .A1(D12834_Y), .B0(D2418_Y), .B1(D13001_Y),     .Y(D2369_Y), .A0(D12879_Y));
KC_AOI22_X1 D2368 ( .A1(D11950_Y), .B0(D12976_Q), .B1(D11953_Y),     .Y(D2368_Y), .A0(D2387_Q));
KC_AOI22_X1 D2367 ( .A1(D1308_Q), .B0(D12025_Y), .B1(D128_Q),     .Y(D2367_Y), .A0(D2301_Y));
KC_AOI22_X1 D2366 ( .A1(D12047_Y), .B0(D128_Q), .B1(D12015_Y),     .Y(D2366_Y), .A0(D1308_Q));
KC_AOI22_X1 D2324 ( .A1(D12987_Q), .B0(D11991_Y), .B1(D2389_Q),     .Y(D2324_Y), .A0(D2277_Y));
KC_AOI22_X1 D2323 ( .A1(D2351_Q), .B0(D11929_Y), .B1(D2352_Q),     .Y(D2323_Y), .A0(D11930_Y));
KC_AOI22_X1 D2322 ( .A1(D2271_Y), .B0(D12467_Q), .B1(D2273_Y),     .Y(D2322_Y), .A0(D12468_Q));
KC_AOI22_X1 D2320 ( .A1(D12450_Q), .B0(D11951_Y), .B1(D12453_Q),     .Y(D2320_Y), .A0(D11981_Y));
KC_AOI22_X1 D2319 ( .A1(D11989_Y), .B0(D12453_Q), .B1(D11949_Y),     .Y(D2319_Y), .A0(D12450_Q));
KC_AOI22_X1 D2318 ( .A1(D2321_Y), .B0(D8340_Y), .B1(D13056_Y),     .Y(D2318_Y), .A0(D8348_Y));
KC_AOI22_X1 D2317 ( .A1(D1031_Q), .B0(D11929_Y), .B1(D12977_Q),     .Y(D2317_Y), .A0(D11930_Y));
KC_AOI22_X1 D2316 ( .A1(D2271_Y), .B0(D12977_Q), .B1(D2273_Y),     .Y(D2316_Y), .A0(D1031_Q));
KC_AOI22_X1 D2315 ( .A1(D12452_Q), .B0(D11952_Y), .B1(D12458_Q),     .Y(D2315_Y), .A0(D2272_Y));
KC_AOI22_X1 D2314 ( .A1(D12455_Q), .B0(D11952_Y), .B1(D12454_Q),     .Y(D2314_Y), .A0(D2272_Y));
KC_AOI22_X1 D2313 ( .A1(D12483_Y), .B0(D8340_Y), .B1(D13066_Y),     .Y(D2313_Y), .A0(D8348_Y));
KC_AOI22_X1 D2275 ( .A1(D2293_Q), .B0(D11991_Y), .B1(D2350_Q),     .Y(D2275_Y), .A0(D2277_Y));
KC_AOI22_X1 D2274 ( .A1(D11863_Q), .B0(D11926_Q), .B1(D11991_Y),     .Y(D2274_Y), .A0(D2277_Y));
KC_AOI22_X1 D2268 ( .A1(D11980_Q), .B0(D11929_Y), .B1(D11978_Q),     .Y(D2268_Y), .A0(D11930_Y));
KC_AOI22_X1 D2267 ( .A1(D11888_Y), .B0(D8340_Y), .B1(D12072_Y),     .Y(D2267_Y), .A0(D8348_Y));
KC_AOI22_X1 D2266 ( .A1(D2270_Y), .B0(D8340_Y), .B1(D12567_Y),     .Y(D2266_Y), .A0(D8348_Y));
KC_AOI22_X1 D2265 ( .A1(D2271_Y), .B0(D11978_Q), .B1(D2273_Y),     .Y(D2265_Y), .A0(D11980_Q));
KC_AOI22_X1 D2264 ( .A1(D10766_Y), .B0(D2288_Q), .B1(D10727_Y),     .Y(D2264_Y), .A0(D11725_Q));
KC_AOI22_X1 D2232 ( .A1(D11834_Y), .B0(D135_Q), .B1(D11232_Y),     .Y(D2232_Y), .A0(D8211_Y));
KC_AOI22_X1 D2231 ( .A1(D11887_Y), .B0(D11389_Q), .B1(D2235_Y),     .Y(D2231_Y), .A0(D8211_Y));
KC_AOI22_X1 D2207 ( .A1(D10766_Y), .B0(D10631_Q), .B1(D10727_Y),     .Y(D2207_Y), .A0(D10630_Q));
KC_AOI22_X1 D2201 ( .A1(D11754_Y), .B0(D2221_Q), .B1(D2208_Y),     .Y(D2201_Y), .A0(D8211_Y));
KC_AOI22_X1 D2199 ( .A1(D10884_Q), .B0(D10903_Y), .B1(D914_Q),     .Y(D2199_Y), .A0(D2184_Y));
KC_AOI22_X1 D2198 ( .A1(D10892_Q), .B0(D10903_Y), .B1(D10891_Q),     .Y(D2198_Y), .A0(D2184_Y));
KC_AOI22_X1 D2197 ( .A1(D1043_Q), .B0(D2189_Y), .B1(D2255_Q),     .Y(D2197_Y), .A0(D10917_Y));
KC_AOI22_X1 D2196 ( .A1(D10394_Y), .B0(D11330_Q), .B1(D10913_Y),     .Y(D2196_Y), .A0(D10889_Q));
KC_AOI22_X1 D2195 ( .A1(D11350_Y), .B0(D8348_Y), .B1(D11815_Y),     .Y(D2195_Y), .A0(D8345_Y));
KC_AOI22_X1 D2194 ( .A1(D10394_Y), .B0(D10954_Q), .B1(D10913_Y),     .Y(D2194_Y), .A0(D10951_Q));
KC_AOI22_X1 D2193 ( .A1(D10990_Y), .B0(D10956_Q), .B1(D10912_Y),     .Y(D2193_Y), .A0(D2220_Q));
KC_AOI22_X1 D2192 ( .A1(D10881_Q), .B0(D2183_Y), .B1(D10883_Q),     .Y(D2192_Y), .A0(D11005_Y));
KC_AOI22_X1 D2191 ( .A1(D2220_Q), .B0(D2190_Y), .B1(D10956_Q),     .Y(D2191_Y), .A0(D2242_Y));
KC_AOI22_X1 D2187 ( .A1(D11006_Y), .B0(D1137_Q), .B1(D10902_Y),     .Y(D2187_Y), .A0(D10999_Q));
KC_AOI22_X1 D2186 ( .A1(D10394_Y), .B0(D2252_Q), .B1(D10913_Y),     .Y(D2186_Y), .A0(D11474_Q));
KC_AOI22_X1 D2185 ( .A1(D11474_Q), .B0(D2189_Y), .B1(D2252_Q),     .Y(D2185_Y), .A0(D10917_Y));
KC_AOI22_X1 D2182 ( .A1(D11006_Y), .B0(D10997_Q), .B1(D10902_Y),     .Y(D2182_Y), .A0(D10998_Q));
KC_AOI22_X1 D2181 ( .A1(D10998_Q), .B0(D2183_Y), .B1(D10997_Q),     .Y(D2181_Y), .A0(D11005_Y));
KC_AOI22_X1 D2180 ( .A1(D11428_Y), .B0(D11541_Q), .B1(D1194_Y),     .Y(D2180_Y), .A0(D9725_Y));
KC_AOI22_X1 D2179 ( .A1(D5461_Y), .B0(D2217_Q), .B1(D10541_Y),     .Y(D2179_Y), .A0(D11031_Q));
KC_AOI22_X1 D2178 ( .A1(D9555_Y), .B0(D11034_Q), .B1(D10541_Y),     .Y(D2178_Y), .A0(D11033_Q));
KC_AOI22_X1 D2177 ( .A1(D2216_Q), .B0(D11013_Y), .B1(D2215_Q),     .Y(D2177_Y), .A0(D10985_Y));
KC_AOI22_X1 D2172 ( .A1(D10353_Q), .B0(D2190_Y), .B1(D10354_Q),     .Y(D2172_Y), .A0(D2242_Y));
KC_AOI22_X1 D2169 ( .A1(D1983_Y), .B0(D10701_Y), .B1(D9393_Y),     .Y(D2169_Y), .A0(D10311_Q));
KC_AOI22_X1 D2134 ( .A1(D10431_Q), .B0(D2190_Y), .B1(D10430_Q),     .Y(D2134_Y), .A0(D2242_Y));
KC_AOI22_X1 D2133 ( .A1(D10990_Y), .B0(D917_Q), .B1(D10912_Y),     .Y(D2133_Y), .A0(D10352_Q));
KC_AOI22_X1 D2130 ( .A1(D11014_Y), .B0(D10991_Q), .B1(D11012_Y),     .Y(D2130_Y), .A0(D10512_Q));
KC_AOI22_X1 D2129 ( .A1(D1144_Y), .B0(D2156_Q), .B1(D10535_Y),     .Y(D2129_Y), .A0(D10546_Q));
KC_AOI22_X1 D2128 ( .A1(D2170_Y), .B0(D10991_Q), .B1(D10560_Y),     .Y(D2128_Y), .A0(D10512_Q));
KC_AOI22_X1 D2126 ( .A1(D10033_Q), .B0(D8901_Y), .B1(D9983_Q),     .Y(D2126_Y), .A0(D9990_Y));
KC_AOI22_X1 D2125 ( .A1(D10047_Q), .B0(D8901_Y), .B1(D10049_Q),     .Y(D2125_Y), .A0(D9990_Y));
KC_AOI22_X1 D2124 ( .A1(D10049_Q), .B0(D8901_Y), .B1(D10051_Q),     .Y(D2124_Y), .A0(D8900_Y));
KC_AOI22_X1 D2116 ( .A1(D1983_Y), .B0(D10216_Y), .B1(D9393_Y),     .Y(D2116_Y), .A0(D10294_Q));
KC_AOI22_X1 D2115 ( .A1(D10348_Q), .B0(D2190_Y), .B1(D10351_Q),     .Y(D2115_Y), .A0(D2242_Y));
KC_AOI22_X1 D2114 ( .A1(D10990_Y), .B0(D10351_Q), .B1(D10912_Y),     .Y(D2114_Y), .A0(D10348_Q));
KC_AOI22_X1 D2113 ( .A1(D1016_Q), .B0(D2183_Y), .B1(D10418_Q),     .Y(D2113_Y), .A0(D11005_Y));
KC_AOI22_X1 D2112 ( .A1(D10554_Q), .B0(D11009_Y), .B1(D10551_Q),     .Y(D2112_Y), .A0(D11003_Y));
KC_AOI22_X1 D2019 ( .A1(D7313_Y), .B0(D7394_Y), .B1(D1472_Y),     .Y(D2019_Y), .A0(D8899_Q));
KC_AOI22_X1 D2018 ( .A1(D8824_Q), .B0(D7394_Y), .B1(D2086_Y),     .Y(D2018_Y), .A0(D7313_Y));
KC_AOI22_X1 D2017 ( .A1(D7313_Y), .B0(D7393_Y), .B1(D9023_Q),     .Y(D2017_Y), .A0(D272_Y));
KC_AOI22_X1 D2014 ( .A1(D8989_Y), .B0(D9018_Y), .B1(D8976_Y),     .Y(D2014_Y), .A0(D7490_Y));
KC_AOI22_X1 D2011 ( .A1(D7362_Y), .B0(D8061_Y), .B1(D8996_Y),     .Y(D2011_Y), .A0(D9481_Y));
KC_AOI22_X1 D2010 ( .A1(D9190_Y), .B0(D308_Y), .B1(D7959_Y),     .Y(D2010_Y), .A0(D9068_Y));
KC_AOI22_X1 D2009 ( .A1(D7958_Y), .B0(D308_Y), .B1(D8062_Y),     .Y(D2009_Y), .A0(D7473_Y));
KC_AOI22_X1 D2006 ( .A1(D334_Q), .B0(D2007_Y), .B1(D9227_Q),     .Y(D2006_Y), .A0(D9041_Y));
KC_AOI22_X1 D2005 ( .A1(D9150_Q), .B0(D9277_Q), .B1(D7494_Y),     .Y(D2005_Y), .A0(D9054_Y));
KC_AOI22_X1 D2004 ( .A1(D2043_Y), .B0(D9054_Y), .B1(D9148_Q),     .Y(D2004_Y), .A0(D9068_Y));
KC_AOI22_X1 D2000 ( .A1(D2093_Q), .B0(D9102_Y), .B1(D421_Q),     .Y(D2000_Y), .A0(D9114_Y));
KC_AOI22_X1 D1999 ( .A1(D7638_Y), .B0(D7631_Y), .B1(D453_Y),     .Y(D1999_Y), .A0(D7702_Y));
KC_AOI22_X1 D1996 ( .A1(D10145_Q), .B0(D9181_Y), .B1(D9275_Q),     .Y(D1996_Y), .A0(D7631_Y));
KC_AOI22_X1 D1882 ( .A1(D4375_Y), .B0(D1883_Y), .B1(D5864_Y),     .Y(D1882_Y), .A0(D5698_Y));
KC_AOI22_X1 D1881 ( .A1(D7181_Y), .B0(D1883_Y), .B1(D5864_Y),     .Y(D1881_Y), .A0(D7194_Y));
KC_AOI22_X1 D1875 ( .A1(D8917_Y), .B0(D1877_Y), .B1(D5864_Y),     .Y(D1875_Y), .A0(D9478_Y));
KC_AOI22_X1 D1874 ( .A1(D7362_Y), .B0(D7318_Y), .B1(D1877_Y),     .Y(D1874_Y), .A0(D9478_Y));
KC_AOI22_X1 D1866 ( .A1(D21_Y), .B0(D1870_Y), .B1(D360_Y), .Y(D1866_Y),     .A0(D12300_Y));
KC_AOI22_X1 D1842 ( .A1(D6589_Y), .B0(D676_Q), .B1(D8023_Y),     .Y(D1842_Y), .A0(D6759_Y));
KC_AOI22_X1 D1833 ( .A1(D3783_Y), .B0(D8345_Y), .B1(D10911_Y),     .Y(D1833_Y), .A0(D8278_Y));
KC_AOI22_X1 D1830 ( .A1(D7039_Y), .B0(D8538_Q), .B1(D6996_Y),     .Y(D1830_Y), .A0(D2032_Y));
KC_AOI22_X1 D1829 ( .A1(D5600_Y), .B0(D8344_Y), .B1(D1252_Y),     .Y(D1829_Y), .A0(D8346_Y));
KC_AOI22_X1 D1701 ( .A1(D1654_Q), .B0(D1453_Y), .B1(D6383_Q),     .Y(D1701_Y), .A0(D3231_Y));
KC_AOI22_X1 D1691 ( .A1(D1801_Y), .B0(D6669_Q), .B1(D157_Y),     .Y(D1691_Y), .A0(D6668_Q));
KC_AOI22_X1 D1687 ( .A1(D5461_Y), .B0(D6823_Q), .B1(D6868_Y),     .Y(D1687_Y), .A0(D6824_Q));
KC_AOI22_X1 D1686 ( .A1(D5461_Y), .B0(D6821_Q), .B1(D6868_Y),     .Y(D1686_Y), .A0(D6820_Q));
KC_AOI22_X1 D1679 ( .A1(D7010_Q), .B0(D5497_Y), .B1(D1207_Q),     .Y(D1679_Y), .A0(D1082_Y));
KC_AOI22_X1 D1678 ( .A1(D1682_Y), .B0(D1207_Q), .B1(D6991_Y),     .Y(D1678_Y), .A0(D7010_Q));
KC_AOI22_X1 D1587 ( .A1(D4356_Y), .B0(D4243_Y), .B1(D4370_Y),     .Y(D1587_Y), .A0(D4131_Y));
KC_AOI22_X1 D1566 ( .A1(D4953_Y), .B0(D1567_Y), .B1(D3378_Y),     .Y(D1566_Y), .A0(D7968_Q));
KC_AOI22_X1 D1560 ( .A1(D1565_Y), .B0(D4872_Y), .B1(D1446_Y),     .Y(D1560_Y), .A0(D4920_Y));
KC_AOI22_X1 D1559 ( .A1(D4963_Y), .B0(D4907_Y), .B1(D1600_Y),     .Y(D1559_Y), .A0(D4883_Y));
KC_AOI22_X1 D1558 ( .A1(D3533_Y), .B0(D5009_Y), .B1(D3502_Y),     .Y(D1558_Y), .A0(D3426_Y));
KC_AOI22_X1 D1551 ( .A1(D5356_Y), .B0(D1124_Q), .B1(D5354_Y),     .Y(D1551_Y), .A0(D3965_Q));
KC_AOI22_X1 D1550 ( .A1(D5405_Y), .B0(D5463_Q), .B1(D5413_Y),     .Y(D1550_Y), .A0(D5526_Q));
KC_AOI22_X1 D1549 ( .A1(D5405_Y), .B0(D1634_Q), .B1(D5413_Y),     .Y(D1549_Y), .A0(D5529_Q));
KC_AOI22_X1 D1548 ( .A1(D6915_Y), .B0(D114_Q), .B1(D6973_Y),     .Y(D1548_Y), .A0(D5570_Q));
KC_AOI22_X1 D1547 ( .A1(D5562_Q), .B0(D5542_Y), .B1(D5564_Q),     .Y(D1547_Y), .A0(D5543_Y));
KC_AOI22_X1 D1546 ( .A1(D5543_Y), .B0(D5565_Q), .B1(D5542_Y),     .Y(D1546_Y), .A0(D5571_Q));
KC_AOI22_X1 D1545 ( .A1(D5570_Q), .B0(D5542_Y), .B1(D114_Q),     .Y(D1545_Y), .A0(D5543_Y));
KC_AOI22_X1 D1544 ( .A1(D6915_Y), .B0(D5565_Q), .B1(D6973_Y),     .Y(D1544_Y), .A0(D5571_Q));
KC_AOI22_X1 D1543 ( .A1(D6915_Y), .B0(D5564_Q), .B1(D6973_Y),     .Y(D1543_Y), .A0(D5562_Q));
KC_AOI22_X1 D1542 ( .A1(D120_Q), .B0(D5509_Y), .B1(D1206_Q),     .Y(D1542_Y), .A0(D5540_Y));
KC_AOI22_X1 D1541 ( .A1(D6972_Y), .B0(D1206_Q), .B1(D6974_Y),     .Y(D1541_Y), .A0(D120_Q));
KC_AOI22_X1 D1540 ( .A1(D6915_Y), .B0(D5609_Q), .B1(D6973_Y),     .Y(D1540_Y), .A0(D1639_Q));
KC_AOI22_X1 D1539 ( .A1(D1639_Q), .B0(D5542_Y), .B1(D5609_Q),     .Y(D1539_Y), .A0(D5543_Y));
KC_AOI22_X1 D1410 ( .A1(D5405_Y), .B0(D3941_Q), .B1(D5413_Y),     .Y(D1410_Y), .A0(D3874_Q));
KC_AOI22_X1 D1409 ( .A1(D3963_Q), .B0(D5340_Y), .B1(D3974_Q),     .Y(D1409_Y), .A0(D1628_Y));
KC_AOI22_X1 D1408 ( .A1(D5449_Y), .B0(D3967_Q), .B1(D5355_Y),     .Y(D1408_Y), .A0(D3960_Q));
KC_AOI22_X1 D1339 ( .A1(D15241_Y), .B0(D15239_Y), .B1(D15239_Y),     .Y(D1339_Y), .A0(D15239_Y));
KC_AOI22_X1 D1337 ( .A1(D11990_Y), .B0(D1369_Q), .B1(D12011_Y),     .Y(D1337_Y), .A0(D13145_Q));
KC_AOI22_X1 D1336 ( .A1(D5522_Y), .B0(D7043_Q), .B1(D6921_Y),     .Y(D1336_Y), .A0(D7042_Q));
KC_AOI22_X1 D1335 ( .A1(D1349_Q), .B0(D5498_Y), .B1(D7076_Q),     .Y(D1335_Y), .A0(D1596_Y));
KC_AOI22_X1 D1334 ( .A1(D10610_Q), .B0(D11013_Y), .B1(D10613_Q),     .Y(D1334_Y), .A0(D10985_Y));
KC_AOI22_X1 D1333 ( .A1(D5522_Y), .B0(D7079_Q), .B1(D6921_Y),     .Y(D1333_Y), .A0(D1352_Q));
KC_AOI22_X1 D1332 ( .A1(D5522_Y), .B0(D7076_Q), .B1(D6921_Y),     .Y(D1332_Y), .A0(D1349_Q));
KC_AOI22_X1 D1331 ( .A1(D5522_Y), .B0(D4081_Q), .B1(D6921_Y),     .Y(D1331_Y), .A0(D4080_Q));
KC_AOI22_X1 D1280 ( .A1(D13524_Y), .B0(D15233_Q), .B1(D14224_Y),     .Y(D1280_Y), .A0(D1325_Q));
KC_AOI22_X1 D1279 ( .A1(D14257_Y), .B0(D15994_Q), .B1(D14254_Y),     .Y(D1279_Y), .A0(D15993_Q));
KC_AOI22_X1 D1278 ( .A1(D14253_Y), .B0(D15233_Q), .B1(D936_Y),     .Y(D1278_Y), .A0(D15213_Q));
KC_AOI22_X1 D1277 ( .A1(D14255_Y), .B0(D1383_Q), .B1(D14252_Y),     .Y(D1277_Y), .A0(D1380_Q));
KC_AOI22_X1 D1266 ( .A1(D11073_Q), .B0(D11011_Y), .B1(D11075_Q),     .Y(D1266_Y), .A0(D11010_Y));
KC_AOI22_X1 D1265 ( .A1(D13117_Q), .B0(D12012_Y), .B1(D13119_Q),     .Y(D1265_Y), .A0(D12052_Y));
KC_AOI22_X1 D1263 ( .A1(D2170_Y), .B0(D11080_Q), .B1(D10560_Y),     .Y(D1263_Y), .A0(D11079_Q));
KC_AOI22_X1 D1262 ( .A1(D12016_Y), .B0(D13119_Q), .B1(D12026_Y),     .Y(D1262_Y), .A0(D13117_Q));
KC_AOI22_X1 D1261 ( .A1(D11584_Q), .B0(D12012_Y), .B1(D1317_Q),     .Y(D1261_Y), .A0(D12052_Y));
KC_AOI22_X1 D1260 ( .A1(D9265_Y), .B0(D11012_Y), .B1(D11082_Q),     .Y(D1260_Y), .A0(D11014_Y));
KC_AOI22_X1 D1259 ( .A1(D7053_Q), .B0(D5498_Y), .B1(D7052_Q),     .Y(D1259_Y), .A0(D1596_Y));
KC_AOI22_X1 D1258 ( .A1(D1290_Q), .B0(D11011_Y), .B1(D1297_Q),     .Y(D1258_Y), .A0(D11010_Y));
KC_AOI22_X1 D1257 ( .A1(D1296_Q), .B0(D11009_Y), .B1(D8639_Q),     .Y(D1257_Y), .A0(D11003_Y));
KC_AOI22_X1 D1256 ( .A1(D5522_Y), .B0(D7052_Q), .B1(D6921_Y),     .Y(D1256_Y), .A0(D7053_Q));
KC_AOI22_X1 D1254 ( .A1(D8634_Q), .B0(D5497_Y), .B1(D8641_Q),     .Y(D1254_Y), .A0(D1082_Y));
KC_AOI22_X1 D1253 ( .A1(D1292_Q), .B0(D5498_Y), .B1(D7045_Q),     .Y(D1253_Y), .A0(D1596_Y));
KC_AOI22_X1 D1251 ( .A1(D5522_Y), .B0(D7045_Q), .B1(D6921_Y),     .Y(D1251_Y), .A0(D1292_Q));
KC_AOI22_X1 D1250 ( .A1(D5522_Y), .B0(D7082_Q), .B1(D6921_Y),     .Y(D1250_Y), .A0(D7085_Q));
KC_AOI22_X1 D1183 ( .A1(D13525_Y), .B0(D15231_Q), .B1(D2475_Y),     .Y(D1183_Y), .A0(D1232_Q));
KC_AOI22_X1 D1181 ( .A1(D13717_Y), .B0(D14308_Q), .B1(D13727_Y),     .Y(D1181_Y), .A0(D1401_Q));
KC_AOI22_X1 D1180 ( .A1(D14258_Y), .B0(D13759_Q), .B1(D2519_Y),     .Y(D1180_Y), .A0(D1375_Q));
KC_AOI22_X1 D1178 ( .A1(D14258_Y), .B0(D13813_Q), .B1(D2519_Y),     .Y(D1178_Y), .A0(D13805_Q));
KC_AOI22_X1 D1175 ( .A1(D13103_Y), .B0(D12043_Q), .B1(D11524_Y),     .Y(D1175_Y), .A0(D9725_Y));
KC_AOI22_X1 D1174 ( .A1(D12047_Y), .B0(D1222_Q), .B1(D12015_Y),     .Y(D1174_Y), .A0(D132_Q));
KC_AOI22_X1 D1173 ( .A1(D13058_Y), .B0(D1246_Q), .B1(D11515_Y),     .Y(D1173_Y), .A0(D9725_Y));
KC_AOI22_X1 D1172 ( .A1(D12570_Y), .B0(D8589_Q), .B1(D1193_Y),     .Y(D1172_Y), .A0(D2032_Y));
KC_AOI22_X1 D1171 ( .A1(D13072_Y), .B0(D12042_Q), .B1(D11526_Y),     .Y(D1171_Y), .A0(D2032_Y));
KC_AOI22_X1 D1170 ( .A1(D7006_Q), .B0(D5497_Y), .B1(D7007_Q),     .Y(D1170_Y), .A0(D1082_Y));
KC_AOI22_X1 D1169 ( .A1(D10544_Q), .B0(D11012_Y), .B1(D2159_Q),     .Y(D1169_Y), .A0(D11014_Y));
KC_AOI22_X1 D1168 ( .A1(D10559_Y), .B0(D1303_Q), .B1(D10558_Y),     .Y(D1168_Y), .A0(D1302_Q));
KC_AOI22_X1 D1167 ( .A1(D1211_Q), .B0(D5509_Y), .B1(D7004_Q),     .Y(D1167_Y), .A0(D5540_Y));
KC_AOI22_X1 D1094 ( .A1(D14253_Y), .B0(D2474_Q), .B1(D936_Y),     .Y(D1094_Y), .A0(D13704_Q));
KC_AOI22_X1 D1093 ( .A1(D1073_Y), .B0(D15874_Q), .B1(D13636_Y),     .Y(D1093_Y), .A0(D1155_Q));
KC_AOI22_X1 D1090 ( .A1(D13634_Y), .B0(D14298_Q), .B1(D1071_Y),     .Y(D1090_Y), .A0(D13704_Q));
KC_AOI22_X1 D1089 ( .A1(D1072_Y), .B0(D14308_Q), .B1(D13710_Y),     .Y(D1089_Y), .A0(D1235_Q));
KC_AOI22_X1 D1088 ( .A1(D11969_Y), .B0(D13032_Q), .B1(D11948_Y),     .Y(D1088_Y), .A0(D13034_Q));
KC_AOI22_X1 D1086 ( .A1(D10917_Y), .B0(D11473_Q), .B1(D2189_Y),     .Y(D1086_Y), .A0(D11472_Q));
KC_AOI22_X1 D1085 ( .A1(D10904_Y), .B0(D11467_Q), .B1(D979_Y),     .Y(D1085_Y), .A0(D11471_Q));
KC_AOI22_X1 D1083 ( .A1(D113_Q), .B0(D5498_Y), .B1(D5573_Q),     .Y(D1083_Y), .A0(D1596_Y));
KC_AOI22_X1 D1081 ( .A1(D5522_Y), .B0(D5573_Q), .B1(D6921_Y),     .Y(D1081_Y), .A0(D113_Q));
KC_AOI22_X1 D1080 ( .A1(D6915_Y), .B0(D1773_Q), .B1(D6973_Y),     .Y(D1080_Y), .A0(D7009_Q));
KC_AOI22_X1 D1079 ( .A1(D5522_Y), .B0(D1202_Q), .B1(D6921_Y),     .Y(D1079_Y), .A0(D1121_Q));
KC_AOI22_X1 D989 ( .A1(D14253_Y), .B0(D14265_Q), .B1(D936_Y),     .Y(D989_Y), .A0(D2391_Q));
KC_AOI22_X1 D987 ( .A1(D13636_Y), .B0(D15711_Q), .B1(D1073_Y),     .Y(D987_Y), .A0(D924_Q));
KC_AOI22_X1 D986 ( .A1(D1073_Y), .B0(D15793_Q), .B1(D13636_Y),     .Y(D986_Y), .A0(D16317_Q));
KC_AOI22_X1 D982 ( .A1(D12985_Q), .B0(D11991_Y), .B1(D12986_Q),     .Y(D982_Y), .A0(D2277_Y));
KC_AOI22_X1 D978 ( .A1(D12979_Q), .B0(D11952_Y), .B1(D12978_Q),     .Y(D978_Y), .A0(D2272_Y));
KC_AOI22_X1 D977 ( .A1(D5461_Y), .B0(D902_Q), .B1(D6868_Y), .Y(D977_Y),     .A0(D118_Q));
KC_AOI22_X1 D975 ( .A1(D3923_Y), .B0(D1930_Q), .B1(D8433_Y),     .Y(D975_Y), .A0(D6759_Y));
KC_AOI22_X1 D974 ( .A1(D11006_Y), .B0(D10420_Q), .B1(D10902_Y),     .Y(D974_Y), .A0(D1021_Q));
KC_AOI22_X1 D971 ( .A1(D5450_Y), .B0(D1775_Q), .B1(D5437_Y),     .Y(D971_Y), .A0(D1012_Q));
KC_AOI22_X1 D969 ( .A1(D6964_Q), .B0(D5437_Y), .B1(D6968_Q),     .Y(D969_Y), .A0(D5450_Y));
KC_AOI22_X1 D967 ( .A1(D3965_Q), .B0(D5349_Y), .B1(D1124_Q),     .Y(D967_Y), .A0(D5347_Y));
KC_AOI22_X1 D873 ( .A1(D14841_Y), .B0(D2604_Y), .B1(D14850_Y),     .Y(D873_Y), .A0(D15472_Y));
KC_AOI22_X1 D871 ( .A1(D14146_Y), .B0(D14109_Q), .B1(D14147_Y),     .Y(D871_Y), .A0(D817_Q));
KC_AOI22_X1 D867 ( .A1(D12391_Y), .B0(D11859_Q), .B1(D11310_Y),     .Y(D867_Y), .A0(D11255_Y));
KC_AOI22_X1 D864 ( .A1(D12381_Y), .B0(D8340_Y), .B1(D12520_Y),     .Y(D864_Y), .A0(D8348_Y));
KC_AOI22_X1 D859 ( .A1(D6918_Y), .B0(D8278_Y), .B1(D5258_Y),     .Y(D859_Y), .A0(D8346_Y));
KC_AOI22_X1 D858 ( .A1(D10990_Y), .B0(D905_Q), .B1(D10912_Y),     .Y(D858_Y), .A0(D904_Q));
KC_AOI22_X1 D759 ( .A1(D15425_Y), .B0(D16800_Y), .B1(D15529_Y),     .Y(D759_Y), .A0(D14750_Y));
KC_AOI22_X1 D758 ( .A1(D12687_Q), .B0(D14033_Y), .B1(D13259_Y),     .Y(D758_Y), .A0(D14077_Y));
KC_AOI22_X1 D750 ( .A1(D13293_Y), .B0(D13378_Y), .B1(D768_Y),     .Y(D750_Y), .A0(D13478_Y));
KC_AOI22_X1 D748 ( .A1(D683_Q), .B0(D10743_Y), .B1(D806_Q), .Y(D748_Y),     .A0(D10805_Y));
KC_AOI22_X1 D747 ( .A1(D801_Q), .B0(D10808_Y), .B1(D805_Q), .Y(D747_Y),     .A0(D10809_Y));
KC_AOI22_X1 D745 ( .A1(D10699_Y), .B0(D797_Q), .B1(D11236_Y),     .Y(D745_Y), .A0(D8211_Y));
KC_AOI22_X1 D742 ( .A1(D11753_Y), .B0(D11260_Q), .B1(D11775_Y),     .Y(D742_Y), .A0(D11255_Y));
KC_AOI22_X1 D736 ( .A1(D5366_Y), .B0(D6754_Q), .B1(D8217_Y),     .Y(D736_Y), .A0(D6759_Y));
KC_AOI22_X1 D735 ( .A1(D5356_Y), .B0(D5311_Q), .B1(D5354_Y),     .Y(D735_Y), .A0(D792_Q));
KC_AOI22_X1 D734 ( .A1(D6625_Y), .B0(D784_Q), .B1(D6726_Y), .Y(D734_Y),     .A0(D6759_Y));
KC_AOI22_X1 D732 ( .A1(D787_Q), .B0(D5345_Y), .B1(D119_Q), .Y(D732_Y),     .A0(D5346_Y));
KC_AOI22_X1 D731 ( .A1(D5353_Y), .B0(D119_Q), .B1(D5344_Y), .Y(D731_Y),     .A0(D787_Q));
KC_AOI22_X1 D638 ( .A1(D15067_Y), .B0(D2508_Y), .B1(D15449_Y),     .Y(D638_Y), .A0(D13400_Y));
KC_AOI22_X1 D633 ( .A1(D14615_Y), .B0(D15348_Y), .B1(D771_Y),     .Y(D633_Y), .A0(D15345_Y));
KC_AOI22_X1 D630 ( .A1(D11182_Q), .B0(D10808_Y), .B1(D689_Q),     .Y(D630_Y), .A0(D10809_Y));
KC_AOI22_X1 D629 ( .A1(D10672_Y), .B0(D10719_Q), .B1(D10757_Y),     .Y(D629_Y), .A0(D688_Q));
KC_AOI22_X1 D628 ( .A1(D803_Q), .B0(D10742_Y), .B1(D677_Q), .Y(D628_Y),     .A0(D10745_Y));
KC_AOI22_X1 D626 ( .A1(D682_Q), .B0(D10742_Y), .B1(D11177_Q),     .Y(D626_Y), .A0(D10745_Y));
KC_AOI22_X1 D623 ( .A1(D6661_Q), .B0(D6689_Y), .B1(D6659_Q),     .Y(D623_Y), .A0(D5322_Y));
KC_AOI22_X1 D611 ( .A1(D10766_Y), .B0(D10183_Q), .B1(D10727_Y),     .Y(D611_Y), .A0(D10185_Q));
KC_AOI22_X1 D571 ( .A1(D530_Q), .B0(D13955_Y), .B1(D14759_Y),     .Y(D571_Y), .A0(D13904_Y));
KC_AOI22_X1 D565 ( .A1(D12681_Q), .B0(D2461_Y), .B1(D607_Q),     .Y(D565_Y), .A0(D2462_Y));
KC_AOI22_X1 D563 ( .A1(D13908_Q), .B0(D13955_Y), .B1(D14772_Y),     .Y(D563_Y), .A0(D13904_Y));
KC_AOI22_X1 D562 ( .A1(D13199_Q), .B0(D13281_Y), .B1(D13198_Q),     .Y(D562_Y), .A0(D13254_Y));
KC_AOI22_X1 D559 ( .A1(D11661_Q), .B0(D10818_Y), .B1(D11656_Q),     .Y(D559_Y), .A0(D10765_Y));
KC_AOI22_X1 D557 ( .A1(D526_Q), .B0(D10818_Y), .B1(D10632_Q),     .Y(D557_Y), .A0(D10765_Y));
KC_AOI22_X1 D556 ( .A1(D10766_Y), .B0(D10184_Q), .B1(D10727_Y),     .Y(D556_Y), .A0(D127_Q));
KC_AOI22_X1 D555 ( .A1(D10766_Y), .B0(D10632_Q), .B1(D10727_Y),     .Y(D555_Y), .A0(D526_Q));
KC_AOI22_X1 D554 ( .A1(D10766_Y), .B0(D2213_Q), .B1(D10727_Y),     .Y(D554_Y), .A0(D525_Q));
KC_AOI22_X1 D551 ( .A1(D5408_Y), .B0(D6612_Q), .B1(D1555_Y),     .Y(D551_Y), .A0(D6611_Q));
KC_AOI22_X1 D550 ( .A1(D5408_Y), .B0(D6596_Q), .B1(D1555_Y),     .Y(D550_Y), .A0(D591_Q));
KC_AOI22_X1 D549 ( .A1(D5408_Y), .B0(D6606_Q), .B1(D1555_Y),     .Y(D549_Y), .A0(D6598_Q));
KC_AOI22_X1 D403 ( .A1(D4817_Q), .B0(D1453_Y), .B1(D6387_Q),     .Y(D403_Y), .A0(D3231_Y));
KC_AOI22_X1 D400 ( .A1(D4824_Q), .B0(D1453_Y), .B1(D6385_Q),     .Y(D400_Y), .A0(D3231_Y));
KC_AOI22_X1 D342 ( .A1(D1864_Y), .B0(D7473_Y), .B1(D8072_Y),     .Y(D342_Y), .A0(D363_Q));
KC_AOI22_X1 D340 ( .A1(D7576_Y), .B0(D7613_Y), .B1(D9086_Y),     .Y(D340_Y), .A0(D8072_Y));
KC_AOI22_X1 D337 ( .A1(D3321_Y), .B0(D3048_Y), .B1(D4620_Y),     .Y(D337_Y), .A0(D4687_Y));
KC_AOI22_X1 D289 ( .A1(D7345_Y), .B0(D8953_Q), .B1(D7456_Y),     .Y(D289_Y), .A0(D7_Y));
KC_AOI22_X1 D279 ( .A1(D15439_Y), .B0(D7313_Y), .B1(D10047_Q),     .Y(D279_Y), .A0(D7394_Y));
KC_AOI22_X1 D278 ( .A1(D7315_Y), .B0(D8974_Y), .B1(D7529_Y),     .Y(D278_Y), .A0(D303_Q));
KC_AOI22_X1 D252 ( .A1(D4131_Y), .B0(D4243_Y), .B1(D5904_Y),     .Y(D252_Y), .A0(D5881_Y));
KC_AOI22_X1 D251 ( .A1(D7343_Y), .B0(D6039_Y), .B1(D213_Y), .Y(D251_Y),     .A0(D7318_Y));
KC_AOI22_X1 D250 ( .A1(D40_Q), .B0(D2070_Y), .B1(D9982_Q), .Y(D250_Y),     .A0(D7393_Y));
KC_AOI22_X1 D248 ( .A1(D36_Y), .B0(D2070_Y), .B1(D147_Q), .Y(D248_Y),     .A0(D7393_Y));
KC_AOI22_X1 D207 ( .A1(D8832_Y), .B0(D209_Y), .B1(D7269_Y), .Y(D207_Y),     .A0(D2095_Y));
KC_AOI22_X1 D178 ( .A1(D7345_Y), .B0(D5645_Y), .B1(D5680_Y),     .Y(D178_Y), .A0(D4129_Y));
KC_AOI22_X1 D88 ( .A1(D2543_Y), .B0(D15479_Y), .B1(D14867_Y),     .Y(D88_Y), .A0(D2609_Y));
KC_AOI22_X1 D87 ( .A1(D2431_Y), .B0(D13375_Y), .B1(D13378_Y),     .Y(D87_Y), .A0(D13478_Y));
KC_AOI22_X1 D85 ( .A1(D2372_Y), .B0(D12879_Y), .B1(D13028_Y),     .Y(D85_Y), .A0(D13393_Y));
KC_AOI22_X1 D83 ( .A1(D694_Q), .B0(D13281_Y), .B1(D13204_Y), .Y(D83_Y),     .A0(D13254_Y));
KC_AOI22_X1 D82 ( .A1(D11969_Y), .B0(D12913_Q), .B1(D11948_Y),     .Y(D82_Y), .A0(D12912_Q));
KC_AOI22_X1 D81 ( .A1(D2387_Q), .B0(D11952_Y), .B1(D12976_Q),     .Y(D81_Y), .A0(D2272_Y));
KC_AOI22_X1 D80 ( .A1(D1087_Y), .B0(D8340_Y), .B1(D13111_Y), .Y(D80_Y),     .A0(D8348_Y));
KC_AOI22_X1 D79 ( .A1(D10394_Y), .B0(D11473_Q), .B1(D10913_Y),     .Y(D79_Y), .A0(D11472_Q));
KC_AOI22_X1 D74 ( .A1(D6081_Y), .B0(D8974_Y), .B1(D9090_Y), .Y(D74_Y),     .A0(D5936_Y));
KC_AOI22_X1 D72 ( .A1(D3009_Y), .B0(D47_Y), .B1(D148_Q), .Y(D72_Y),     .A0(D9345_Y));
KC_AOI22_X1 D66 ( .A1(D5420_Y), .B0(D6825_Q), .B1(D1893_Y), .Y(D66_Y),     .A0(D6759_Y));
KC_AOI22_X1 D63 ( .A1(D5356_Y), .B0(D1494_Q), .B1(D5354_Y), .Y(D63_Y),     .A0(D1493_Q));
KC_AOI22_X1 D62 ( .A1(D1783_Q), .B0(D5542_Y), .B1(D1784_Q), .Y(D62_Y),     .A0(D5543_Y));
KC_AOI211_X1 D16606 ( .A(D16573_Y), .Y(D16606_Y), .C1(D16611_Q),     .C0(D16603_Y), .B(D16607_Y));
KC_AOI211_X1 D16605 ( .A(D16572_Y), .Y(D16605_Y), .C1(D16613_Q),     .C0(D1374_Q), .B(D16573_Y));
KC_AOI211_X1 D16601 ( .A(D16603_Y), .Y(D16601_Y), .C1(D16595_Y),     .C0(D16600_Y), .B(D16573_Y));
KC_AOI211_X1 D16562 ( .A(D16563_Y), .Y(D16562_Y), .C1(D16561_Y),     .C0(D1340_Y), .B(D16573_Y));
KC_AOI211_X1 D16486 ( .A(D16540_Y), .Y(D16486_Y), .C1(D16513_Y),     .C0(D16511_Y), .B(D13392_Y));
KC_AOI211_X1 D16480 ( .A(D16418_Y), .Y(D16480_Y), .C1(D16481_Y),     .C0(D16410_Y), .B(D13392_Y));
KC_AOI211_X1 D16462 ( .A(D16415_Y), .Y(D16462_Y), .C1(D16463_Y),     .C0(D1378_Q), .B(D16372_Y));
KC_AOI211_X1 D16418 ( .A(D16470_Q), .Y(D16418_Y), .C1(D16424_Y),     .C0(D16423_Y), .B(D16417_Y));
KC_AOI211_X1 D16189 ( .A(D16264_Y), .Y(D16189_Y), .C1(D16226_Q),     .C0(D16252_Y), .B(D13392_Y));
KC_AOI211_X1 D16186 ( .A(D16112_Y), .Y(D16186_Y), .C1(D16170_Y),     .C0(D16188_Y), .B(D16134_Y));
KC_AOI211_X1 D16003 ( .A(D16010_Q), .Y(D16003_Y), .C1(D16007_Y),     .C0(D15228_Y), .B(D1339_Y));
KC_AOI211_X1 D15722 ( .A(D15777_Y), .Y(D15722_Y), .C1(D2641_Q),     .C0(D15728_Y), .B(D15819_Y));
KC_AOI211_X1 D15477 ( .A(D15544_Y), .Y(D15477_Y), .C1(D15633_Y),     .C0(D15485_Y), .B(D15481_Y));
KC_AOI211_X1 D15369 ( .A(D15417_Y), .Y(D15369_Y), .C1(D15513_Y),     .C0(D15378_Y), .B(D15372_Y));
KC_AOI211_X1 D15341 ( .A(D15414_Y), .Y(D15341_Y), .C1(D15378_Y),     .C0(D15551_Y), .B(D15427_Y));
KC_AOI211_X1 D14925 ( .A(D96_Y), .Y(D14925_Y), .C1(D14828_Y),     .C0(D14926_Y), .B(D14923_Y));
KC_AOI211_X1 D14849 ( .A(D14848_Y), .Y(D14849_Y), .C1(D14815_Q),     .C0(D14726_Y), .B(D14909_Y));
KC_AOI211_X1 D14736 ( .A(D14734_Y), .Y(D14736_Y), .C1(D14735_Y),     .C0(D12856_Q), .B(D14775_Y));
KC_AOI211_X1 D14731 ( .A(D13392_Y), .Y(D14731_Y), .C1(D16398_Y),     .C0(D13330_Y), .B(D14807_Y));
KC_AOI211_X1 D14545 ( .A(D14567_Y), .Y(D14545_Y), .C1(D2546_Y),     .C0(D2548_Y), .B(D14553_Y));
KC_AOI211_X1 D14485 ( .A(D15227_Y), .Y(D14485_Y), .C1(D1376_Q),     .C0(D15226_Y), .B(D14484_Y));
KC_AOI211_X1 D14480 ( .A(D14479_Y), .Y(D14480_Y), .C1(D14490_Q),     .C0(D14486_Y), .B(D14488_Y));
KC_AOI211_X1 D14432 ( .A(D14358_Y), .Y(D14432_Y), .C1(D13771_Q),     .C0(D14440_Y), .B(D14372_Y));
KC_AOI211_X1 D14427 ( .A(D14399_Y), .Y(D14427_Y), .C1(D1321_Q),     .C0(D14430_Y), .B(D14468_Y));
KC_AOI211_X1 D14419 ( .A(D14441_Y), .Y(D14419_Y), .C1(D13815_Q),     .C0(D14413_Y), .B(D1274_Y));
KC_AOI211_X1 D14415 ( .A(D15197_Y), .Y(D14415_Y), .C1(D1323_Q),     .C0(D14418_Y), .B(D14454_Y));
KC_AOI211_X1 D14410 ( .A(D14451_Y), .Y(D14410_Y), .C1(D14475_Q),     .C0(D14414_Y), .B(D14467_Y));
KC_AOI211_X1 D14406 ( .A(D14443_Y), .Y(D14406_Y), .C1(D13814_Q),     .C0(D14424_Y), .B(D14465_Y));
KC_AOI211_X1 D14405 ( .A(D15975_Y), .Y(D14405_Y), .C1(D1325_Q),     .C0(D1269_Y), .B(D14407_Y));
KC_AOI211_X1 D14404 ( .A(D15205_Y), .Y(D14404_Y), .C1(D15213_Q),     .C0(D15165_Y), .B(D14431_Y));
KC_AOI211_X1 D14360 ( .A(D15203_Y), .Y(D14360_Y), .C1(D15218_Q),     .C0(D15107_Y), .B(D14439_Y));
KC_AOI211_X1 D14351 ( .A(D14352_Y), .Y(D14351_Y), .C1(D14375_Q),     .C0(D14356_Y), .B(D14371_Y));
KC_AOI211_X1 D14344 ( .A(D15118_Y), .Y(D14344_Y), .C1(D2524_Q),     .C0(D14348_Y), .B(D14349_Y));
KC_AOI211_X1 D14329 ( .A(D15923_Y), .Y(D14329_Y), .C1(D1232_Q),     .C0(D15106_Y), .B(D14336_Y));
KC_AOI211_X1 D14275 ( .A(D14289_Y), .Y(D14275_Y), .C1(D15890_Y),     .C0(D14295_Y), .B(D14204_Y));
KC_AOI211_X1 D14128 ( .A(D14906_Y), .Y(D14128_Y), .C1(D13983_Y),     .C0(D14852_Y), .B(D14843_Y));
KC_AOI211_X1 D14124 ( .A(D14203_Y), .Y(D14124_Y), .C1(D13975_Y),     .C0(D872_Y), .B(D14208_Y));
KC_AOI211_X1 D13936 ( .A(D14017_Y), .Y(D13936_Y), .C1(D13848_Y),     .C0(D13933_Y), .B(D13890_Y));
KC_AOI211_X1 D13718 ( .A(D13752_Y), .Y(D13718_Y), .C1(D10266_Y),     .C0(D13730_Y), .B(D13769_Y));
KC_AOI211_X1 D13658 ( .A(D14072_Y), .Y(D13658_Y), .C1(D14249_Y),     .C0(D14859_Y), .B(D13691_Y));
KC_AOI211_X1 D13657 ( .A(D14072_Y), .Y(D13657_Y), .C1(D14220_Y),     .C0(D14859_Y), .B(D2442_Y));
KC_AOI211_X1 D13654 ( .A(D14072_Y), .Y(D13654_Y), .C1(D14220_Y),     .C0(D14786_Y), .B(D13690_Y));
KC_AOI211_X1 D13653 ( .A(D14072_Y), .Y(D13653_Y), .C1(D14250_Y),     .C0(D14859_Y), .B(D13689_Y));
KC_AOI211_X1 D13652 ( .A(D14072_Y), .Y(D13652_Y), .C1(D14250_Y),     .C0(D14786_Y), .B(D13581_Y));
KC_AOI211_X1 D13651 ( .A(D14072_Y), .Y(D13651_Y), .C1(D984_Y),     .C0(D14786_Y), .B(D2441_Y));
KC_AOI211_X1 D13650 ( .A(D14072_Y), .Y(D13650_Y), .C1(D14249_Y),     .C0(D14786_Y), .B(D13582_Y));
KC_AOI211_X1 D13574 ( .A(D769_Y), .Y(D13574_Y), .C1(D13557_Y),     .C0(D10216_Y), .B(D13592_Y));
KC_AOI211_X1 D13573 ( .A(D13421_Y), .Y(D13573_Y), .C1(D13027_Y),     .C0(D12813_Y), .B(D2371_Y));
KC_AOI211_X1 D13568 ( .A(D769_Y), .Y(D13568_Y), .C1(D13556_Y),     .C0(D14246_Q), .B(D13600_Y));
KC_AOI211_X1 D13564 ( .A(D769_Y), .Y(D13564_Y), .C1(D13550_Y),     .C0(D14241_Q), .B(D13591_Y));
KC_AOI211_X1 D13563 ( .A(D769_Y), .Y(D13563_Y), .C1(D13561_Y),     .C0(D14239_Q), .B(D13597_Y));
KC_AOI211_X1 D13438 ( .A(D13421_Y), .Y(D13438_Y), .C1(D13696_Y),     .C0(D12813_Y), .B(D13467_Y));
KC_AOI211_X1 D13433 ( .A(D769_Y), .Y(D13433_Y), .C1(D13450_Y),     .C0(D926_Q), .B(D13489_Y));
KC_AOI211_X1 D13432 ( .A(D769_Y), .Y(D13432_Y), .C1(D13449_Y),     .C0(D14166_Q), .B(D13496_Y));
KC_AOI211_X1 D13431 ( .A(D13456_Y), .Y(D13431_Y), .C1(D13512_Y),     .C0(D12813_Y), .B(D13421_Y));
KC_AOI211_X1 D13425 ( .A(D14072_Y), .Y(D13425_Y), .C1(D984_Y),     .C0(D14859_Y), .B(D13486_Y));
KC_AOI211_X1 D13424 ( .A(D13421_Y), .Y(D13424_Y), .C1(D13697_Y),     .C0(D12813_Y), .B(D13430_Y));
KC_AOI211_X1 D13415 ( .A(D769_Y), .Y(D13415_Y), .C1(D13422_Y),     .C0(D14167_Q), .B(D13485_Y));
KC_AOI211_X1 D13414 ( .A(D13421_Y), .Y(D13414_Y), .C1(D12970_Y),     .C0(D12813_Y), .B(D12950_Y));
KC_AOI211_X1 D13324 ( .A(D13320_Y), .Y(D13324_Y), .C1(D13332_Y),     .C0(D13376_Y), .B(D16203_Y));
KC_AOI211_X1 D13232 ( .A(D7609_Y), .Y(D13232_Y), .C1(D14043_Y),     .C0(D13243_Y), .B(D13252_Y));
KC_AOI211_X1 D13219 ( .A(D12739_Y), .Y(D13219_Y), .C1(D13380_Y),     .C0(D13323_Y), .B(D16608_Y));
KC_AOI211_X1 D12937 ( .A(D12895_Y), .Y(D12937_Y), .C1(D12889_Y),     .C0(D12894_Y), .B(D13003_Y));
KC_AOI211_X1 D12866 ( .A(D12797_Y), .Y(D12866_Y), .C1(D783_Y),     .C0(D12794_Y), .B(D12855_Q));
KC_AOI211_X1 D12768 ( .A(D12712_Y), .Y(D12768_Y), .C1(D12769_Y),     .C0(D13349_Y), .B(D12735_Y));
KC_AOI211_X1 D12766 ( .A(D12708_Y), .Y(D12766_Y), .C1(D12767_Y),     .C0(D12732_Y), .B(D12735_Y));
KC_AOI211_X1 D12697 ( .A(D12765_Y), .Y(D12697_Y), .C1(D12204_Y),     .C0(D12717_Y), .B(D12728_Y));
KC_AOI211_X1 D12623 ( .A(D13154_Y), .Y(D12623_Y), .C1(D12631_Y),     .C0(D13287_Y), .B(D12624_Y));
KC_AOI211_X1 D12298 ( .A(D14806_Y), .Y(D12298_Y), .C1(D12299_Y),     .C0(D12203_Y), .B(D12190_Y));
KC_AOI211_X1 D11677 ( .A(D10179_Y), .Y(D11677_Y), .C1(D11678_Y),     .C0(D553_Y), .B(D4747_Y));
KC_AOI211_X1 D10101 ( .A(D10085_Y), .Y(D10101_Y), .C1(D10102_Y),     .C0(D10073_Y), .B(D10067_Y));
KC_AOI211_X1 D10065 ( .A(D10059_Q), .Y(D10065_Y), .C1(D10066_Y),     .C0(D11114_Y), .B(D10054_Y));
KC_AOI211_X1 D9420 ( .A(D9418_Y), .Y(D9420_Y), .C1(D9463_Y),     .C0(D9484_Y), .B(D9408_Y));
KC_AOI211_X1 D9396 ( .A(D9441_Y), .Y(D9396_Y), .C1(D8151_Q),     .C0(D9404_Y), .B(D1989_Y));
KC_AOI211_X1 D9389 ( .A(D9442_Y), .Y(D9389_Y), .C1(D8151_Q),     .C0(D9390_Y), .B(D2062_Y));
KC_AOI211_X1 D9110 ( .A(D9111_Y), .Y(D9110_Y), .C1(D5966_Y),     .C0(D386_Q), .B(D1903_Y));
KC_AOI211_X1 D9100 ( .A(D9106_Y), .Y(D9100_Y), .C1(D6075_Y),     .C0(D12305_Y), .B(D1903_Y));
KC_AOI211_X1 D59 ( .A(D2064_Y), .Y(D59_Y), .C1(D7473_Y), .C0(D8071_Y),     .B(D9055_Y));
KC_AOI211_X1 D9072 ( .A(D9077_Y), .Y(D9072_Y), .C1(D9163_Q),     .C0(D1864_Y), .B(D2012_Y));
KC_AOI211_X1 D9065 ( .A(D9079_Y), .Y(D9065_Y), .C1(D2095_Y),     .C0(D7362_Y), .B(D2047_Y));
KC_AOI211_X1 D9064 ( .A(D9069_Y), .Y(D9064_Y), .C1(D7473_Y),     .C0(D7959_Y), .B(D9066_Y));
KC_AOI211_X1 D9058 ( .A(D8942_Y), .Y(D9058_Y), .C1(D9068_Y),     .C0(D9178_Y), .B(D9083_Y));
KC_AOI211_X1 D9053 ( .A(D8994_Y), .Y(D9053_Y), .C1(D9068_Y),     .C0(D9334_Y), .B(D2046_Y));
KC_AOI211_X1 D9052 ( .A(D9076_Y), .Y(D9052_Y), .C1(D9068_Y),     .C0(D9155_Y), .B(D9082_Y));
KC_AOI211_X1 D9045 ( .A(D9075_Y), .Y(D9045_Y), .C1(D9068_Y),     .C0(D9202_Y), .B(D9050_Y));
KC_AOI211_X1 D9039 ( .A(D8881_Y), .Y(D9039_Y), .C1(D9068_Y),     .C0(D9332_Y), .B(D9093_Y));
KC_AOI211_X1 D8968 ( .A(D1707_Y), .Y(D8968_Y), .C1(D8974_Y),     .C0(D1476_Y), .B(D9042_Y));
KC_AOI211_X1 D8739 ( .A(D9958_Y), .Y(D8739_Y), .C1(D8821_Q),     .C0(D201_Y), .B(D9957_Y));
KC_AOI211_X1 D8673 ( .A(D190_Y), .Y(D8673_Y), .C1(D7132_Y),     .C0(D7133_Y), .B(D8690_Y));
KC_AOI211_X1 D8397 ( .A(D8476_Y), .Y(D8397_Y), .C1(D8382_Y),     .C0(D8384_Y), .B(D8449_Y));
KC_AOI211_X1 D8194 ( .A(D8250_Q), .Y(D8194_Y), .C1(D7655_Y),     .C0(D9528_Y), .B(D9525_Y));
KC_AOI211_X1 D8089 ( .A(D8088_Y), .Y(D8089_Y), .C1(D1984_Y),     .C0(D8153_Y), .B(D642_Y));
KC_AOI211_X1 D7987 ( .A(D7915_Y), .Y(D7987_Y), .C1(D7988_Y),     .C0(D7926_Y), .B(D7921_Y));
KC_AOI211_X1 D7931 ( .A(D1852_Y), .Y(D7931_Y), .C1(D7948_Y),     .C0(D7947_Y), .B(D7916_Y));
KC_AOI211_X1 D7840 ( .A(D6434_Y), .Y(D7840_Y), .C1(D7827_Y),     .C0(D7839_Y), .B(D7916_Y));
KC_AOI211_X1 D7836 ( .A(D1852_Y), .Y(D7836_Y), .C1(D7850_Y),     .C0(D7863_Y), .B(D7837_Y));
KC_AOI211_X1 D7825 ( .A(D7828_Y), .Y(D7825_Y), .C1(D7929_Y),     .C0(D8257_Y), .B(D1857_Y));
KC_AOI211_X1 D7770 ( .A(D7769_Y), .Y(D7770_Y), .C1(D272_Y),     .C0(D7768_Y), .B(D7760_Y));
KC_AOI211_X1 D7681 ( .A(D7721_Y), .Y(D7681_Y), .C1(D7713_Y),     .C0(D6350_Q), .B(D7705_Y));
KC_AOI211_X1 D7632 ( .A(D12305_Y), .Y(D7632_Y), .C1(D7677_Y),     .C0(D6095_Y), .B(D382_Y));
KC_AOI211_X1 D7354 ( .A(D7356_Y), .Y(D7354_Y), .C1(D5671_Y),     .C0(D7369_Y), .B(D5892_Y));
KC_AOI211_X1 D7341 ( .A(D7192_Y), .Y(D7341_Y), .C1(D7338_Y),     .C0(D7385_Y), .B(D5849_Y));
KC_AOI211_X1 D7340 ( .A(D7348_Y), .Y(D7340_Y), .C1(D249_Y),     .C0(D7094_Y), .B(D7233_Y));
KC_AOI211_X1 D7336 ( .A(D4311_Y), .Y(D7336_Y), .C1(D7225_Y),     .C0(D8841_Y), .B(D7352_Y));
KC_AOI211_X1 D7330 ( .A(D7335_Y), .Y(D7330_Y), .C1(D7382_Y),     .C0(D5908_Y), .B(D583_Co));
KC_AOI211_X1 D7312 ( .A(D5936_Y), .Y(D7312_Y), .C1(D9482_Y),     .C0(D7342_Y), .B(D7393_Y));
KC_AOI211_X1 D7309 ( .A(D7224_Y), .Y(D7309_Y), .C1(D7634_Y),     .C0(D7226_Y), .B(D1885_Y));
KC_AOI211_X1 D7230 ( .A(D7376_Y), .Y(D7230_Y), .C1(D7248_Y),     .C0(D7231_Y), .B(D7304_Y));
KC_AOI211_X1 D7223 ( .A(D5760_Y), .Y(D7223_Y), .C1(D8899_Q),     .C0(D4171_Y), .B(D5795_Y));
KC_AOI211_X1 D7222 ( .A(D7187_Y), .Y(D7222_Y), .C1(D7476_Q),     .C0(D7276_Y), .B(D7224_Y));
KC_AOI211_X1 D7202 ( .A(D7179_Y), .Y(D7202_Y), .C1(D7634_Y),     .C0(D220_Y), .B(D7198_Y));
KC_AOI211_X1 D6510 ( .A(D6512_Y), .Y(D6510_Y), .C1(D6555_Q),     .C0(D6514_Y), .B(D6511_Y));
KC_AOI211_X1 D6442 ( .A(D6458_Y), .Y(D6442_Y), .C1(D4900_Y),     .C0(D6445_Y), .B(D6464_Y));
KC_AOI211_X1 D6440 ( .A(D6433_Y), .Y(D6440_Y), .C1(D485_Q),     .C0(D6481_Q), .B(D6444_Y));
KC_AOI211_X1 D6435 ( .A(D6483_Y), .Y(D6435_Y), .C1(D3408_Y),     .C0(D4885_Y), .B(D475_Y));
KC_AOI211_X1 D6425 ( .A(D6458_Y), .Y(D6425_Y), .C1(D4885_Y),     .C0(D6430_Y), .B(D4989_Y));
KC_AOI211_X1 D6424 ( .A(D1852_Y), .Y(D6424_Y), .C1(D7920_Y),     .C0(D6555_Q), .B(D7841_Y));
KC_AOI211_X1 D6366 ( .A(D4951_Y), .Y(D6366_Y), .C1(D446_Q),     .C0(D6365_Y), .B(D6367_Y));
KC_AOI211_X1 D6224 ( .A(D6263_Y), .Y(D6224_Y), .C1(D6254_Y),     .C0(D6247_Y), .B(D6280_Y));
KC_AOI211_X1 D6088 ( .A(D6105_Y), .Y(D6088_Y), .C1(D6500_Y),     .C0(D6106_Y), .B(D16143_Y));
KC_AOI211_X1 D6015 ( .A(D6018_Y), .Y(D6015_Y), .C1(D4243_Y),     .C0(D6017_Y), .B(D6052_Y));
KC_AOI211_X1 D5994 ( .A(D6067_Y), .Y(D5994_Y), .C1(D6000_Y),     .C0(D284_Y), .B(D6053_Y));
KC_AOI211_X1 D5993 ( .A(D213_Y), .Y(D5993_Y), .C1(D5984_Y),     .C0(D5745_Y), .B(D6067_Y));
KC_AOI211_X1 D5979 ( .A(D6046_Y), .Y(D5979_Y), .C1(D7295_Y),     .C0(D6023_Y), .B(D5972_Y));
KC_AOI211_X1 D5946 ( .A(D5741_Y), .Y(D5946_Y), .C1(D5947_Y),     .C0(D7305_Y), .B(D6059_Y));
KC_AOI211_X1 D5945 ( .A(D1908_Y), .Y(D5945_Y), .C1(D6033_Y),     .C0(D6029_Y), .B(D5861_Y));
KC_AOI211_X1 D5891 ( .A(D5858_Y), .Y(D5891_Y), .C1(D7360_Y),     .C0(D7192_Y), .B(D5873_Y));
KC_AOI211_X1 D5879 ( .A(D1727_Y), .Y(D5879_Y), .C1(D6033_Y),     .C0(D5887_Y), .B(D1816_Y));
KC_AOI211_X1 D5860 ( .A(D1727_Y), .Y(D5860_Y), .C1(D5738_Y),     .C0(D5922_Y), .B(D1737_Y));
KC_AOI211_X1 D5844 ( .A(D5845_Y), .Y(D5844_Y), .C1(D6033_Y),     .C0(D1750_Y), .B(D5862_Y));
KC_AOI211_X1 D5843 ( .A(D7386_Y), .Y(D5843_Y), .C1(D7470_Y),     .C0(D7366_Y), .B(D5910_Y));
KC_AOI211_X1 D5836 ( .A(D5829_Y), .Y(D5836_Y), .C1(D5841_Y),     .C0(D7103_Y), .B(D5921_Y));
KC_AOI211_X1 D5824 ( .A(D5714_Y), .Y(D5824_Y), .C1(D9481_Y),     .C0(D7193_Y), .B(D5821_Y));
KC_AOI211_X1 D5767 ( .A(D5714_Y), .Y(D5767_Y), .C1(D5882_Y),     .C0(D4131_Y), .B(D7220_Y));
KC_AOI211_X1 D5766 ( .A(D5717_Y), .Y(D5766_Y), .C1(D4132_Y),     .C0(D5787_Y), .B(D5790_Y));
KC_AOI211_X1 D5759 ( .A(D5716_Y), .Y(D5759_Y), .C1(D8824_Q),     .C0(D4171_Y), .B(D5778_Y));
KC_AOI211_X1 D5758 ( .A(D1728_Y), .Y(D5758_Y), .C1(D6039_Y),     .C0(D4382_Y), .B(D5788_Y));
KC_AOI211_X1 D5748 ( .A(D5779_Y), .Y(D5748_Y), .C1(D177_Y),     .C0(D7373_Y), .B(D5780_Y));
KC_AOI211_X1 D5734 ( .A(D7207_Y), .Y(D5734_Y), .C1(D5698_Y),     .C0(D4353_Y), .B(D5735_Y));
KC_AOI211_X1 D5711 ( .A(D5777_Y), .Y(D5711_Y), .C1(D5646_Y),     .C0(D5755_Y), .B(D5820_Y));
KC_AOI211_X1 D5027 ( .A(D5059_Y), .Y(D5027_Y), .C1(D4883_Y),     .C0(D3582_Y), .B(D4861_Y));
KC_AOI211_X1 D5026 ( .A(D5061_Y), .Y(D5026_Y), .C1(D1562_Y),     .C0(D3416_Y), .B(D5065_Y));
KC_AOI211_X1 D5015 ( .A(D5061_Y), .Y(D5015_Y), .C1(D5028_Y),     .C0(D1562_Y), .B(D5016_Y));
KC_AOI211_X1 D4988 ( .A(D5053_Y), .Y(D4988_Y), .C1(D5033_Y),     .C0(D6449_Y), .B(D5080_Y));
KC_AOI211_X1 D4987 ( .A(D5010_Y), .Y(D4987_Y), .C1(D3484_Q),     .C0(D5056_Y), .B(D4931_Y));
KC_AOI211_X1 D4870 ( .A(D4950_Y), .Y(D4870_Y), .C1(D3400_Y),     .C0(D4978_Y), .B(D4980_Y));
KC_AOI211_X1 D4769 ( .A(D4785_Y), .Y(D4769_Y), .C1(D4698_Y),     .C0(D4779_Y), .B(D6329_Y));
KC_AOI211_X1 D4744 ( .A(D4662_Y), .Y(D4744_Y), .C1(D4745_Y),     .C0(D3302_Q), .B(D4663_Y));
KC_AOI211_X1 D4688 ( .A(D4574_Y), .Y(D4688_Y), .C1(D4694_Y),     .C0(D4575_Y), .B(D4690_Y));
KC_AOI211_X1 D4674 ( .A(D4680_Y), .Y(D4674_Y), .C1(D4670_Y),     .C0(D4724_Y), .B(D92_Y));
KC_AOI211_X1 D4600 ( .A(D47_Y), .Y(D4600_Y), .C1(D4604_Y), .C0(D371_Y),     .B(D50_Y));
KC_AOI211_X1 D4584 ( .A(D4650_Y), .Y(D4584_Y), .C1(D4581_Y),     .C0(D4586_Y), .B(D4594_Y));
KC_AOI211_X1 D4583 ( .A(D4650_Y), .Y(D4583_Y), .C1(D1574_Y),     .C0(D4582_Y), .B(D4588_Y));
KC_AOI211_X1 D4577 ( .A(D4637_Q), .Y(D4577_Y), .C1(D4640_Q),     .C0(D4638_Q), .B(D4582_Y));
KC_AOI211_X1 D4514 ( .A(D4466_Y), .Y(D4514_Y), .C1(D4513_Y),     .C0(D4411_Y), .B(D4481_Y));
KC_AOI211_X1 D4407 ( .A(D4450_Y), .Y(D4407_Y), .C1(D4234_Y),     .C0(D4389_Y), .B(D4404_Y));
KC_AOI211_X1 D4403 ( .A(D4288_Y), .Y(D4403_Y), .C1(D5837_Y),     .C0(D4291_Y), .B(D5853_Y));
KC_AOI211_X1 D4352 ( .A(D4373_Y), .Y(D4352_Y), .C1(D7243_Y),     .C0(D249_Y), .B(D4384_Y));
KC_AOI211_X1 D4332 ( .A(D5928_Y), .Y(D4332_Y), .C1(D4345_Y),     .C0(D4327_Y), .B(D4331_Y));
KC_AOI211_X1 D4321 ( .A(D4393_Y), .Y(D4321_Y), .C1(D5863_Y),     .C0(D4333_Y), .B(D5911_Y));
KC_AOI211_X1 D4297 ( .A(D5833_Y), .Y(D4297_Y), .C1(D4299_Y),     .C0(D4317_Y), .B(D4365_Y));
KC_AOI211_X1 D4296 ( .A(D4311_Y), .Y(D4296_Y), .C1(D8865_Y),     .C0(D7164_Y), .B(D4314_Y));
KC_AOI211_X1 D4295 ( .A(D4414_Y), .Y(D4295_Y), .C1(D3038_Y),     .C0(D4306_Y), .B(D8861_Y));
KC_AOI211_X1 D4286 ( .A(D7315_Y), .Y(D4286_Y), .C1(D3038_Y),     .C0(D5833_Y), .B(D4364_Y));
KC_AOI211_X1 D4273 ( .A(D5833_Y), .Y(D4273_Y), .C1(D4465_Y),     .C0(D4299_Y), .B(D5936_Y));
KC_AOI211_X1 D3601 ( .A(D1953_Y), .Y(D3601_Y), .C1(D3646_Q),     .C0(D1474_Y), .B(D3600_Y));
KC_AOI211_X1 D3530 ( .A(D3553_Y), .Y(D3530_Y), .C1(D3406_Y),     .C0(D4916_Y), .B(D3409_Y));
KC_AOI211_X1 D3518 ( .A(D3578_Y), .Y(D3518_Y), .C1(D3531_Y),     .C0(D3527_Y), .B(D3547_Y));
KC_AOI211_X1 D3506 ( .A(D3578_Y), .Y(D3506_Y), .C1(D3531_Y),     .C0(D3522_Y), .B(D3557_Y));
KC_AOI211_X1 D3496 ( .A(D68_Y), .Y(D3496_Y), .C1(D3497_Y),     .C0(D4926_Y), .B(D4911_Y));
KC_AOI211_X1 D3495 ( .A(D3496_Y), .Y(D3495_Y), .C1(D4891_Y),     .C0(D4969_Y), .B(D3450_Y));
KC_AOI211_X1 D3435 ( .A(D3411_Y), .Y(D3435_Y), .C1(D3432_Y),     .C0(D3488_Y), .B(D4939_Y));
KC_AOI211_X1 D3434 ( .A(D3439_Y), .Y(D3434_Y), .C1(D3372_Q),     .C0(D5033_Y), .B(D3474_Y));
KC_AOI211_X1 D3397 ( .A(D1453_Y), .Y(D3397_Y), .C1(D3346_Y),     .C0(D4815_Y), .B(D3362_Y));
KC_AOI211_X1 D3310 ( .A(D3396_Y), .Y(D3310_Y), .C1(D3337_Y),     .C0(D3313_Y), .B(D3312_Y));
KC_AOI211_X1 D3300 ( .A(D3327_Y), .Y(D3300_Y), .C1(D3301_Y),     .C0(D3258_Y), .B(D3246_Y));
KC_AOI211_X1 D3236 ( .A(D1423_Y), .Y(D3236_Y), .C1(D3283_Q),     .C0(D1425_Y), .B(D3238_Y));
KC_AOI211_X1 D3211 ( .A(D3277_Y), .Y(D3211_Y), .C1(D3261_Y),     .C0(D4815_Y), .B(D3213_Y));
KC_AOI211_X1 D3199 ( .A(D3113_Y), .Y(D3199_Y), .C1(D3200_Y),     .C0(D3194_Y), .B(D3125_Y));
KC_AOI211_X1 D3197 ( .A(D3125_Y), .Y(D3197_Y), .C1(D3198_Y),     .C0(D3165_Y), .B(D3131_Y));
KC_AOI211_X1 D3121 ( .A(D3123_Y), .Y(D3121_Y), .C1(D3122_Y),     .C0(D3123_Y), .B(D3123_Y));
KC_AOI211_X1 D3111 ( .A(D3172_Y), .Y(D3111_Y), .C1(D3165_Y),     .C0(D3048_Y), .B(D7641_Y));
KC_AOI211_X1 D3110 ( .A(D3172_Y), .Y(D3110_Y), .C1(D3108_Y),     .C0(D3252_Y), .B(D3120_Y));
KC_AOI211_X1 D3103 ( .A(D3128_Y), .Y(D3103_Y), .C1(D3252_Y),     .C0(D3108_Y), .B(D3107_Y));
KC_AOI211_X1 D3102 ( .A(D1421_Y), .Y(D3102_Y), .C1(D4592_Y),     .C0(D3165_Y), .B(D3157_Y));
KC_AOI211_X1 D3100 ( .A(D3157_Y), .Y(D3100_Y), .C1(D4773_Y),     .C0(D3194_Y), .B(D4575_Y));
KC_AOI211_X1 D3095 ( .A(D345_Y), .Y(D3095_Y), .C1(D3061_Y),     .C0(D3167_Y), .B(D3104_Y));
KC_AOI211_X1 D2903 ( .A(D2955_Y), .Y(D2903_Y), .C1(D2952_Y),     .C0(D2996_Y), .B(D28_Y));
KC_AOI211_X1 D2841 ( .A(D2843_Y), .Y(D2841_Y), .C1(D2847_Y),     .C0(D2839_Y), .B(D2804_Y));
KC_AOI211_X1 D2840 ( .A(D2804_Y), .Y(D2840_Y), .C1(D2888_Q),     .C0(D2843_Y), .B(D2842_Y));
KC_AOI211_X1 D2759 ( .A(D2764_Y), .Y(D2759_Y), .C1(D1441_Y),     .C0(D2848_Y), .B(D2757_Y));
KC_AOI211_X1 D2754 ( .A(D2755_Y), .Y(D2754_Y), .C1(D2801_Q),     .C0(D2886_Q), .B(D2756_Y));
KC_AOI211_X1 D2748 ( .A(D1442_Y), .Y(D2748_Y), .C1(D2750_Y),     .C0(D2754_Y), .B(D2749_Y));
KC_AOI211_X1 D2743 ( .A(D2772_Y), .Y(D2743_Y), .C1(D2783_Y),     .C0(D2901_Y), .B(D2801_Q));
KC_AOI211_X1 D2611 ( .A(D15545_Y), .Y(D2611_Y), .C1(D15485_Y),     .C0(D15657_Y), .B(D15546_Y));
KC_AOI211_X1 D2592 ( .A(D15405_Y), .Y(D2592_Y), .C1(D16047_Y),     .C0(D2593_Y), .B(D15406_Y));
KC_AOI211_X1 D2423 ( .A(D769_Y), .Y(D2423_Y), .C1(D2428_Y),     .C0(D14164_Q), .B(D2445_Y));
KC_AOI211_X1 D2422 ( .A(D13421_Y), .Y(D2422_Y), .C1(D13699_Y),     .C0(D12813_Y), .B(D2401_Y));
KC_AOI211_X1 D1970 ( .A(D7172_Y), .Y(D1970_Y), .C1(D1971_Y),     .C0(D355_Y), .B(D1910_Y));
KC_AOI211_X1 D1867 ( .A(D1868_Y), .Y(D1867_Y), .C1(D1870_Y),     .C0(D1952_Y), .B(D7511_Y));
KC_AOI211_X1 D1862 ( .A(D18_Y), .Y(D1862_Y), .C1(D7631_Y),     .C0(D5981_Y), .B(D382_Y));
KC_AOI211_X1 D1850 ( .A(D7839_Y), .Y(D1850_Y), .C1(D7946_Y),     .C0(D7955_Y), .B(D7924_Y));
KC_AOI211_X1 D1826 ( .A(D1966_Y), .Y(D1826_Y), .C1(D1935_Y),     .C0(D1828_Y), .B(D105_Y));
KC_AOI211_X1 D1725 ( .A(D7192_Y), .Y(D1725_Y), .C1(D291_Y),     .C0(D1728_Y), .B(D1768_Y));
KC_AOI211_X1 D1715 ( .A(D1723_Y), .Y(D1715_Y), .C1(D6026_Y),     .C0(D240_Y), .B(D1752_Y));
KC_AOI211_X1 D1693 ( .A(D7974_Y), .Y(D1693_Y), .C1(D6426_Y),     .C0(D468_Y), .B(D1820_Y));
KC_AOI211_X1 D1589 ( .A(D4402_Y), .Y(D1589_Y), .C1(D4356_Y),     .C0(D4245_Y), .B(D1616_Y));
KC_AOI211_X1 D1588 ( .A(D1627_Y), .Y(D1588_Y), .C1(D4172_Y),     .C0(D4119_Q), .B(D4313_Y));
KC_AOI211_X1 D1561 ( .A(D1415_Y), .Y(D1561_Y), .C1(D5012_Y),     .C0(D3599_Y), .B(D3413_Y));
KC_AOI211_X1 D1532 ( .A(D1443_Y), .Y(D1532_Y), .C1(D1533_Y),     .C0(D3527_Y), .B(D3457_Y));
KC_AOI211_X1 D1420 ( .A(D1422_Y), .Y(D1420_Y), .C1(D1426_Y),     .C0(D3237_Y), .B(D1423_Y));
KC_AOI211_X1 D1418 ( .A(D1480_Y), .Y(D1418_Y), .C1(D1506_Y),     .C0(D3265_Y), .B(D3288_Y));
KC_AOI211_X1 D1416 ( .A(D3484_Q), .Y(D1416_Y), .C1(D4925_Y),     .C0(D1451_Y), .B(D1467_Y));
KC_AOI211_X1 D1414 ( .A(D3455_Y), .Y(D1414_Y), .C1(D1562_Y),     .C0(D1448_Y), .B(D3490_Y));
KC_AOI211_X1 D1405 ( .A(D16530_Y), .Y(D1405_Y), .C1(D16482_Y),     .C0(D16511_Y), .B(D13392_Y));
KC_AOI211_X1 D1182 ( .A(D14334_Y), .Y(D1182_Y), .C1(D13761_Q),     .C0(D13719_Y), .B(D13746_Y));
KC_AOI211_X1 D751 ( .A(D14762_Y), .Y(D751_Y), .C1(D15483_Y),     .C0(D14867_Y), .B(D15542_Y));
KC_AOI211_X1 D641 ( .A(D14656_Y), .Y(D641_Y), .C1(D15395_Y),     .C0(D14656_Y), .B(D2565_Y));
KC_AOI211_X1 D634 ( .A(D14660_Y), .Y(D634_Y), .C1(D15350_Y),     .C0(D771_Y), .B(D15413_Y));
KC_AOI211_X1 D624 ( .A(D9418_Y), .Y(D624_Y), .C1(D10214_Y),     .C0(D10310_Y), .B(D10195_Y));
KC_AOI211_X1 D552 ( .A(D2379_Y), .Y(D552_Y), .C1(D161_Y),     .C0(D12661_Y), .B(D12663_Y));
KC_AOI211_X1 D494 ( .A(D7919_Y), .Y(D494_Y), .C1(D6426_Y),     .C0(D4982_Y), .B(D7918_Y));
KC_AOI211_X1 D470 ( .A(D5008_Y), .Y(D470_Y), .C1(D1563_Y),     .C0(D4996_Y), .B(D5072_Y));
KC_AOI211_X1 D467 ( .A(D1858_Y), .Y(D467_Y), .C1(D7935_Y),     .C0(D6421_Y), .B(D7952_Y));
KC_AOI211_X1 D433 ( .A(D436_Y), .Y(D433_Y), .C1(D432_Y), .C0(D4906_Y),     .B(D1449_Y));
KC_AOI211_X1 D406 ( .A(D4662_Y), .Y(D406_Y), .C1(D3298_Y),     .C0(D4763_Y), .B(D3381_Y));
KC_AOI211_X1 D398 ( .A(D3248_Y), .Y(D398_Y), .C1(D397_Y), .C0(D3298_Y),     .B(D3327_Y));
KC_AOI211_X1 D341 ( .A(D1945_Y), .Y(D341_Y), .C1(D4629_Y), .C0(D166_Y),     .B(D4593_Y));
KC_AOI211_X1 D269 ( .A(D7356_Y), .Y(D269_Y), .C1(D7348_Y),     .C0(D5768_Y), .B(D7343_Y));
KC_AOI211_X1 D246 ( .A(D93_Y), .Y(D246_Y), .C1(D4243_Y), .C0(D260_Y),     .B(D4379_Y));
KC_AOI211_X1 D241 ( .A(D93_Y), .Y(D241_Y), .C1(D240_Y), .C0(D280_Y),     .B(D4376_Y));
KC_AOI211_X1 D206 ( .A(D7195_Y), .Y(D206_Y), .C1(D7193_Y), .C0(D214_Y),     .B(D1737_Y));
KC_AOI211_X1 D200 ( .A(D7263_Y), .Y(D200_Y), .C1(D5881_Y),     .C0(D3573_Y), .B(D4221_Y));
KC_AOI211_X1 D170 ( .A(D13421_Y), .Y(D170_Y), .C1(D13028_Y),     .C0(D12813_Y), .B(D2372_Y));
KC_AOI211_X1 D76 ( .A(D1883_Y), .Y(D76_Y), .C1(D5671_Y), .C0(D7395_Y),     .B(D5940_Y));
KC_AOI211_X1 D75 ( .A(D6071_Y), .Y(D75_Y), .C1(D7263_Y), .C0(D291_Y),     .B(D6055_Y));
KC_AOI211_X1 D61 ( .A(D8671_Y), .Y(D61_Y), .C1(D8759_Y), .C0(D1977_Y),     .B(D8717_Y));

endmodule
