// Library - lyt_9160734, Cell - lyt, View - schematic
// LAST TIME SAVED: Feb  4 16:06:55 2017
// NETLIST TIME: Feb  4 16:07:23 2017
`timescale 1ns / 1ns 

module lyt_top (
T13053_SN,
T9218_B  ,
T15168_CK,
T9484_B  ,
T9495_B  ,
T9496_B  ,
T9493_B  ,
T9494_B  ,
T2377_A  ,
T2378_A  ,
T1845_A  ,
T1835_A  ,
T1855_A  ,
T15190_A ,
T15167_A ,
T1283_RN ,
T209_A   ,
T15004_A ,
T9198_B  ,
T9197_B  ,
T9214_B  ,
T9215_B  ,
T9216_B  ,
T9217_B  ,
T9209_B  ,
T9210_B  ,
T9211_B  ,
T9212_B  ,
T9213_B  ,
T9237_B  ,
T9236_B  ,
T9238_B  ,
T9250_B  ,
T9248_B  ,
T9206_B  ,
T9207_B  ,
T9205_B  ,
T9201_B  ,
T9208_B  ,
T9203_B  ,
T9204_B  ,
T9202_B  ,
T9249_B  ,
T9134_B  ,
T9499_B  ,
T9492_B  ,
T9491_B  ,
T9183_B  ,
T9084_B  ,
T9083_B  ,
T9179_B  ,
T238_AN  ,    //up input  
T5422_Y  ,
T16170_Y ,
T4929_Y  ,
T4879_Y  ,
T2075_Y  ,
T1851_Y  ,
T1853_Y  ,
T1852_Y  ,
T1854_Y  ,
T1848_Y  ,
T1849_Y  ,
T15717_Y ,
T15716_Y ,
T6497_Y  ,
T15925_Y ,
T1754_Y  ,
T1756_Y  ,
T1755_Y  ,
T1747_Y  ,
T1745_Y  ,
T845_Y   ,
T1616_Y  ,
T1170_Y  ,
T1169_Y  ,
T1145_Y  ,
T213_Y   ,
T1023_Y  ,
T1024_Y  ,
T586_Y   ,
T593_Y   ,
T11900_Y ,
T16188_Y ,
T141_Q   ,
T13264_Y ,
T429_Y   ,
T428_Y   ,
T395_Y   ,
T199_Y   ,
T15718_Y ,
T16487_Q ,
T16488_Q ,
T16483_Q ,
T16486_Q ,
T2091_Q  ,
T16485_Q ,
T2125_Y  ,
T5443_Y  ,
T1746_Y  ,
T1006_Y  ,
T4409_Y  ,
T211_Q   ,
T6359_Q  ,
T6417_Q  ,
T6730_Q  ,
T6425_Q  ,
T6364_Q  ,
T6432_Q  ,
T6361_Q  ,
T6415_Q  ,
T6423_Q  ,
T6371_Q  ,
T6479_Q  ,
T6358_Q  ,
T6424_Q  ,
T6391_Q  ,
T7899_Y  ,
T7815_Y  ,
T7811_Y  ,
T7853_Y  ,
T7854_Y  ,
T7859_Y  ,
T7809_Y  ,
T16480_Q ,
T152_Y


  );
input  T13053_SN;
input  T9218_B  ;
input  T15168_CK;
input  T9484_B  ;
input  T9495_B  ;
input  T9496_B  ;
input  T9493_B  ;
input  T9494_B  ;
input  T2377_A  ;
input  T2378_A  ;
input  T1845_A  ;
input  T1835_A  ;
input  T1855_A  ;
input  T15190_A ;
input  T15167_A ;
input  T1283_RN ;
input  T209_A   ;
input  T15004_A ;
input  T9198_B  ;
input  T9197_B  ;
input  T9214_B  ;
input  T9215_B  ;
input  T9216_B  ;
input  T9217_B  ;
input  T9209_B  ;
input  T9210_B  ;
input  T9211_B  ;
input  T9212_B  ;
input  T9213_B  ;
input  T9237_B  ;
input  T9236_B  ;
input  T9238_B  ;
input  T9250_B  ;
input  T9248_B  ;
input  T9206_B  ;
input  T9207_B  ;
input  T9205_B  ;
input  T9201_B  ;
input  T9208_B  ;
input  T9203_B  ;
input  T9204_B  ;
input  T9202_B  ;
input  T9249_B  ;
input  T9134_B  ;
input  T9499_B  ;
input  T9492_B  ;
input  T9491_B  ;
input  T9183_B  ;
input  T9084_B  ;
input  T9083_B  ;
input  T9179_B  ;
input  T238_AN  ;    //up input  
output T5422_Y  ;
output T16170_Y ;
output T4929_Y  ;
output T4879_Y  ;
output T2075_Y  ;
output T1851_Y  ;
output T1853_Y  ;
output T1852_Y  ;
output T1854_Y  ;
output T1848_Y  ;
output T1849_Y  ;
output T15717_Y ;
output T15716_Y ;
output T6497_Y  ;
output T15925_Y ;
output T1754_Y  ;
output T1756_Y  ;
output T1755_Y  ;
output T1747_Y  ;
output T1745_Y  ;
output T845_Y   ;
output T1616_Y  ;
output T1170_Y  ;
output T1169_Y  ;
output T1145_Y  ;
output T213_Y   ;
output T1023_Y  ;
output T1024_Y  ;
output T586_Y   ;
output T593_Y   ;
output T11900_Y ;
output T16188_Y ;
output T141_Q   ;
output T13264_Y ;
output T429_Y   ;
output T428_Y   ;
output T395_Y   ;
output T199_Y   ;
output T15718_Y ;  ////
output T16487_Q ;
output T16488_Q ;
output T16483_Q ;
output T16486_Q ;
output T2091_Q  ;
output T16485_Q ;
output T2125_Y  ;
output T5443_Y  ;
output T1746_Y  ;
output T1006_Y  ;
output T4409_Y  ;
output T211_Q   ;
output T6359_Q  ;
output T6417_Q  ;
output T6730_Q  ;
output T6425_Q  ;
output T6364_Q  ;
output T6432_Q  ;
output T6361_Q  ;
output T6415_Q  ;
output T6423_Q  ;
output T6371_Q  ;
output T6479_Q  ;
output T6358_Q  ;
output T6424_Q  ;
output T6391_Q  ;
output T7899_Y  ;
output T7815_Y  ;
output T7811_Y  ;
output T7853_Y  ;
output T7854_Y  ;
output T7859_Y  ;
output T7809_Y  ;
output T16480_Q ;
output T152_Y   ;


//specify 
//    specparam CDS_LIBNAME  = "lyt_9160734";
//    specparam CDS_CELLNAME = "lyt";
//    specparam CDS_VIEWNAME = "schematic";
//endspecify


KC_NAND3_X3 T350 ( .Y(T350_Y), .B(T9271_Y), .C(T6318_Y), .A(T8579_Y));
KC_INV_X8 T187 ( .Y(T187_Y), .A(T15407_Y));
KC_OAI21B_X4 T1345 ( .A0N(T11274_Y), .B(T1446_Y), .A1(T8268_Y),     .Y(T1345_Y));
KC_AO2222_X2 T15839 ( .Y(T15839_Y), .A0(T11188_Y), .A1(T8741_Y),     .B0(T8697_Y), .B1(T16320_Y), .C0(T8742_Y), .C1(T9178_Y),     .D0(T8740_Y), .D1(T9333_Y));
KC_AO2222_X2 T736 ( .Y(T736_Y), .A0(T11214_Y), .A1(T8697_Y),     .B0(T11187_Y), .B1(T8741_Y), .C0(T8649_Y), .C1(T8740_Y),     .D0(T8107_Y), .D1(T8742_Y));
KC_AO2222_X2 T16162 ( .Y(T16162_Y), .A0(T682_Y), .A1(T8741_Y),     .B0(T8703_Y), .B1(T8697_Y), .C0(T9020_Y), .C1(T8742_Y),     .D0(T8637_Y), .D1(T8740_Y));
KC_AO2222_X2 T7813 ( .Y(T7813_Y), .A0(T11184_Y), .A1(T8697_Y),     .B0(T11893_Y), .B1(T8741_Y), .C0(T9344_Y), .C1(T8740_Y),     .D0(T8143_Y), .D1(T8742_Y));
KC_AO2222_X2 T7812 ( .Y(T7812_Y), .A0(T11187_Y), .A1(T8697_Y),     .B0(T11184_Y), .B1(T8741_Y), .C0(T8108_Y), .C1(T8742_Y),     .D0(T9511_Y), .D1(T8740_Y));
KC_AO2222_X2 T15840 ( .Y(T15840_Y), .A0(T11247_Y), .A1(T8868_Y),     .B0(T8812_Y), .B1(T12455_Y), .C0(T8867_Y), .C1(T9489_Y),     .D0(T8811_Y), .D1(T8710_Y));
KC_AO2222_X2 T8808 ( .Y(T8808_Y), .A0(T11269_Y), .A1(T8812_Y),     .B0(T11266_Y), .B1(T8868_Y), .C0(T8666_Y), .C1(T8811_Y),     .D0(T9068_Y), .D1(T8867_Y));
KC_AO2222_X2 T16376 ( .Y(T16376_Y), .A0(T11246_Y), .A1(T8812_Y),     .B0(T11269_Y), .B1(T8868_Y), .C0(T9018_Y), .C1(T8867_Y),     .D0(T8646_Y), .D1(T8811_Y));
KC_MXI2B_X1 T15377 ( .Y(T15377_Y), .A(T6855_S), .BN(T433_Y),     .S0(T280_Y));
KC_MXI2B_X1 T10138 ( .Y(T10138_Y), .A(T4917_Y), .BN(T957_Y),     .S0(T9199_Y));
KC_BUF_X15 T10211 ( .Y(T10211_Y), .A(T9472_Q));
KC_OAI112_X2 T16463 ( .A(T8805_Y), .B(T7645_Y), .C0(T15654_Y),     .C1(T7801_Y), .Y(T16463_Y));
KC_AOI22BB_X1 T15771 ( .Y(T15771_Y), .A0N(T7672_Y), .A1(T16332_Y),     .B0N(T7570_Y), .B1(T9375_Y));
KC_AOI22BB_X1 T15764 ( .Y(T15764_Y), .A0N(T7567_Y), .A1(T9375_Y),     .B0N(T7674_Y), .B1(T16332_Y));
KC_AOI22BB_X1 T16389 ( .Y(T16389_Y), .A0N(T7906_Y), .A1(T8948_Y),     .B0N(T7904_Y), .B1(T1213_Y));
KC_AOI22BB_X1 T15791 ( .Y(T15791_Y), .A0N(T7903_Y), .A1(T1213_Y),     .B0N(T7857_Y), .B1(T8948_Y));
KC_AOI22BB_X1 T6815 ( .Y(T6815_Y), .A0N(T155_Q), .A1(T179_Q),     .B0N(T360_Q), .B1(T9338_Q));
KC_AOI22BB_X1 T15768 ( .Y(T15768_Y), .A0N(T529_Q), .A1(T4827_Q),     .B0N(T517_Q), .B1(T4840_Q));
KC_AOI22BB_X1 T15789 ( .Y(T15789_Y), .A0N(T13260_Y), .A1(T8860_Y),     .B0N(T9445_Y), .B1(T8859_Y));
KC_AOI22BB_X1 T15788 ( .Y(T15788_Y), .A0N(T8895_Y), .A1(T8860_Y),     .B0N(T8899_Y), .B1(T8859_Y));
KC_AOI22BB_X1 T15787 ( .Y(T15787_Y), .A0N(T8894_Y), .A1(T8860_Y),     .B0N(T8898_Y), .B1(T8859_Y));
KC_XOR2_X6 T4353 ( .B(T958_Y), .A(T7870_Y), .Y(T4353_Y));
KC_BUF_X12 T213 ( .Y(T213_Y), .A(T13065_Q));
KC_AO22_X3 T16302 ( .B0(T2073_Y), .B1(T10041_Y), .A1(T10160_Y),     .A0(T15800_Y), .Y(T16302_Y));
KC_NAND2B_X2 T6819 ( .B(T7599_Y), .Y(T6819_Y), .AN(T9374_Y));
KC_NAND2B_X2 T16159 ( .B(T1257_Y), .Y(T16159_Y), .AN(T10142_Y));
KC_DFFSNHQ_X4 T13064 ( .Q(T13064_Q), .D(T10227_Y), .CK(T15168_Q),     .SN(T13053_SN));
KC_DFFSNHQ_X4 T13057 ( .Q(T13057_Q), .D(T1377_Y), .CK(T15176_Y),     .SN(T13053_SN));
KC_NOR3_X3 T845 ( .Y(T845_Y), .B(T16407_Y), .C(T2539_Y), .A(T1675_Q));
KC_NOR2B_X5 T3926 ( .B(T15989_Y), .AN(T1789_Q), .Y(T3926_Y));
KC_OAI21B_X3 T8189 ( .BN(T1764_Y), .A0(T1765_Y), .A1(T15941_Y),     .Y(T8189_Y));
KC_NOR2B_X4 T15924 ( .B(T15036_Y), .AN(T1763_Y), .Y(T15924_Y));
KC_AND2BB_X1 T15925 ( .BN(T148_Y), .Y(T15925_Y), .AN(T1764_Y));
KC_AND2BB_X1 T15923 ( .BN(T15036_Y), .Y(T15923_Y), .AN(T1763_Y));
KC_NOR2B_X2 T13088 ( .B(T15904_Y), .AN(T1826_Q), .Y(T13088_Y));
KC_NOR2B_X2 T16150 ( .B(T15989_Y), .AN(T1787_Q), .Y(T16150_Y));
KC_NOR2B_X2 T15921 ( .B(T15989_Y), .AN(T4925_Q), .Y(T15921_Y));
KC_NOR2B_X2 T15920 ( .B(T15989_Y), .AN(T1823_Q), .Y(T15920_Y));
KC_NOR2B_X2 T15914 ( .B(T15989_Y), .AN(T1806_Q), .Y(T15914_Y));
KC_NOR2B_X2 T15905 ( .B(T15989_Y), .AN(T1785_Q), .Y(T15905_Y));
KC_AND2B_X1 T2599 ( .B(T9880_Y), .A(T6686_Co), .Y(T2599_Y));
KC_OR2_X3 T15006 ( .Y(T15006_Y), .A(T8395_Y), .B(T5389_Q));
KC_OR2_X3 T14965 ( .Y(T14965_Y), .A(T2076_Y), .B(T10253_Y));
KC_INV_X5 T14967 ( .Y(T14967_Y), .A(T1855_Y));
KC_NAND3_X5 T16151 ( .Y(T16151_Y), .B(T11416_Y), .C(T11415_Y),     .A(T2165_Y));
KC_AOI21BB_X1 T6556 ( .BN(T2359_Q), .A1N(T8412_Y), .Y(T6556_Y),     .A0(T2355_Q));
KC_MXI2B_X6 T15507 ( .Y(T15507_Y), .A(T2540_Y), .BN(T2523_Y),     .S0(T16169_Y));
KC_MXI2B_X3 T15957 ( .Y(T15957_Y), .B(T8253_Y), .AN(T10088_Y),     .S0(T1773_Y));
KC_MXI2B_X3 T16447 ( .Y(T16447_Y), .B(T10942_Y), .AN(T14501_Q),     .S0(T2640_Q));
KC_OAI211B_X3 T16244 ( .C0N(T16266_Y), .B(T4896_Y), .A(T16264_Y),     .C1(T4868_Y), .Y(T16244_Y));
KC_AO22_X2 T16235 ( .B0(T10203_Y), .B1(T2484_Y), .A1(T12089_Y),     .A0(T16236_Y), .Y(T16235_Y));
KC_AO22_X2 T9162 ( .B0(T10203_Y), .B1(T2455_Y), .A1(T3669_Y),     .A0(T16236_Y), .Y(T9162_Y));
KC_OAI112B_X1 T16164 ( .C0(T2663_Y), .BN(T14984_Y), .A(T16161_Y),     .C1(T2655_Y), .Y(T16164_Y));
KC_NAND3B_X2 T10263 ( .CN(T10275_Y), .Y(T10263_Y), .B(T5750_Y),     .A(T2657_Y));
KC_AOI32_X2 T15786 ( .E(T7855_Y), .B(T7855_Y), .C(T7818_Y),     .Y(T15786_Y), .D(T968_Y), .A(T8138_Y));
KC_AOI32_X2 T6821 ( .E(T7357_Y), .B(T7357_Y), .C(T7418_Y), .Y(T6821_Y),     .D(T886_Y), .A(T11140_Y));
KC_AOI32_X2 T15892 ( .E(T15804_Q), .B(T15804_Q), .C(T5813_Y),     .Y(T15892_Y), .D(T2707_Y), .A(T11432_Y));
KC_XNOR2_X5 T16452 ( .Y(T16452_Y), .A(T11582_Y), .B(T1708_Y));
KC_BUF_X7 T13211 ( .Y(T13211_Y), .A(T15180_Y));
KC_BUF_X7 T13288 ( .Y(T13288_Y), .A(T14983_Y));
KC_BUF_X7 T13262 ( .Y(T13262_Y), .A(T15177_Q));
KC_BUF_X7 T13266 ( .Y(T13266_Y), .A(T15183_Q));
KC_BUF_X7 T13261 ( .Y(T13261_Y), .A(T1510_Y));
KC_BUF_X7 T13268 ( .Y(T13268_Y), .A(T2097_Y));
KC_TINV_X2 T2183 ( .B(T11498_Y), .Y(T2183_Y), .A(T2184_Y));
KC_TINV_X2 T2831 ( .B(T5013_Y), .Y(T2831_Y), .A(T8467_Y));
KC_NAND4_X3 T6334 ( .D(T2823_Y), .C(T12047_Y), .B(T11676_Y),     .A(T6086_Y), .Y(T6334_Y));
KC_OR4_X2 T8395 ( .Y(T8395_Y), .C(T3524_Q), .B(T2839_Y), .D(T10978_Y),     .A(T2949_Q));
KC_OR4_X2 T8394 ( .Y(T8394_Y), .C(T2878_Q), .B(T2949_Q), .D(T16081_Q),     .A(T16458_Q));
KC_OAI211B_X2 T9057 ( .B(T10174_Y), .C0(T10143_Y), .AN(T10069_Y),     .C1(T1257_Y), .Y(T9057_Y));
KC_OAI211B_X2 T16121 ( .B(T6493_Y), .C0(T6077_Y), .AN(T5503_Y),     .C1(T15989_Y), .Y(T16121_Y));
KC_AND4_X2 T16120 ( .D(T10978_Y), .C(T6161_Y), .B(T6159_Y),     .A(T6086_Y), .Y(T16120_Y));
KC_NAND2_X3 T12067 ( .B(T6561_Y), .A(T12065_Y), .Y(T12067_Y));
KC_OAI21BB_X2 T6830 ( .BN(T9412_Y), .A1N(T690_Q), .A0(T7365_Y),     .Y(T6830_Y));
KC_OAI21BB_X2 T16052 ( .BN(T5500_Y), .A1N(T11666_Y), .A0(T11678_Y),     .Y(T16052_Y));
KC_OAI21BB_X2 T15862 ( .BN(T3242_Q), .A1N(T5074_Q), .A0(T12148_Y),     .Y(T15862_Y));
KC_MXI2B_X5 T8268 ( .Y(T8268_Y), .A(T8989_Y), .BN(T15490_Y),     .S0(T15489_Y));
KC_MXI2B_X5 T3352 ( .Y(T3352_Y), .A(T2734_Y), .BN(T2762_Y),     .S0(T2758_Y));
KC_MXI2B_X5 T3345 ( .Y(T3345_Y), .A(T3991_Y), .BN(T6230_Co),     .S0(T3315_Y));
KC_XNOR2_X4 T12461 ( .A(T11397_Y), .B(T10638_Y), .Y(T12461_Y));
KC_XNOR2_X4 T12460 ( .A(T11581_Y), .B(T8286_Y), .Y(T12460_Y));
KC_XNOR2_X4 T12462 ( .A(T8224_Y), .B(T11455_Y), .Y(T12462_Y));
KC_XNOR2_X4 T12463 ( .A(T11561_Y), .B(T13135_Q), .Y(T12463_Y));
KC_AND2B_X2 T4468 ( .B(T8324_Y), .A(T3351_Y), .Y(T4468_Y));
KC_NOR2_X5 T16148 ( .Y(T16148_Y), .A(T15636_Y), .B(T2917_Y));
KC_NOR2_X5 T16156 ( .Y(T16156_Y), .A(T2848_Y), .B(T3411_Y));
KC_NOR3B_X2 T15951 ( .Y(T15951_Y), .B(T5911_Y), .A(T1766_Y),     .CN(T1835_Y));
KC_NOR3B_X2 T16033 ( .Y(T16033_Y), .B(T3385_Y), .A(T3354_Y),     .CN(T12003_Y));
KC_NAND3_X4 T6515 ( .Y(T6515_Y), .B(T3525_Q), .C(T3527_Y),     .A(T3520_Q));
KC_OAI22B_X1 T9099 ( .A1(T9157_Y), .B0(T9156_Y), .A0(T9114_Y),     .B1N(T9124_Y), .Y(T9099_Y));
KC_OAI22B_X1 T16313 ( .A1(T914_Y), .B0(T741_Q), .A0(T528_Q),     .B1N(T714_Q), .Y(T16313_Y));
KC_OAI22B_X1 T16439 ( .A1(T7866_Y), .B0(T12677_Y), .A0(T7868_Y),     .B1N(T5343_Q), .Y(T16439_Y));
KC_OAI22B_X1 T16438 ( .A1(T7869_Y), .B0(T8761_Y), .A0(T7867_Y),     .B1N(T5360_Q), .Y(T16438_Y));
KC_OAI22B_X1 T1696 ( .A1(T7866_Y), .B0(T12678_Y), .A0(T15654_Y),     .B1N(T5359_Q), .Y(T1696_Y));
KC_OAI22B_X1 T16432 ( .A1(T10329_Y), .B0(T8025_Y), .A0(T16377_Y),     .B1N(T1216_Q), .Y(T16432_Y));
KC_OAI22B_X1 T6553 ( .A1(T2339_Y), .B0(T11751_Y), .A0(T6522_Y),     .B1N(T1832_Q), .Y(T6553_Y));
KC_OAI22B_X1 T6544 ( .A1(T2339_Y), .B0(T11046_Y), .A0(T6518_Y),     .B1N(T2364_Q), .Y(T6544_Y));
KC_OAI22B_X1 T9882 ( .A1(T2005_Q), .B0(T9973_Y), .A0(T2028_Q),     .B1N(T10523_Y), .Y(T9882_Y));
KC_OAI22B_X1 T15848 ( .A1(T3845_Y), .B0(T5427_Y), .A0(T15699_Y),     .B1N(T14536_Q), .Y(T15848_Y));
KC_OAI22B_X1 T15901 ( .A1(T5106_Y), .B0(T3824_Y), .A0(T145_Q),     .B1N(T12181_Y), .Y(T15901_Y));
KC_OAI22B_X1 T15889 ( .A1(T3833_Y), .B0(T3834_Y), .A0(T11969_Y),     .B1N(T14544_Q), .Y(T15889_Y));
KC_OAI22B_X1 T15887 ( .A1(T5806_Y), .B0(T3832_Y), .A0(T5801_Y),     .B1N(T11393_Y), .Y(T15887_Y));
KC_NAND3BB_X1 T5897 ( .CN(T11512_Y), .Y(T5897_Y), .BN(T5459_Y),     .A(T5100_Y));
KC_AND4B_X1 T40 ( .D(T8561_Y), .C(T5630_Y), .B(T878_Y), .Y(T40_Y),     .AN(T5608_Y));
KC_AND4B_X1 T6849 ( .D(T2482_Y), .C(T2478_Y), .B(T2476_Y), .Y(T6849_Y),     .AN(T9745_Y));
KC_AND4B_X1 T5984 ( .D(T15968_Y), .C(T15945_Y), .B(T11505_Y),     .Y(T5984_Y), .AN(T11588_Y));
KC_AND3_X1 T16375 ( .C(T8767_Y), .B(T8829_Y), .A(T7645_Y),     .Y(T16375_Y));
KC_AND3_X1 T15843 ( .C(T2572_Q), .B(T2592_Q), .A(T2591_Q),     .Y(T15843_Y));
KC_AND3_X1 T15831 ( .C(T10251_Y), .B(T3218_Q), .A(T14522_Q),     .Y(T15831_Y));
KC_AND3_X1 T8385 ( .C(T6098_Y), .B(T15620_Y), .A(T4022_Y),     .Y(T8385_Y));
KC_DFFHQ_X2 T16445 ( .Q(T16445_Q), .CK(T991_Y), .D1(T8111_Y),     .D2(T15491_Y));
KC_DFFHQ_X2 T9048 ( .Q(T9048_Q), .CK(T1163_Y), .D1(T1150_Y),     .D2(T15521_Y));
KC_DFFHQ_X2 T16467 ( .Q(T16467_Q), .CK(T4282_Y), .D1(T12664_Y),     .D2(T15450_Y));
KC_TIEH_X1 T13068 ( .Y(T13068_Y));
KC_TIEH_X1 T13075 ( .Y(T13075_Y));
KC_TIEH_X1 T70 ( .Y(T70_Y));
KC_TIEH_X1 T15321 ( .Y(T15321_Y));
KC_TIEH_X1 T15407 ( .Y(T15407_Y));
KC_TIEH_X1 T15369 ( .Y(T15369_Y));
KC_TIEH_X1 T15484 ( .Y(T15484_Y));
KC_TIEH_X1 T15335 ( .Y(T15335_Y));
KC_TIEH_X1 T15673 ( .Y(T15673_Y));
KC_TIEH_X1 T15411 ( .Y(T15411_Y));
KC_TIEH_X1 T15496 ( .Y(T15496_Y));
KC_TIEH_X1 T15545 ( .Y(T15545_Y));
KC_TIEH_X1 T15342 ( .Y(T15342_Y));
KC_TIEH_X1 T15415 ( .Y(T15415_Y));
KC_TIEH_X1 T8671 ( .Y(T8671_Y));
KC_TIEH_X1 T984 ( .Y(T984_Y));
KC_TIEH_X1 T15480 ( .Y(T15480_Y));
KC_TIEH_X1 T15347 ( .Y(T15347_Y));
KC_TIEH_X1 T15381 ( .Y(T15381_Y));
KC_TIEH_X1 T6848 ( .Y(T6848_Y));
KC_TIEH_X1 T7837 ( .Y(T7837_Y));
KC_TIEH_X1 T16303 ( .Y(T16303_Y));
KC_TIEH_X1 T15551 ( .Y(T15551_Y));
KC_TIEH_X1 T15565 ( .Y(T15565_Y));
KC_TIEH_X1 T15639 ( .Y(T15639_Y));
KC_TIEH_X1 T3290 ( .Y(T3290_Y));
KC_TIEH_X1 T15594 ( .Y(T15594_Y));
KC_TIEH_X1 T4352 ( .Y(T4352_Y));
KC_TIEH_X1 T15366 ( .Y(T15366_Y));
KC_TIEH_X1 T6455 ( .Y(T6455_Y));
KC_TIEH_X1 T2724 ( .Y(T2724_Y));
KC_AOI22_X2 T8636 ( .Y(T8636_Y), .B1(T649_Q), .B0(T12415_Y),     .A1(T621_Q), .A0(T12417_Y));
KC_AOI22_X2 T8633 ( .Y(T8633_Y), .B1(T847_Q), .B0(T12414_Y),     .A1(T653_Q), .A0(T12416_Y));
KC_AOI22_X2 T8183 ( .Y(T8183_Y), .B1(T16488_Q), .B0(T12248_Y),     .A1(T15860_Q), .A0(T5848_Y));
KC_AOI22_X2 T8182 ( .Y(T8182_Y), .B1(T5432_Q), .B0(T5909_Y),     .A1(T2091_Q), .A0(T11499_Y));
KC_AOI22_X2 T8175 ( .Y(T8175_Y), .B1(T11410_Y), .B0(T5798_Y),     .A1(T11365_Y), .A0(T11408_Y));
KC_AOI22_X2 T8174 ( .Y(T8174_Y), .B1(T6742_Y), .B0(T15869_Y),     .A1(T11371_Y), .A0(T3826_Y));
KC_TLAT_X3 T106 ( .Q(T106_Q), .D(T134_Q), .G(T8804_Y));
KC_TLAT_X3 T141 ( .Q(T141_Q), .D(T16190_Y), .G(T9469_Q));
KC_TLAT_X3 T124 ( .Q(T124_Q), .D(T667_Y), .G(T8650_Y));
KC_TLAT_X3 T125 ( .Q(T125_Q), .D(T9853_Y), .G(T15054_Y));
KC_TLAT_X3 T145 ( .Q(T145_Q), .D(T15121_Y), .G(T4454_Q));
KC_TLAT_X3 T144 ( .Q(T144_Q), .D(T4456_Q), .G(T5044_Y));
KC_XOR2_X2 T16154 ( .Y(T16154_Y), .A(T16147_Y), .B(T5164_Q));
KC_MX2_X2 T16078 ( .Y(T16078_Y), .A(T1290_Y), .S0(T15544_Y),     .B(T15168_Q));
KC_MX2_X2 T8358 ( .Y(T8358_Y), .A(T15055_Y), .S0(T9855_Y),     .B(T5849_Y));
KC_MX2_X2 T16004 ( .Y(T16004_Y), .A(T10952_Y), .S0(T3294_Y),     .B(T15997_Y));
KC_MX2_X2 T16011 ( .Y(T16011_Y), .A(T8349_Y), .S0(T3294_Y),     .B(T15997_Y));
KC_MX2_X2 T16147 ( .Y(T16147_Y), .A(T3222_Y), .S0(T15909_Y),     .B(T12180_Y));
KC_MX2_X2 T15954 ( .Y(T15954_Y), .A(T5888_Y), .S0(T4533_Y),     .B(T8252_Y));
KC_AND4_X1 T15769 ( .D(T743_Y), .C(T647_Y), .B(T7581_Y), .A(T212_Q),     .Y(T15769_Y));
KC_AND4_X1 T15765 ( .D(T645_Y), .C(T647_Y), .B(T802_Y), .A(T223_Q),     .Y(T15765_Y));
KC_AND4_X1 T1096 ( .D(T954_Y), .C(T318_Y), .B(T321_Y), .A(T332_Y),     .Y(T1096_Y));
KC_AND4_X1 T6601 ( .D(T15388_Y), .C(T396_Y), .B(T386_Y), .A(T6608_Y),     .Y(T6601_Y));
KC_AND4_X1 T6808 ( .D(T164_Q), .C(T165_Q), .B(T664_Q), .A(T4837_Q),     .Y(T6808_Y));
KC_AND4_X1 T6249 ( .D(T15355_Y), .C(T6289_Y), .B(T15171_Y), .A(T345_Y),     .Y(T6249_Y));
KC_AND4_X1 T6248 ( .D(T6313_Y), .C(T304_Y), .B(T249_Y), .A(T6266_Y),     .Y(T6248_Y));
KC_AND4_X1 T6252 ( .D(T6257_Y), .C(T301_Y), .B(T245_Y), .A(T317_Y),     .Y(T6252_Y));
KC_AND4_X1 T6480 ( .D(T377_Y), .C(T379_Y), .B(T15390_Y), .A(T15391_Y),     .Y(T6480_Y));
KC_AND4_X1 T15817 ( .D(T10137_Y), .C(T5147_Y), .B(T10153_Y),     .A(T10136_Y), .Y(T15817_Y));
KC_AND4_X1 T15851 ( .D(T16474_Y), .C(T15881_Y), .B(T15882_Y),     .A(T2127_Y), .Y(T15851_Y));
KC_AND4_X1 T16016 ( .D(T2215_Y), .C(T2211_Y), .B(T2796_Y), .A(T2225_Y),     .Y(T16016_Y));
KC_AND4_X1 T6569 ( .D(T15633_Y), .C(T12103_Y), .B(T12107_Y),     .A(T12101_Y), .Y(T6569_Y));
KC_AND4_X1 T16051 ( .D(T6048_Y), .C(T12004_Y), .B(T15760_Q),     .A(T11641_Y), .Y(T16051_Y));
KC_AND4_X1 T6550 ( .D(T6517_Y), .C(T11813_Y), .B(T15637_Y),     .A(T11736_Y), .Y(T6550_Y));
KC_AND4_X1 T15782 ( .D(T4272_Y), .C(T5173_Y), .B(T4271_Y),     .A(T16444_Y), .Y(T15782_Y));
KC_AND4_X1 T15934 ( .D(T4483_Y), .C(T10629_Y), .B(T4497_Y),     .A(T4492_Q), .Y(T15934_Y));
KC_AND4_X1 T16013 ( .D(T6344_Y), .C(T4602_Q), .B(T5159_Q), .A(T4608_Q),     .Y(T16013_Y));
KC_NOR3B_X1 T5611 ( .Y(T5611_Y), .B(T5588_Y), .A(T48_Q), .CN(T5189_Q));
KC_NOR3B_X1 T58 ( .Y(T58_Y), .B(T5636_Y), .A(T5184_Q), .CN(T80_Y));
KC_NOR3B_X1 T6911 ( .Y(T6911_Y), .B(T6935_Y), .A(T8602_Y),     .CN(T8597_Y));
KC_NOR3B_X1 T8123 ( .Y(T8123_Y), .B(T8127_Y), .A(T8063_Y),     .CN(T8120_Y));
KC_NOR3B_X1 T15800 ( .Y(T15800_Y), .B(T745_Y), .A(T13241_Q),     .CN(T9028_Y));
KC_NOR3B_X1 T8037 ( .Y(T8037_Y), .B(T8117_Y), .A(T12368_Y),     .CN(T12456_Y));
KC_NOR3B_X1 T10660 ( .Y(T10660_Y), .B(T9983_Y), .A(T11914_Y),     .CN(T10163_Y));
KC_NOR3B_X1 T6216 ( .Y(T6216_Y), .B(T1773_Y), .A(T1769_Y),     .CN(T15923_Y));
KC_NOR3B_X1 T5906 ( .Y(T5906_Y), .B(T8394_Y), .A(T2001_Q),     .CN(T2054_Q));
KC_NOR3B_X1 T6235 ( .Y(T6235_Y), .B(T2755_Y), .A(T10928_Y),     .CN(T11449_Y));
KC_NOR3B_X1 T6579 ( .Y(T6579_Y), .B(T3514_Y), .A(T8417_Y),     .CN(T10547_Y));
KC_NOR3B_X1 T6722 ( .Y(T6722_Y), .B(T5433_Y), .A(T3202_Y),     .CN(T3204_Y));
KC_NOR3B_X1 T6035 ( .Y(T6035_Y), .B(T10243_Y), .A(T10241_Y),     .CN(T11959_Y));
KC_NOR3B_X1 T6352 ( .Y(T6352_Y), .B(T6022_Y), .A(T4606_Q),     .CN(T4590_Y));
KC_NOR3B_X1 T6219 ( .Y(T6219_Y), .B(T4535_Y), .A(T4489_Y),     .CN(T11453_Y));
KC_NOR3B_X1 T6344 ( .Y(T6344_Y), .B(T5158_Q), .A(T4606_Q),     .CN(T4607_Q));
KC_TINV_X1 T2521 ( .Y(T2521_Y), .A(T4641_Y), .OE(T4668_Y));
KC_OA21_X1 T8398 ( .B(T5145_Y), .A0(T6169_Y), .A1(T5152_Y),     .Y(T8398_Y));
KC_OAI21B_X2 T15047 ( .BN(T8851_Y), .A0(T659_Y), .A1(T9510_Y),     .Y(T15047_Y));
KC_OAI21B_X2 T15085 ( .BN(T10025_Y), .A0(T10006_Y), .A1(T10042_Y),     .Y(T15085_Y));
KC_OAI21B_X2 T15048 ( .BN(T1675_Q), .A0(T1665_Q), .A1(T7702_Y),     .Y(T15048_Y));
KC_OAI21B_X2 T15124 ( .BN(T11492_Y), .A0(T15916_Y), .A1(T15895_Y),     .Y(T15124_Y));
KC_OAI21B_X2 T15123 ( .BN(T11492_Y), .A0(T15916_Y), .A1(T15912_Y),     .Y(T15123_Y));
KC_OAI21B_X2 T15122 ( .BN(T11501_Y), .A0(T15916_Y), .A1(T2719_Y),     .Y(T15122_Y));
KC_OAI21B_X2 T15040 ( .BN(T11501_Y), .A0(T15916_Y), .A1(T15858_Y),     .Y(T15040_Y));
KC_OAI21B_X2 T15070 ( .BN(T15255_Y), .A0(T5027_Q), .A1(T15443_Y),     .Y(T15070_Y));
KC_OAI21B_X2 T15139 ( .BN(T5567_Q), .A0(T2854_Y), .A1(T4104_Y),     .Y(T15139_Y));
KC_OAI21B_X2 T15137 ( .BN(T12276_Y), .A0(T6077_Y), .A1(T11704_Y),     .Y(T15137_Y));
KC_OAI21B_X2 T15044 ( .BN(T2905_Y), .A0(T5517_Y), .A1(T10980_Y),     .Y(T15044_Y));
KC_OAI21B_X2 T15141 ( .BN(T11778_Y), .A0(T4704_Y), .A1(T10981_Y),     .Y(T15141_Y));
KC_INV_X3 T9 ( .Y(T9_Y), .A(T4003_Y));
KC_INV_X3 T8 ( .Y(T8_Y), .A(T4618_Y));
KC_INV_X3 T7 ( .Y(T7_Y), .A(T4004_Y));
KC_INV_X3 T2 ( .Y(T2_Y), .A(T4013_Y));
KC_INV_X3 T3 ( .Y(T3_Y), .A(T5482_Y));
KC_INV_X3 T4 ( .Y(T4_Y), .A(T1824_Y));
KC_INV_X3 T5 ( .Y(T5_Y), .A(T3994_Y));
KC_INV_X3 T6 ( .Y(T6_Y), .A(T4002_Y));
KC_INV_X3 T10 ( .Y(T10_Y), .A(T4619_Y));
KC_INV_X3 T11 ( .Y(T11_Y), .A(T4012_Y));
KC_INV_X3 T12 ( .Y(T12_Y), .A(T3995_Y));
KC_INV_X3 T13 ( .Y(T13_Y), .A(T4005_Y));
KC_INV_X3 T14 ( .Y(T14_Y), .A(T4000_Y));
KC_INV_X3 T15 ( .Y(T15_Y), .A(T4620_Y));
KC_INV_X3 T16 ( .Y(T16_Y), .A(T4001_Y));
KC_INV_X3 T17 ( .Y(T17_Y), .A(T4610_Y));
KC_INV_X3 T1748 ( .Y(T1748_Y), .A(T15805_Q));
KC_INV_X3 T2751 ( .Y(T2751_Y), .A(T15807_Q));
KC_INV_X3 T16238 ( .Y(T16238_Y), .A(T13_Y));
KC_INV_X3 T16200 ( .Y(T16200_Y), .A(T4_Y));
KC_INV_X3 T16199 ( .Y(T16199_Y), .A(T15_Y));
KC_INV_X3 T16198 ( .Y(T16198_Y), .A(T12_Y));
KC_INV_X3 T16197 ( .Y(T16197_Y), .A(T14_Y));
KC_INV_X3 T16196 ( .Y(T16196_Y), .A(T16_Y));
KC_INV_X3 T16174 ( .Y(T16174_Y), .A(T3_Y));
KC_INV_X3 T16155 ( .Y(T16155_Y), .A(T7_Y));
KC_INV_X3 T4796 ( .Y(T4796_Y), .A(T6_Y));
KC_INV_X3 T4428 ( .Y(T4428_Y), .A(T10_Y));
KC_INV_X3 T4408 ( .Y(T4408_Y), .A(T9_Y));
KC_INV_X3 T4407 ( .Y(T4407_Y), .A(T11_Y));
KC_INV_X3 T4413 ( .Y(T4413_Y), .A(T17_Y));
KC_INV_X3 T4414 ( .Y(T4414_Y), .A(T2_Y));
KC_INV_X3 T4423 ( .Y(T4423_Y), .A(T8_Y));
KC_INV_X3 T4422 ( .Y(T4422_Y), .A(T5_Y));
KC_INV_X3 T4795 ( .Y(T4795_Y), .A(T4422_Y));
KC_INV_X3 T4792 ( .Y(T4792_Y), .A(T4414_Y));
KC_INV_X3 T4791 ( .Y(T4791_Y), .A(T16200_Y));
KC_INV_X3 T298 ( .Y(T298_Y), .A(T16198_Y));
KC_INV_X3 T15949 ( .Y(T15949_Y), .A(T4796_Y));
KC_INV_X3 T15687 ( .Y(T15687_Y), .A(T16174_Y));
KC_INV_X3 T4794 ( .Y(T4794_Y), .A(T4413_Y));
KC_INV_X3 T4793 ( .Y(T4793_Y), .A(T16199_Y));
KC_INV_X3 T4790 ( .Y(T4790_Y), .A(T16155_Y));
KC_INV_X3 T4789 ( .Y(T4789_Y), .A(T4428_Y));
KC_INV_X3 T4785 ( .Y(T4785_Y), .A(T4407_Y));
KC_INV_X3 T4786 ( .Y(T4786_Y), .A(T16197_Y));
KC_INV_X3 T4779 ( .Y(T4779_Y), .A(T4423_Y));
KC_INV_X3 T4781 ( .Y(T4781_Y), .A(T4408_Y));
KC_INV_X3 T4778 ( .Y(T4778_Y), .A(T16196_Y));
KC_INV_X3 T4780 ( .Y(T4780_Y), .A(T16238_Y));
KC_BUF_X16 T4409 ( .Y(T4409_Y), .A(T13263_Q));
KC_DFFRNHQ_X5 T16410 ( .Q(T16410_Q), .D(T15469_Y), .RN(T16182_Y),     .CK(T1055_Y));
KC_DFFRNHQ_X5 T16409 ( .Q(T16409_Q), .D(T15467_Y), .RN(T16182_Y),     .CK(T15167_Y));
KC_DFFRNHQ_X5 T16468 ( .Q(T16468_Q), .D(T16436_Y), .RN(T16182_Y),     .CK(T15469_Y));
KC_DFFRNHQ_X5 T16464 ( .Q(T16464_Q), .D(T1055_Y), .RN(T16182_Y),     .CK(T15467_Y));
KC_DFFRNHQ_X5 T16470 ( .Q(T16470_Q), .D(T1690_Q), .RN(T14988_Y),     .CK(T1598_Y));
KC_DFFHQ_X3 T16446 ( .Q(T16446_Q), .CK(T13057_Q), .D(T15006_Y));
KC_AND2_X4 T225 ( .B(T15333_Y), .A(T662_Y), .Y(T225_Y));
KC_AND2_X4 T118 ( .B(T15333_Y), .A(T662_Y), .Y(T118_Y));
KC_AND2_X4 T16407 ( .B(T16434_Q), .A(T4922_Y), .Y(T16407_Y));
KC_AO112BB_X1 T6750 ( .D(T10261_Y), .Y(T6750_Y), .C(T10918_Y),     .A(T2474_Y), .B(T4887_Y));
KC_AO112BB_X1 T16254 ( .D(T16244_Y), .Y(T16254_Y), .C(T10906_Y),     .A(T2566_Y), .B(T16261_Y));
KC_MXI2_X3 T13264 ( .Y(T13264_Y), .A(T4813_Y), .B(T4814_Y),     .S0(T9166_Y));
KC_MXI2_X3 T13260 ( .Y(T13260_Y), .A(T997_Q), .B(T9457_Q),     .S0(T15795_Q));
KC_MXI2_X3 T13060 ( .Y(T13060_Y), .A(T15855_Y), .B(T15796_Q),     .S0(T1025_Y));
KC_MXI2_X3 T13082 ( .Y(T13082_Y), .A(T2835_Q), .B(T11447_Y),     .S0(T15014_Y));
KC_MXI2_X3 T13113 ( .Y(T13113_Y), .A(T2281_Q), .B(T11467_Y),     .S0(T3294_Y));
KC_MXI2_X3 T13105 ( .Y(T13105_Y), .A(T5380_Q), .B(T15912_Y),     .S0(T3256_Q));
KC_MXI2_X3 T13097 ( .Y(T13097_Y), .A(T2249_Q), .B(T11469_Y),     .S0(T3294_Y));
KC_MXI2_X3 T13131 ( .Y(T13131_Y), .A(T5525_Q), .B(T3927_Y),     .S0(T3294_Y));
KC_MXI2_X3 T13121 ( .Y(T13121_Y), .A(T4147_Q), .B(T16500_Y),     .S0(T3294_Y));
KC_MXI2_X3 T12982 ( .Y(T12982_Y), .A(T4176_Q), .B(T3928_Y),     .S0(T3294_Y));
KC_MXI2_X3 T13125 ( .Y(T13125_Y), .A(T4179_Q), .B(T5459_Y),     .S0(T3294_Y));
KC_MXI2_X3 T13300 ( .Y(T13300_Y), .A(T2275_Q), .B(T3869_Y),     .S0(T15014_Y));
KC_XNOR2_X6 T16456 ( .Y(T16456_Y), .A(T12838_Y), .B(T11479_Y));
KC_AOI222_X1 T12808 ( .A0(T11499_Y), .Y(T12808_Y), .C1(T2382_Q),     .C0(T5944_Y), .B1(T2161_Q), .B0(T5909_Y), .A1(T2125_Y));
KC_AOI222_X1 T12871 ( .A0(T8422_Y), .Y(T12871_Y), .C1(T15138_Q),     .C0(T10995_Y), .B1(T12105_Y), .B0(T10553_Y), .A1(T6238_Y));
KC_AOI222_X1 T12567 ( .A0(T3020_Y), .Y(T12567_Y), .C1(T2991_Y),     .C0(T9669_Y), .B1(T2448_Y), .B0(T3020_Y), .A1(T478_Y));
KC_AOI222_X1 T12559 ( .A0(T5080_Y), .Y(T12559_Y), .C1(T2962_Y),     .C0(T9655_Y), .B1(T2448_Y), .B0(T5080_Y), .A1(T431_Y));
KC_AOI222_X1 T12556 ( .A0(T5080_Y), .Y(T12556_Y), .C1(T3549_Y),     .C0(T9655_Y), .B1(T2448_Y), .B0(T5080_Y), .A1(T423_Y));
KC_AOI222_X1 T12466 ( .A0(T4101_Y), .Y(T12466_Y), .C1(T10584_Y),     .C0(T3435_Y), .B1(T10585_Y), .B0(T4079_Y), .A1(T11746_Y));
KC_AOI222_X1 T12864 ( .A0(T3469_Y), .Y(T12864_Y), .C1(T15631_Y),     .C0(T8408_Y), .B1(T6503_S), .B0(T6210_Y), .A1(T5530_Q));
KC_AOI222_X1 T12860 ( .A0(T3469_Y), .Y(T12860_Y), .C1(T4540_Y),     .C0(T6574_Y), .B1(T15631_Y), .B0(T2927_Y), .A1(T4176_Q));
KC_AOI222_X1 T12467 ( .A0(T3469_Y), .Y(T12467_Y), .C1(T6842_S),     .C0(T6210_Y), .B1(T6193_Y), .B0(T3480_Y), .A1(T15760_Q));
KC_AOI222_X1 T12800 ( .A0(T3850_Y), .Y(T12800_Y), .C1(T11410_Y),     .C0(T5553_Y), .B1(T5830_Y), .B0(T14551_Q), .A1(T15907_Y));
KC_AOI222_X1 T12798 ( .A0(T11398_Y), .Y(T12798_Y), .C1(T11371_Y),     .C0(T4439_Y), .B1(T4487_Q), .B0(T11399_Y), .A1(T4457_Y));
KC_AOI222_X1 T12972 ( .A0(T12465_Y), .Y(T12972_Y), .C1(T6214_Y),     .C0(T15233_Y), .B1(T10551_Y), .B0(T10555_Y), .A1(T12317_Y));
KC_AOI222_X1 T12943 ( .A0(T2629_Y), .Y(T12943_Y), .C1(T5321_Y),     .C0(T1508_Y), .B1(T16363_Y), .B0(T2629_Y), .A1(T1508_Y));
KC_AOI222_X1 T12964 ( .A0(T16108_Y), .Y(T12964_Y), .C1(T12290_Y),     .C0(T4059_Y), .B1(T4016_Y), .B0(T16108_Y), .A1(T16107_Y));
KC_NAND3B_X1 T5622 ( .CN(T15213_Y), .Y(T5622_Y), .B(T16176_Y),     .A(T878_Y));
KC_NAND3B_X1 T9286 ( .CN(T9288_Y), .Y(T9286_Y), .B(T260_Y),     .A(T133_Q));
KC_NAND3B_X1 T9269 ( .CN(T6321_Y), .Y(T9269_Y), .B(T133_Q),     .A(T8579_Y));
KC_NAND3B_X1 T9025 ( .CN(T1448_Y), .Y(T9025_Y), .B(T9455_Y),     .A(T15492_Y));
KC_NAND3B_X1 T8994 ( .CN(T8992_Y), .Y(T8994_Y), .B(T15099_Y),     .A(T1386_Y));
KC_NAND3B_X1 T7913 ( .CN(T7917_Y), .Y(T7913_Y), .B(T8080_Y),     .A(T7916_Y));
KC_NAND3B_X1 T7892 ( .CN(T16388_Y), .Y(T7892_Y), .B(T758_Y),     .A(T8946_Y));
KC_NAND3B_X1 T7866 ( .CN(T16159_Y), .Y(T7866_Y), .B(T10941_Y),     .A(T988_Y));
KC_NAND3B_X1 T7835 ( .CN(T7834_Y), .Y(T7835_Y), .B(T952_Y),     .A(T7844_Y));
KC_NAND3B_X1 T7834 ( .CN(T8790_Y), .Y(T7834_Y), .B(T8849_Y),     .A(T9402_Y));
KC_NAND3B_X1 T6889 ( .CN(T6893_Y), .Y(T6889_Y), .B(T1521_Y),     .A(T1521_Y));
KC_NAND3B_X1 T10318 ( .CN(T9782_Y), .Y(T10318_Y), .B(T9782_Y),     .A(T1563_Y));
KC_NAND3B_X1 T1834 ( .CN(T11046_Y), .Y(T1834_Y), .B(T1847_Y),     .A(T11845_Y));
KC_NAND3B_X1 T2107 ( .CN(T3339_Y), .Y(T2107_Y), .B(T2148_Y),     .A(T12794_Y));
KC_NAND3B_X1 T2166 ( .CN(T10928_Y), .Y(T2166_Y), .B(T11436_Y),     .A(T11597_Y));
KC_NAND3B_X1 T2321 ( .CN(T15713_Y), .Y(T2321_Y), .B(T2348_Y),     .A(T10562_Y));
KC_NAND3B_X1 T2371 ( .CN(T2369_Y), .Y(T2371_Y), .B(T12072_Y),     .A(T2369_Y));
KC_NAND3B_X1 T2374 ( .CN(T2369_Y), .Y(T2374_Y), .B(T2369_Y),     .A(T6500_Y));
KC_NAND3B_X1 T2504 ( .CN(T16195_Y), .Y(T2504_Y), .B(T882_Y),     .A(T16447_Y));
KC_NAND3B_X1 T2505 ( .CN(T16447_Y), .Y(T2505_Y), .B(T882_Y),     .A(T16195_Y));
KC_NAND3B_X1 T2551 ( .CN(T2545_Y), .Y(T2551_Y), .B(T16363_Y),     .A(T2571_Q));
KC_NAND3B_X1 T2593 ( .CN(T16245_Y), .Y(T2593_Y), .B(T1544_Y),     .A(T3741_Y));
KC_NAND3B_X1 T2604 ( .CN(T10104_Y), .Y(T2604_Y), .B(T15518_Y),     .A(T10101_Y));
KC_NAND3B_X1 T2665 ( .CN(T10244_Y), .Y(T2665_Y), .B(T12128_Y),     .A(T15442_Y));
KC_NAND3B_X1 T2705 ( .CN(T8198_Y), .Y(T2705_Y), .B(T15886_Y),     .A(T2703_Y));
KC_NAND3B_X1 T2723 ( .CN(T2721_Y), .Y(T2723_Y), .B(T2740_Y),     .A(T2739_Y));
KC_NAND3B_X1 T2852 ( .CN(T3404_Y), .Y(T2852_Y), .B(T12267_Y),     .A(T12046_Y));
KC_NAND3B_X1 T2862 ( .CN(T6556_Y), .Y(T2862_Y), .B(T3424_Y),     .A(T6237_Y));
KC_NAND3B_X1 T2914 ( .CN(T2891_Y), .Y(T2914_Y), .B(T6576_Y),     .A(T2330_Y));
KC_NAND3B_X1 T3208 ( .CN(T3201_Y), .Y(T3208_Y), .B(T3213_Q),     .A(T5428_Q));
KC_NAND3B_X1 T3285 ( .CN(T6230_Co), .Y(T3285_Y), .B(T3309_Y),     .A(T12210_Y));
KC_NAND3B_X1 T3287 ( .CN(T3286_Y), .Y(T3287_Y), .B(T3298_Y),     .A(T3289_Y));
KC_NAND3B_X1 T3391 ( .CN(T11662_Y), .Y(T3391_Y), .B(T3384_Y),     .A(T3369_Y));
KC_NAND3B_X1 T3403 ( .CN(T3401_Y), .Y(T3403_Y), .B(T12002_Y),     .A(T6123_Y));
KC_NAND3B_X1 T3421 ( .CN(T11725_Y), .Y(T3421_Y), .B(T3436_Y),     .A(T11676_Y));
KC_NAND3B_X1 T3915 ( .CN(T5936_Y), .Y(T3915_Y), .B(T10202_Y),     .A(T15130_Y));
KC_NAND3B_X1 T4158 ( .CN(T8163_Y), .Y(T4158_Y), .B(T4761_Y),     .A(T3996_Y));
KC_NAND3B_X1 T4467 ( .CN(T4488_Y), .Y(T4467_Y), .B(T5142_Y),     .A(T4470_Y));
KC_NAND3B_X1 T4547 ( .CN(T4572_Q), .Y(T4547_Y), .B(T15584_Y),     .A(T12016_Y));
KC_NAND3B_X1 T4705 ( .CN(T13165_Q), .Y(T4705_Y), .B(T5464_Y),     .A(T5512_Q));
KC_NAND3B_X1 T4737 ( .CN(T4749_Y), .Y(T4737_Y), .B(T6187_Y),     .A(T4747_Y));
KC_NAND3B_X1 T5057 ( .CN(T12215_Y), .Y(T5057_Y), .B(T15162_Y),     .A(T3344_Y));
KC_NAND3B_X1 T5114 ( .CN(T3984_Y), .Y(T5114_Y), .B(T4928_Y),     .A(T4928_Y));
KC_NAND2_X1 T27 ( .B(T13068_Y), .A(T29_Y), .Y(T27_Y));
KC_NAND2_X1 T5592 ( .B(T13075_Y), .A(T35_Y), .Y(T5592_Y));
KC_NAND2_X1 T5581 ( .B(T13075_Y), .A(T5593_Y), .Y(T5581_Y));
KC_NAND2_X1 T68 ( .B(T70_Y), .A(T82_Y), .Y(T68_Y));
KC_NAND2_X1 T73 ( .B(T70_Y), .A(T56_Y), .Y(T73_Y));
KC_NAND2_X1 T92 ( .B(T15321_Y), .A(T90_Y), .Y(T92_Y));
KC_NAND2_X1 T93 ( .B(T15321_Y), .A(T97_Y), .Y(T93_Y));
KC_NAND2_X1 T201 ( .B(T15407_Y), .A(GND), .Y(T201_Y));
KC_NAND2_X1 T468 ( .B(T15369_Y), .A(T465_Y), .Y(T468_Y));
KC_NAND2_X1 T480 ( .B(T15369_Y), .A(T466_Y), .Y(T480_Y));
KC_NAND2_X1 T576 ( .B(T15484_Y), .A(T575_Y), .Y(T576_Y));
KC_NAND2_X1 T584 ( .B(T15484_Y), .A(T582_Y), .Y(T584_Y));
KC_NAND2_X1 T16310 ( .B(T747_Q), .A(T977_Q), .Y(T16310_Y));
KC_NAND2_X1 T800 ( .B(T15335_Y), .A(T798_Y), .Y(T800_Y));
KC_NAND2_X1 T801 ( .B(T15335_Y), .A(T792_Y), .Y(T801_Y));
KC_NAND2_X1 T6835 ( .B(T7599_Y), .A(T9360_Y), .Y(T6835_Y));
KC_NAND2_X1 T6803 ( .B(T7599_Y), .A(T9359_Y), .Y(T6803_Y));
KC_NAND2_X1 T894 ( .B(T15411_Y), .A(T891_Y), .Y(T894_Y));
KC_NAND2_X1 T895 ( .B(T15411_Y), .A(T890_Y), .Y(T895_Y));
KC_NAND2_X1 T896 ( .B(T7599_Y), .A(T553_Y), .Y(T896_Y));
KC_NAND2_X1 T1028 ( .B(T15673_Y), .A(T5557_Y), .Y(T1028_Y));
KC_NAND2_X1 T1032 ( .B(T15673_Y), .A(T1030_Y), .Y(T1032_Y));
KC_NAND2_X1 T1230 ( .B(T15496_Y), .A(T1229_Y), .Y(T1230_Y));
KC_NAND2_X1 T1242 ( .B(T15496_Y), .A(T1240_Y), .Y(T1242_Y));
KC_NAND2_X1 T1320 ( .B(T15342_Y), .A(T1318_Y), .Y(T1320_Y));
KC_NAND2_X1 T1398 ( .B(T15342_Y), .A(T1390_Y), .Y(T1398_Y));
KC_NAND2_X1 T1467 ( .B(T15415_Y), .A(T1464_Y), .Y(T1467_Y));
KC_NAND2_X1 T1468 ( .B(T15415_Y), .A(T1463_Y), .Y(T1468_Y));
KC_NAND2_X1 T1536 ( .B(T8671_Y), .A(T1534_Y), .Y(T1536_Y));
KC_NAND2_X1 T1541 ( .B(T8671_Y), .A(T1540_Y), .Y(T1541_Y));
KC_NAND2_X1 T1572 ( .B(T984_Y), .A(T1569_Y), .Y(T1572_Y));
KC_NAND2_X1 T1591 ( .B(T984_Y), .A(T1589_Y), .Y(T1591_Y));
KC_NAND2_X1 T1863 ( .B(T15347_Y), .A(T1862_Y), .Y(T1863_Y));
KC_NAND2_X1 T1870 ( .B(T15347_Y), .A(T1866_Y), .Y(T1870_Y));
KC_NAND2_X1 T1966 ( .B(T6848_Y), .A(T1965_Y), .Y(T1966_Y));
KC_NAND2_X1 T2442 ( .B(T15381_Y), .A(T2441_Y), .Y(T2442_Y));
KC_NAND2_X1 T2445 ( .B(T15381_Y), .A(T2443_Y), .Y(T2445_Y));
KC_NAND2_X1 T6481 ( .B(T2449_Y), .A(T14984_Y), .Y(T6481_Y));
KC_NAND2_X1 T10261 ( .B(T9780_Y), .A(T10493_Y), .Y(T10261_Y));
KC_NAND2_X1 T10254 ( .B(T9780_Y), .A(T9747_Y), .Y(T10254_Y));
KC_NAND2_X1 T2490 ( .B(T6848_Y), .A(T2488_Y), .Y(T2490_Y));
KC_NAND2_X1 T2492 ( .B(T9874_Y), .A(T9854_Y), .Y(T2492_Y));
KC_NAND2_X1 T16245 ( .B(T10239_Y), .A(T2564_Y), .Y(T16245_Y));
KC_NAND2_X1 T3155 ( .B(T16303_Y), .A(GND), .Y(T3155_Y));
KC_NAND2_X1 T3160 ( .B(T16303_Y), .A(T3158_Y), .Y(T3160_Y));
KC_NAND2_X1 T3189 ( .B(T15551_Y), .A(T3188_Y), .Y(T3189_Y));
KC_NAND2_X1 T3194 ( .B(T15551_Y), .A(T3191_Y), .Y(T3194_Y));
KC_NAND2_X1 T3236 ( .B(T15565_Y), .A(T3239_Y), .Y(T3236_Y));
KC_NAND2_X1 T3237 ( .B(T15565_Y), .A(T3234_Y), .Y(T3237_Y));
KC_NAND2_X1 T3504 ( .B(T15639_Y), .A(T5531_Y), .Y(T3504_Y));
KC_NAND2_X1 T3505 ( .B(T15639_Y), .A(T5542_Y), .Y(T3505_Y));
KC_NAND2_X1 T3641 ( .B(T3290_Y), .A(T3638_Y), .Y(T3641_Y));
KC_NAND2_X1 T3644 ( .B(T3290_Y), .A(T3643_Y), .Y(T3644_Y));
KC_NAND2_X1 T15835 ( .B(T11985_Y), .A(T11389_Y), .Y(T15835_Y));
KC_NAND2_X1 T15825 ( .B(T11322_Y), .A(T5763_Y), .Y(T15825_Y));
KC_NAND2_X1 T3929 ( .B(T15594_Y), .A(T3938_Y), .Y(T3929_Y));
KC_NAND2_X1 T3958 ( .B(T15594_Y), .A(T3957_Y), .Y(T3958_Y));
KC_NAND2_X1 T4041 ( .B(T4352_Y), .A(T4039_Y), .Y(T4041_Y));
KC_NAND2_X1 T4199 ( .B(T15366_Y), .A(T4190_Y), .Y(T4199_Y));
KC_NAND2_X1 T4200 ( .B(T15366_Y), .A(T4198_Y), .Y(T4200_Y));
KC_NAND2_X1 T4208 ( .B(T6455_Y), .A(T5175_Y), .Y(T4208_Y));
KC_NAND2_X1 T4229 ( .B(T6455_Y), .A(T4227_Y), .Y(T4229_Y));
KC_NAND2_X1 T4334 ( .B(T2724_Y), .A(T4332_Y), .Y(T4334_Y));
KC_NAND2_X1 T4335 ( .B(T2724_Y), .A(T4331_Y), .Y(T4335_Y));
KC_NAND2_X1 T4797 ( .B(T13068_Y), .A(T4798_Y), .Y(T4797_Y));
KC_NAND2_X1 T15740 ( .B(T7599_Y), .A(T9362_Y), .Y(T15740_Y));
KC_NAND2_X1 T8238 ( .B(T15943_Y), .A(T2848_Y), .Y(T8238_Y));
KC_NAND2_X1 T16005 ( .B(T16004_Y), .A(T16011_Y), .Y(T16005_Y));
KC_NAND2_X1 T16451 ( .B(T14947_Q), .A(T2566_Y), .Y(T16451_Y));
KC_NAND2_X1 T16450 ( .B(T14510_Q), .A(T2566_Y), .Y(T16450_Y));
KC_NAND2_X1 T5128 ( .B(T4352_Y), .A(T5127_Y), .Y(T5128_Y));
KC_XOR2_X1 T16063 ( .Y(T16063_Y), .A(T15537_Y), .B(T5548_Y));
KC_XOR2_X1 T13055 ( .Y(T13055_Y), .A(T9227_Y), .B(T11562_Y));
KC_XOR2_X1 T16083 ( .Y(T16083_Y), .A(T12282_Y), .B(T3336_Y));
KC_XOR2_X1 T6443 ( .Y(T6443_Y), .A(T4189_Y), .B(T9590_Y));
KC_XOR2_X1 T16153 ( .Y(T16153_Y), .A(T15156_Y), .B(T4455_Q));
KC_XOR2_X1 T16152 ( .Y(T16152_Y), .A(T3315_Y), .B(T15043_Y));
KC_XOR2_X1 T15908 ( .Y(T15908_Y), .A(T12151_Y), .B(T5165_Q));
KC_INV_X2 T22 ( .Y(T22_Y), .A(T4797_Y));
KC_INV_X2 T31 ( .Y(T31_Y), .A(T27_Y));
KC_INV_X2 T42 ( .Y(T42_Y), .A(T5581_Y));
KC_INV_X2 T43 ( .Y(T43_Y), .A(T5592_Y));
KC_INV_X2 T67 ( .Y(T67_Y), .A(T68_Y));
KC_INV_X2 T78 ( .Y(T78_Y), .A(T73_Y));
KC_INV_X2 T91 ( .Y(T91_Y), .A(T93_Y));
KC_INV_X2 T99 ( .Y(T99_Y), .A(T92_Y));
KC_INV_X2 T199 ( .Y(T199_Y), .A(T197_Y));
KC_INV_X2 T200 ( .Y(T200_Y), .A(T201_Y));
KC_INV_X2 T467 ( .Y(T467_Y), .A(T468_Y));
KC_INV_X2 T479 ( .Y(T479_Y), .A(T480_Y));
KC_INV_X2 T533 ( .Y(T533_Y), .A(T576_Y));
KC_INV_X2 T583 ( .Y(T583_Y), .A(T584_Y));
KC_INV_X2 T15720 ( .Y(T15720_Y), .A(T801_Y));
KC_INV_X2 T799 ( .Y(T799_Y), .A(T800_Y));
KC_INV_X2 T892 ( .Y(T892_Y), .A(T895_Y));
KC_INV_X2 T893 ( .Y(T893_Y), .A(T894_Y));
KC_INV_X2 T1031 ( .Y(T1031_Y), .A(T1032_Y));
KC_INV_X2 T1194 ( .Y(T1194_Y), .A(T1242_Y));
KC_INV_X2 T1241 ( .Y(T1241_Y), .A(T1230_Y));
KC_INV_X2 T1285 ( .Y(T1285_Y), .A(T192_Y));
KC_INV_X2 T1290 ( .Y(T1290_Y), .A(T16392_Y));
KC_INV_X2 T1319 ( .Y(T1319_Y), .A(T1320_Y));
KC_INV_X2 T1362 ( .Y(T1362_Y), .A(T10936_Y));
KC_INV_X2 T1365 ( .Y(T1365_Y), .A(T13125_Y));
KC_INV_X2 T1366 ( .Y(T1366_Y), .A(T10934_Y));
KC_INV_X2 T1383 ( .Y(T1383_Y), .A(T15188_Y));
KC_INV_X2 T1397 ( .Y(T1397_Y), .A(T1398_Y));
KC_INV_X2 T1465 ( .Y(T1465_Y), .A(T1468_Y));
KC_INV_X2 T1466 ( .Y(T1466_Y), .A(T1467_Y));
KC_INV_X2 T1528 ( .Y(T1528_Y), .A(T1536_Y));
KC_INV_X2 T1530 ( .Y(T1530_Y), .A(T1541_Y));
KC_INV_X2 T1570 ( .Y(T1570_Y), .A(T1572_Y));
KC_INV_X2 T1578 ( .Y(T1578_Y), .A(T13113_Y));
KC_INV_X2 T1590 ( .Y(T1590_Y), .A(T1591_Y));
KC_INV_X2 T1597 ( .Y(T1597_Y), .A(T13097_Y));
KC_INV_X2 T1633 ( .Y(T1633_Y), .A(T3072_Y));
KC_INV_X2 T1709 ( .Y(T1709_Y), .A(T13300_Y));
KC_INV_X2 T1724 ( .Y(T1724_Y), .A(T10912_Y));
KC_INV_X2 T1786 ( .Y(T1786_Y), .A(T2315_Q));
KC_INV_X2 T1788 ( .Y(T1788_Y), .A(T2311_Q));
KC_INV_X2 T1804 ( .Y(T1804_Y), .A(T1820_Q));
KC_INV_X2 T1805 ( .Y(T1805_Y), .A(T1822_Q));
KC_INV_X2 T1864 ( .Y(T1864_Y), .A(T1863_Y));
KC_INV_X2 T1867 ( .Y(T1867_Y), .A(T1870_Y));
KC_INV_X2 T16240 ( .Y(T16240_Y), .A(T2490_Y));
KC_INV_X2 T1962 ( .Y(T1962_Y), .A(T1966_Y));
KC_INV_X2 T2127 ( .Y(T2127_Y), .A(T15798_Q));
KC_INV_X2 T2239 ( .Y(T2239_Y), .A(T2237_Q));
KC_INV_X2 T2240 ( .Y(T2240_Y), .A(T4964_Q));
KC_INV_X2 T2245 ( .Y(T2245_Y), .A(T5494_Q));
KC_INV_X2 T2246 ( .Y(T2246_Y), .A(T5486_Q));
KC_INV_X2 T2247 ( .Y(T2247_Y), .A(T2314_Q));
KC_INV_X2 T2250 ( .Y(T2250_Y), .A(T2313_Q));
KC_INV_X2 T2279 ( .Y(T2279_Y), .A(T6419_Q));
KC_INV_X2 T2280 ( .Y(T2280_Y), .A(T5497_Q));
KC_INV_X2 T2344 ( .Y(T2344_Y), .A(T5566_Q));
KC_INV_X2 T2438 ( .Y(T2438_Y), .A(T2442_Y));
KC_INV_X2 T2444 ( .Y(T2444_Y), .A(T2445_Y));
KC_INV_X2 T2448 ( .Y(T2448_Y), .A(T14984_Y));
KC_INV_X2 T2451 ( .Y(T2451_Y), .A(T3640_Y));
KC_INV_X2 T2620 ( .Y(T2620_Y), .A(T14994_Y));
KC_INV_X2 T2708 ( .Y(T2708_Y), .A(T15894_Q));
KC_INV_X2 T2717 ( .Y(T2717_Y), .A(T8482_Y));
KC_INV_X2 T2719 ( .Y(T2719_Y), .A(T16301_Q));
KC_INV_X2 T2839 ( .Y(T2839_Y), .A(T2879_Y));
KC_INV_X2 T2848 ( .Y(T2848_Y), .A(T6515_Y));
KC_INV_X2 T3154 ( .Y(T3154_Y), .A(T3155_Y));
KC_INV_X2 T3159 ( .Y(T3159_Y), .A(T3160_Y));
KC_INV_X2 T3192 ( .Y(T3192_Y), .A(T3194_Y));
KC_INV_X2 T3193 ( .Y(T3193_Y), .A(T3189_Y));
KC_INV_X2 T16239 ( .Y(T16239_Y), .A(T3236_Y));
KC_INV_X2 T3235 ( .Y(T3235_Y), .A(T3237_Y));
KC_INV_X2 T3317 ( .Y(T3317_Y), .A(T3929_Y));
KC_INV_X2 T3331 ( .Y(T3331_Y), .A(T10949_Y));
KC_INV_X2 T3501 ( .Y(T3501_Y), .A(T3504_Y));
KC_INV_X2 T3534 ( .Y(T3534_Y), .A(T3505_Y));
KC_INV_X2 T3639 ( .Y(T3639_Y), .A(T3641_Y));
KC_INV_X2 T3648 ( .Y(T3648_Y), .A(T3644_Y));
KC_INV_X2 T3683 ( .Y(T3683_Y), .A(T3684_Y));
KC_INV_X2 T3856 ( .Y(T3856_Y), .A(T16154_Y));
KC_INV_X2 T3872 ( .Y(T3872_Y), .A(T10943_Y));
KC_INV_X2 T16242 ( .Y(T16242_Y), .A(T5128_Y));
KC_INV_X2 T4040 ( .Y(T4040_Y), .A(T4041_Y));
KC_INV_X2 T4184 ( .Y(T4184_Y), .A(T4200_Y));
KC_INV_X2 T4192 ( .Y(T4192_Y), .A(T4199_Y));
KC_INV_X2 T4228 ( .Y(T4228_Y), .A(T4229_Y));
KC_INV_X2 T5913 ( .Y(T5913_Y), .A(T4334_Y));
KC_INV_X2 T4333 ( .Y(T4333_Y), .A(T4335_Y));
KC_INV_X2 T4486 ( .Y(T4486_Y), .A(T4463_Y));
KC_INV_X2 T4856 ( .Y(T4856_Y), .A(T1028_Y));
KC_INV_X2 T4872 ( .Y(T4872_Y), .A(T10941_Y));
KC_INV_X2 T4901 ( .Y(T4901_Y), .A(T16079_Q));
KC_INV_X2 T4922 ( .Y(T4922_Y), .A(T16470_Q));
KC_INV_X2 T4926 ( .Y(T4926_Y), .A(T5524_Q));
KC_INV_X2 T4968 ( .Y(T4968_Y), .A(T16082_Q));
KC_INV_X2 T5026 ( .Y(T5026_Y), .A(T16079_Q));
KC_INV_X2 T5070 ( .Y(T5070_Y), .A(T6526_Q));
KC_INV_X2 T5072 ( .Y(T5072_Y), .A(T6549_Q));
KC_INV_X2 T5121 ( .Y(T5121_Y), .A(T3958_Y));
KC_INV_X2 T5176 ( .Y(T5176_Y), .A(T4208_Y));
KC_INV_X4 T24 ( .Y(T24_Y), .A(T26_Y));
KC_INV_X4 T30 ( .Y(T30_Y), .A(T5230_Y));
KC_INV_X4 T37 ( .Y(T37_Y), .A(T39_Y));
KC_INV_X4 T49 ( .Y(T49_Y), .A(T5584_Y));
KC_INV_X4 T63 ( .Y(T63_Y), .A(T65_Y));
KC_INV_X4 T74 ( .Y(T74_Y), .A(T75_Y));
KC_INV_X4 T95 ( .Y(T95_Y), .A(T5186_Y));
KC_INV_X4 T111 ( .Y(T111_Y), .A(T104_Y));
KC_INV_X4 T193 ( .Y(T193_Y), .A(T6359_Q));
KC_INV_X4 T203 ( .Y(T203_Y), .A(T6355_Q));
KC_INV_X4 T462 ( .Y(T462_Y), .A(T481_Y));
KC_INV_X4 T470 ( .Y(T470_Y), .A(T469_Y));
KC_INV_X4 T537 ( .Y(T537_Y), .A(T539_Y));
KC_INV_X4 T580 ( .Y(T580_Y), .A(T534_Y));
KC_INV_X4 T795 ( .Y(T795_Y), .A(T5201_Y));
KC_INV_X4 T804 ( .Y(T804_Y), .A(T117_Y));
KC_INV_X4 T887 ( .Y(T887_Y), .A(T901_Y));
KC_INV_X4 T897 ( .Y(T897_Y), .A(T898_Y));
KC_INV_X4 T1179 ( .Y(T1179_Y), .A(T5235_Y));
KC_INV_X4 T1181 ( .Y(T1181_Y), .A(T1182_Y));
KC_INV_X4 T1226 ( .Y(T1226_Y), .A(T1233_Y));
KC_INV_X4 T1235 ( .Y(T1235_Y), .A(T1234_Y));
KC_INV_X4 T1388 ( .Y(T1388_Y), .A(T1387_Y));
KC_INV_X4 T1392 ( .Y(T1392_Y), .A(T1322_Y));
KC_INV_X4 T1454 ( .Y(T1454_Y), .A(T4888_Y));
KC_INV_X4 T1460 ( .Y(T1460_Y), .A(T5291_Y));
KC_INV_X4 T1529 ( .Y(T1529_Y), .A(T4894_Y));
KC_INV_X4 T1543 ( .Y(T1543_Y), .A(T1531_Y));
KC_INV_X4 T1577 ( .Y(T1577_Y), .A(T1573_Y));
KC_INV_X4 T1595 ( .Y(T1595_Y), .A(T1592_Y));
KC_INV_X4 T1868 ( .Y(T1868_Y), .A(T1871_Y));
KC_INV_X4 T1959 ( .Y(T1959_Y), .A(T5580_Y));
KC_INV_X4 T2409 ( .Y(T2409_Y), .A(T1865_Y));
KC_INV_X4 T2497 ( .Y(T2497_Y), .A(T5285_Y));
KC_INV_X4 T3009 ( .Y(T3009_Y), .A(T3008_Y));
KC_INV_X4 T3149 ( .Y(T3149_Y), .A(T5392_Y));
KC_INV_X4 T3156 ( .Y(T3156_Y), .A(T5398_Y));
KC_INV_X4 T3190 ( .Y(T3190_Y), .A(T3196_Y));
KC_INV_X4 T3197 ( .Y(T3197_Y), .A(T3195_Y));
KC_INV_X4 T3229 ( .Y(T3229_Y), .A(T3232_Y));
KC_INV_X4 T3243 ( .Y(T3243_Y), .A(T3240_Y));
KC_INV_X4 T3366 ( .Y(T3366_Y), .A(T3365_Y));
KC_INV_X4 T3407 ( .Y(T3407_Y), .A(T5073_Y));
KC_INV_X4 T3529 ( .Y(T3529_Y), .A(T3502_Y));
KC_INV_X4 T3532 ( .Y(T3532_Y), .A(T3535_Y));
KC_INV_X4 T3642 ( .Y(T3642_Y), .A(T5133_Y));
KC_INV_X4 T3646 ( .Y(T3646_Y), .A(T3649_Y));
KC_INV_X4 T3955 ( .Y(T3955_Y), .A(T3959_Y));
KC_INV_X4 T4193 ( .Y(T4193_Y), .A(T4185_Y));
KC_INV_X4 T4194 ( .Y(T4194_Y), .A(T4201_Y));
KC_INV_X4 T4206 ( .Y(T4206_Y), .A(T4209_Y));
KC_INV_X4 T4224 ( .Y(T4224_Y), .A(T4223_Y));
KC_INV_X4 T4327 ( .Y(T4327_Y), .A(T1497_Y));
KC_INV_X4 T4336 ( .Y(T4336_Y), .A(T4337_Y));
KC_INV_X4 T5117 ( .Y(T5117_Y), .A(T5475_Y));
KC_INV_X4 T5246 ( .Y(T5246_Y), .A(T5245_Y));
KC_OAI13_X3 T16167 ( .B0(T2807_Y), .A(T4981_Y), .B2(T2669_Q),     .Y(T16167_Y), .B1(T3242_Q));
KC_OAI13_X3 T15311 ( .B0(T886_Y), .A(T9331_Y), .B2(T6648_Y),     .Y(T15311_Y), .B1(T578_Y));
KC_NOR4_X1 T6247 ( .Y(T6247_Y), .D(T277_Q), .C(T284_Q), .B(T278_Q),     .A(T294_Q));
KC_NOR4_X1 T6246 ( .Y(T6246_Y), .D(T5205_Q), .C(T626_Q), .B(T443_Q),     .A(T5198_Q));
KC_NOR4_X1 T15766 ( .Y(T15766_Y), .D(T712_Q), .C(T5300_Q), .B(T705_Q),     .A(T710_Q));
KC_NOR4_X1 T16233 ( .Y(T16233_Y), .D(T12263_Y), .C(T16040_Y),     .B(T1365_Y), .A(T15529_Y));
KC_NOR4_X1 T15910 ( .Y(T15910_Y), .D(T3895_Q), .C(T3883_Q),     .B(T3877_Q), .A(T5129_Q));
KC_NOR4_X1 T15727 ( .Y(T15727_Y), .D(T9353_Q), .C(T5303_Q), .B(T522_Q),     .A(T363_Q));
KC_NOR4_X1 T15756 ( .Y(T15756_Y), .D(T5339_Y), .C(T6091_Y),     .B(T13323_Q), .A(T13324_Q));
KC_NOR4_X1 T15726 ( .Y(T15726_Y), .D(T184_Q), .C(T9354_Q), .B(T359_Q),     .A(T9355_Q));
KC_OAI13_X2 T16177 ( .B0(T15769_Y), .A(T8745_Y), .B2(T7676_Y),     .Y(T16177_Y), .B1(T15213_Y));
KC_OAI13_X2 T6597 ( .B0(T886_Y), .A(T7413_Y), .B2(T6685_Y),     .Y(T6597_Y), .B1(T384_Y));
KC_OAI13_X2 T9889 ( .B0(T2065_Y), .A(T5979_Y), .B2(T2560_Y),     .Y(T9889_Y), .B1(T2068_Y));
KC_OAI13_X2 T15739 ( .B0(T886_Y), .A(T7590_Y), .B2(T7585_Y),     .Y(T15739_Y), .B1(T7593_Y));
KC_OAI13_X2 T6801 ( .B0(T886_Y), .A(T7410_Y), .B2(T6798_Y),     .Y(T6801_Y), .B1(T15408_Y));
KC_OAI13_X2 T6799 ( .B0(T886_Y), .A(T7414_Y), .B2(T7355_Y),     .Y(T6799_Y), .B1(T6693_Y));
KC_OAI13_X2 T6445 ( .B0(T10389_Y), .A(T1419_Y), .B2(T16448_Y),     .Y(T6445_Y), .B1(T4884_Y));
KC_OAI13_X2 T6444 ( .B0(T15670_Y), .A(T1419_Y), .B2(T4884_Y),     .Y(T6444_Y), .B1(T9541_Y));
KC_OAI13_X2 T6818 ( .B0(T886_Y), .A(T7412_Y), .B2(T7407_Y),     .Y(T6818_Y), .B1(T15650_Y));
KC_ADD_C_X1 T6189 ( .B(T167_Q), .A(T6400_Y), .Y(T6189_Y), .C(T6233_Y));
KC_ADD_C_X1 T6724 ( .B(T182_Q), .A(T6410_Y), .Y(T6724_Y), .C(T6727_Y));
KC_ADD_C_X1 T1477 ( .B(T6465_Y), .A(T7071_Y), .Y(T1477_Y),     .C(T5237_Q));
KC_ADD_C_X1 T1487 ( .B(T157_Q), .A(T303_Y), .Y(T1487_Y), .C(T327_Y));
KC_ADD_C_X1 T6353 ( .B(T180_Q), .A(T307_Y), .Y(T6353_Y), .C(T6351_Y));
KC_ADD_C_X1 T6354 ( .B(T154_Q), .A(T300_Y), .Y(T6354_Y), .C(T6471_Y));
KC_ADD_C_X1 T6612 ( .B(T386_Y), .A(T6703_Y), .Y(T6612_Y), .C(T329_Q));
KC_ADD_C_X1 T6607 ( .B(T6608_Y), .A(T6714_Y), .Y(T6607_Y), .C(T326_Q));
KC_ADD_C_X1 T6602 ( .B(T164_Q), .A(T6603_Y), .Y(T6602_Y), .C(T6398_Y));
KC_ADD_C_X1 T6598 ( .B(T173_Q), .A(T389_Y), .Y(T6598_Y), .C(T6724_Y));
KC_ADD_C_X1 T6368 ( .B(T397_Y), .A(T6598_Y), .Y(T6368_Y), .C(T174_Q));
KC_ADD_C_X1 T6377 ( .B(T396_Y), .A(T6602_Y), .Y(T6377_Y), .C(T5263_Q));
KC_ADD_C_X1 T6378 ( .B(T6189_Y), .A(T399_Y), .Y(T6378_Y), .C(T169_Q));
KC_ADD_C_X1 T6714 ( .B(T165_Q), .A(T6723_Y), .Y(T6714_Y), .C(T6409_Y));
KC_ADD_C_X1 T6672 ( .B(T6681_Y), .A(T15725_Y), .Y(T6672_Y),     .C(T9355_Q));
KC_ADD_C_X1 T6389 ( .B(T505_Y), .A(T338_Y), .Y(T6389_Y), .C(T9354_Q));
KC_ADD_C_X1 T6390 ( .B(T5277_Q), .A(T349_Y), .Y(T6390_Y), .C(T506_Y));
KC_ADD_C_X1 T6398 ( .B(T335_Q), .A(T6389_Y), .Y(T6398_Y), .C(T535_Y));
KC_ADD_C_X1 T6409 ( .B(T344_Q), .A(T6672_Y), .Y(T6409_Y), .C(T568_Y));
KC_ADD_C_X1 T6410 ( .B(T507_Y), .A(T8675_Y), .Y(T6410_Y), .C(T5278_Q));
KC_ADD_C_X1 T16077 ( .B(T5228_Y), .A(T9174_Y), .Y(T16077_Y),     .C(T9199_Y));
KC_ADD_C_X1 T1498 ( .B(T155_Q), .A(T476_Y), .Y(T1498_Y), .C(T15371_Y));
KC_ADD_C_X1 T6347 ( .B(T179_Q), .A(T4834_Y), .Y(T6347_Y), .C(T381_Y));
KC_ADD_C_X1 T6618 ( .B(T6613_Y), .A(T6396_Y), .Y(T6618_Y),     .C(T5254_Q));
KC_ADD_C_X1 T6366 ( .B(T385_Y), .A(T6708_Y), .Y(T6366_Y), .C(T5261_Q));
KC_ADD_C_X1 T6375 ( .B(T391_Y), .A(T6706_Y), .Y(T6375_Y), .C(T489_Q));
KC_ADD_C_X1 T6376 ( .B(T4810_Q), .A(T486_Y), .Y(T6376_Y),     .C(T15389_Y));
KC_ADD_C_X1 T6708 ( .B(T664_Q), .A(T6712_Y), .Y(T6708_Y), .C(T6408_Y));
KC_ADD_C_X1 T6706 ( .B(T4799_Q), .A(T6713_Y), .Y(T6706_Y),     .C(T6405_Y));
KC_ADD_C_X1 T6663 ( .B(T6670_Y), .A(T9343_Y), .Y(T6663_Y), .C(T523_Q));
KC_ADD_C_X1 T6384 ( .B(T525_Q), .A(T6663_Y), .Y(T6384_Y), .C(T562_Y));
KC_ADD_C_X1 T6385 ( .B(T502_Y), .A(T509_Y), .Y(T6385_Y), .C(T9338_Q));
KC_ADD_C_X1 T6386 ( .B(T504_Y), .A(T508_Y), .Y(T6386_Y), .C(T359_Q));
KC_ADD_C_X1 T6396 ( .B(T4837_Q), .A(T527_Y), .Y(T6396_Y), .C(T6384_Y));
KC_ADD_C_X1 T6405 ( .B(T500_Q), .A(T6407_Y), .Y(T6405_Y),     .C(T15412_Y));
KC_ADD_C_X1 T6406 ( .B(T343_Q), .A(T6386_Y), .Y(T6406_Y), .C(T6397_Y));
KC_ADD_C_X1 T6407 ( .B(T564_Y), .A(T8662_Y), .Y(T6407_Y), .C(T360_Q));
KC_ADD_C_X1 T6408 ( .B(T5279_Q), .A(T6385_Y), .Y(T6408_Y), .C(T563_Y));
KC_ADD_C_X1 T2391 ( .B(T6172_Y), .A(T8604_Y), .Y(T2391_Y),     .C(T4854_Q));
KC_ADD_C_X1 T5804 ( .B(T15647_Y), .A(T8616_Y), .Y(T5804_Y),     .C(T828_Q));
KC_ADD_C_X1 T6372 ( .B(T15391_Y), .A(T8611_Y), .Y(T6372_Y),     .C(T5258_Q));
KC_ADD_C_X1 T6373 ( .B(T15390_Y), .A(T8584_Y), .Y(T6373_Y),     .C(T5259_Q));
KC_ADD_C_X1 T6374 ( .B(T379_Y), .A(T8569_Y), .Y(T6374_Y), .C(T861_Q));
KC_ADD_C_X1 T16068 ( .B(T5968_Y), .A(T12770_Y), .Y(T16068_Y),     .C(T3342_Y));
KC_ADD_C_X1 T6566 ( .B(T2317_Y), .A(T2358_Y), .Y(T6566_Y),     .C(T15638_Y));
KC_ADD_C_X1 T6501 ( .B(T6500_Y), .A(T6500_Y), .Y(T6501_Y),     .C(T2369_Y));
KC_ADD_C_X1 T15991 ( .B(T2782_Y), .A(T12241_Y), .Y(T15991_Y),     .C(T8280_Y));
KC_ADD_C_X1 T6413 ( .B(T9752_Y), .A(T9773_Y), .Y(T6413_Y),     .C(T11175_Y));
KC_ADD_C_X1 T6429 ( .B(T6846_Y), .A(T3681_Y), .Y(T6429_Y),     .C(T16230_Y));
KC_ADD_C_X1 T15823 ( .B(T6031_Co), .A(T5426_Y), .Y(T15823_Y),     .C(T15554_Y));
KC_ADD_C_X1 T15930 ( .B(T15128_Y), .A(T10927_Y), .Y(T15930_Y),     .C(T12185_Y));
KC_ADD_C_X1 T15963 ( .B(T9487_Y), .A(T4542_Y), .Y(T15963_Y),     .C(T4541_Y));
KC_ADD_C_X1 T15947 ( .B(T12209_Y), .A(T12197_Y), .Y(T15947_Y),     .C(T5884_Y));
KC_ADD_C_X1 T15986 ( .B(T15988_Y), .A(T4570_Y), .Y(T15986_Y),     .C(T11572_Y));
KC_ADD_C_X1 T511 ( .B(T153_Q), .A(T308_Y), .Y(T511_Y), .C(T15372_Y));
KC_ADD_C_X1 T6703 ( .B(T5252_Q), .A(T6609_Y), .Y(T6703_Y),     .C(T6406_Y));
KC_ADD_C_X1 T5782 ( .B(T5938_Y), .A(T8562_Y), .Y(T5782_Y),     .C(T5238_Q));
KC_ADD_C_X1 T6220 ( .B(T15387_Y), .A(T8592_Y), .Y(T6220_Y),     .C(T860_Q));
KC_ADD_C_X1 T16089 ( .B(T7779_Y), .A(T4919_Y), .Y(T16089_Y),     .C(T9781_Y));
KC_ADD_C_X1 T16095 ( .B(T2025_Y), .A(T2007_Y), .Y(T16095_Y),     .C(T2025_Y));
KC_ADD_C_X1 T6356 ( .B(T14969_Y), .A(T4962_Y), .Y(T6356_Y),     .C(T14969_Y));
KC_ADD_C_X1 T16093 ( .B(T634_Y), .A(T2478_Y), .Y(T16093_Y),     .C(T4986_Y));
KC_ADD_C_X1 T6400 ( .B(T183_Q), .A(T6728_Y), .Y(T6400_Y), .C(T6390_Y));
KC_NOR3_X2 T15195 ( .Y(T15195_Y), .B(T84_Q), .C(T5623_Y), .A(T98_Q));
KC_NOR3_X2 T15213 ( .Y(T15213_Y), .B(T647_Y), .C(T7678_Y), .A(T802_Y));
KC_NOR3_X2 T15223 ( .Y(T15223_Y), .B(T1133_Q), .C(T980_Q), .A(T946_Y));
KC_NOR3_X2 T15198 ( .Y(T15198_Y), .B(T3072_Y), .C(T7182_Y),     .A(T3071_Y));
KC_NOR3_X2 T15197 ( .Y(T15197_Y), .B(T2589_Y), .C(T10404_Y),     .A(T14980_Y));
KC_NOR3_X2 T15248 ( .Y(T15248_Y), .B(T2589_Y), .C(T5673_Y),     .A(T1338_Y));
KC_NOR3_X2 T15207 ( .Y(T15207_Y), .B(T3072_Y), .C(T5674_Y),     .A(T3071_Y));
KC_NOR3_X2 T15194 ( .Y(T15194_Y), .B(T5331_Y), .C(T7340_Y),     .A(T10788_Y));
KC_NOR3_X2 T15247 ( .Y(T15247_Y), .B(T5331_Y), .C(T5664_Y),     .A(T7323_Y));
KC_NOR3_X2 T15246 ( .Y(T15246_Y), .B(T3072_Y), .C(T5650_Y),     .A(T3071_Y));
KC_NOR3_X2 T15245 ( .Y(T15245_Y), .B(T2589_Y), .C(T5651_Y),     .A(T1545_Y));
KC_NOR3_X2 T15202 ( .Y(T15202_Y), .B(T5331_Y), .C(T5648_Y),     .A(T7323_Y));
KC_NOR3_X2 T15201 ( .Y(T15201_Y), .B(T3650_Y), .C(T7320_Y),     .A(T3653_Y));
KC_NOR3_X2 T15229 ( .Y(T15229_Y), .B(T5331_Y), .C(T10320_Y),     .A(T8011_Y));
KC_NOR3_X2 T15228 ( .Y(T15228_Y), .B(T2589_Y), .C(T8003_Y),     .A(T8000_Y));
KC_NOR3_X2 T15224 ( .Y(T15224_Y), .B(T3072_Y), .C(T8002_Y),     .A(T3071_Y));
KC_NOR3_X2 T15205 ( .Y(T15205_Y), .B(T3072_Y), .C(T7334_Y),     .A(T3071_Y));
KC_NOR3_X2 T15221 ( .Y(T15221_Y), .B(T16447_Y), .C(T2500_Y),     .A(T16195_Y));
KC_NOR3_X2 T15220 ( .Y(T15220_Y), .B(T2861_Y), .C(T2501_Y),     .A(T5021_Y));
KC_NOR3_X2 T15218 ( .Y(T15218_Y), .B(T16447_Y), .C(T2502_Y),     .A(T16195_Y));
KC_NOR3_X2 T15232 ( .Y(T15232_Y), .B(T11633_Y), .C(T6039_Y),     .A(T6086_Y));
KC_NOR3_X2 T15233 ( .Y(T15233_Y), .B(T15636_Y), .C(T10881_Y),     .A(T2936_Y));
KC_NOR3_X2 T15212 ( .Y(T15212_Y), .B(T3072_Y), .C(T3014_Y),     .A(T3071_Y));
KC_NOR3_X2 T15211 ( .Y(T15211_Y), .B(T2589_Y), .C(T3013_Y),     .A(T3610_Y));
KC_NOR3_X2 T15234 ( .Y(T15234_Y), .B(T3510_Y), .C(T3512_Y),     .A(T3523_Q));
KC_NOR3_X2 T15256 ( .Y(T15256_Y), .B(T5331_Y), .C(T3607_Y),     .A(T5088_Y));
KC_NOR3_X2 T15222 ( .Y(T15222_Y), .B(T5331_Y), .C(T3651_Y),     .A(T16063_Y));
KC_NOR3_X2 T15219 ( .Y(T15219_Y), .B(T2589_Y), .C(T3654_Y),     .A(T3635_Y));
KC_NOR3_X2 T15216 ( .Y(T15216_Y), .B(T3081_Y), .C(T3667_Y),     .A(T3080_Y));
KC_NOR3_X2 T15215 ( .Y(T15215_Y), .B(T2589_Y), .C(T3668_Y),     .A(T3684_Y));
KC_NOR3_X2 T15214 ( .Y(T15214_Y), .B(T3677_Y), .C(T3666_Y),     .A(T3676_Y));
KC_NOR3_X2 T15254 ( .Y(T15254_Y), .B(T5331_Y), .C(T5082_Y),     .A(T3719_Y));
KC_NOR3_X2 T15253 ( .Y(T15253_Y), .B(T3677_Y), .C(T3712_Y),     .A(T3676_Y));
KC_NOR3_X2 T15231 ( .Y(T15231_Y), .B(T5862_Y), .C(T10631_Y),     .A(T15570_Y));
KC_NOR3_X2 T15244 ( .Y(T15244_Y), .B(T3650_Y), .C(T7351_Y),     .A(T3653_Y));
KC_NOR3_X2 T15237 ( .Y(T15237_Y), .B(T5331_Y), .C(T7350_Y),     .A(T7337_Y));
KC_NOR3_X2 T15235 ( .Y(T15235_Y), .B(T3650_Y), .C(T5663_Y),     .A(T3653_Y));
KC_NOR3_X2 T15251 ( .Y(T15251_Y), .B(T3677_Y), .C(T3608_Y),     .A(T3676_Y));
KC_NOR3_X2 T15204 ( .Y(T15204_Y), .B(T2589_Y), .C(T7322_Y),     .A(T1545_Y));
KC_NOR3_X2 T15217 ( .Y(T15217_Y), .B(T3081_Y), .C(T3069_Y),     .A(T3080_Y));
KC_NAND4_X2 T12368 ( .D(T114_Q), .C(T103_Q), .B(T5203_Q), .A(T8543_Y),     .Y(T12368_Y));
KC_NAND4_X2 T16176 ( .D(T743_Y), .C(T15430_Y), .B(T7581_Y), .A(T207_Q),     .Y(T16176_Y));
KC_NAND4_X2 T12446 ( .D(T8863_Y), .C(T15429_Y), .B(T8790_Y),     .A(T7676_Y), .Y(T12446_Y));
KC_NAND4_X2 T15903 ( .D(T12155_Y), .C(T2702_Y), .B(T5380_Q),     .A(T16301_Q), .Y(T15903_Y));
KC_NAND4_X2 T12357 ( .D(T15857_Y), .C(T2719_Y), .B(T15797_Q),     .A(T5380_Q), .Y(T12357_Y));
KC_NAND4_X2 T6511 ( .D(T6490_Y), .C(T11833_Y), .B(T3523_Q),     .A(T3525_Q), .Y(T6511_Y));
KC_NAND4_X2 T12064 ( .D(T6512_Y), .C(T11843_Y), .B(T8150_Y),     .A(T3525_Q), .Y(T12064_Y));
KC_NAND4_X2 T16050 ( .D(T6043_Y), .C(T5070_Y), .B(T11656_Y),     .A(T11638_Y), .Y(T16050_Y));
KC_NAND4_X2 T12089 ( .D(T9961_Y), .C(T4288_Y), .B(T4301_Y),     .A(T4287_Y), .Y(T12089_Y));
KC_NAND4_X2 T12442 ( .D(T743_Y), .C(T7695_Y), .B(T5192_Q), .A(T566_Q),     .Y(T12442_Y));
KC_DFFSNHQ_X3 T16482 ( .CK(T14960_Q), .D(T2088_Y), .Q(T16482_Q),     .SN(T15011_Y));
KC_DFFSNHQ_X3 T16480 ( .CK(T352_Y), .D(T11236_Y), .Q(T16480_Q),     .SN(T14976_Y));
KC_DFFRNHQ_X4 T16462 ( .Q(T16462_Q), .CK1(T1727_Y), .D(T1729_Q),     .RN(T15003_Y), .CK(T1604_Y));
KC_DFFRNHQ_X4 T16461 ( .Q(T16461_Q), .CK1(T2048_Y), .D(T2056_Y),     .RN(T10083_Y), .CK(T14967_Y));
KC_DFFRNHQ_X4 T16469 ( .Q(T16469_Q), .CK1(T16156_Y), .D(T15004_Y),     .RN(T15011_Y), .CK(T14557_Q));
KC_DFFRNHQ_X4 T16471 ( .Q(T16471_Q), .CK1(T16156_Y), .D(T16469_Q),     .RN(T15011_Y), .CK(T14557_Q));
KC_DFFRNHQ_X4 T16458 ( .Q(T16458_Q), .CK1(T11726_Y), .D(T12317_Y),     .RN(T15021_Y), .CK(T4045_Y));
KC_DFFRNHQ_X4 T16455 ( .Q(T16455_Q), .CK1(T4008_Y), .D(T4063_Y),     .RN(T15035_Y), .CK(T4045_Y));
KC_DFFRNHQ_X4 T16454 ( .Q(T16454_Q), .CK1(T5126_Y), .D(T6469_Y),     .RN(T15035_Y), .CK(T4045_Y));
KC_DFFRNHQ_X4 T16453 ( .Q(T16453_Q), .CK1(T4007_Y), .D(T6469_Y),     .RN(T15035_Y), .CK(T4045_Y));
KC_DFFRNHQ_X4 T16457 ( .Q(T16457_Q), .CK1(T10960_Y), .D(T8503_Y),     .RN(T15035_Y), .CK(T14575_Q));
KC_DFFRNHQ_X4 T16466 ( .Q(T16466_Q), .CK1(T4536_Y), .D(T10931_Y),     .RN(T3888_Y), .CK(T3879_Y));
KC_DFFRNHQ_X4 T16460 ( .Q(T16460_Q), .CK1(T12868_Y), .D(T11786_Y),     .RN(T15022_Y), .CK(T4728_Y));
KC_DFFRNHQ_X4 T16459 ( .Q(T16459_Q), .CK1(T5151_Y), .D(T16144_Y),     .RN(T15022_Y), .CK(T2736_Y));
KC_DFFRNHQ_X4 T16465 ( .Q(T16465_Q), .CK1(T1102_Y), .D(T7837_Y),     .RN(T2019_Y), .CK(T2667_Y));
KC_OA22_X1 T16119 ( .A1(T8024_Y), .B0(T9925_Y), .B1(T9895_Y),     .A0(T8023_Y), .Y(T16119_Y));
KC_OA22_X1 T16126 ( .A1(T10042_Y), .B0(T10002_Y), .B1(T1481_Y),     .A0(T9917_Y), .Y(T16126_Y));
KC_OA22_X1 T15846 ( .A1(T4436_Y), .B0(T3840_Y), .B1(T3797_Y),     .A0(T5780_Y), .Y(T15846_Y));
KC_OA22_X1 T15833 ( .A1(T5806_Y), .B0(T3816_Y), .B1(T5101_Y),     .A0(T5780_Y), .Y(T15833_Y));
KC_OA22_X1 T15898 ( .A1(T11408_Y), .B0(T4440_Y), .B1(T3827_Y),     .A0(T5840_Y), .Y(T15898_Y));
KC_OA22_X1 T16128 ( .A1(T10580_Y), .B0(T11710_Y), .B1(T4083_Y),     .A0(T6517_Y), .Y(T16128_Y));
KC_OA22_X1 T16118 ( .A1(T7948_Y), .B0(T10313_Y), .B1(T9914_Y),     .A0(T10314_Y), .Y(T16118_Y));
KC_OA12B_X1 T60 ( .Y(T60_Y), .C(T12470_Y), .A(T12472_Y), .B(T12471_Y));
KC_OA12B_X1 T15816 ( .Y(T15816_Y), .C(T16285_Y), .A(T9072_Y),     .B(T9069_Y));
KC_OA12B_X1 T16408 ( .Y(T16408_Y), .C(T13250_Y), .A(T756_Y),     .B(T8945_Y));
KC_OA12B_X1 T15770 ( .Y(T15770_Y), .C(T791_Y), .A(T7646_Y),     .B(T7844_Y));
KC_OA12B_X1 T15763 ( .Y(T15763_Y), .C(T791_Y), .A(T7563_Y),     .B(T7844_Y));
KC_OA12B_X1 T15941 ( .Y(T15941_Y), .C(T11531_Y), .A(T11532_Y),     .B(T6191_Y));
KC_OA12B_X1 T15814 ( .Y(T15814_Y), .C(T16268_Y), .A(T2029_Y),     .B(T2032_Y));
KC_OA12B_X1 T15812 ( .Y(T15812_Y), .C(T2035_Y), .A(T1721_Y),     .B(T1720_Y));
KC_OA12B_X1 T16057 ( .Y(T16057_Y), .C(T11029_Y), .A(T16305_Y),     .B(T2841_Q));
KC_OA12B_X1 T15961 ( .Y(T15961_Y), .C(T3918_Y), .A(T11024_Y),     .B(T11534_Y));
KC_OA12B_X1 T6589 ( .Y(T6589_Y), .C(T11779_Y), .A(T10989_Y),     .B(T4704_Y));
KC_OA12B_X1 T15993 ( .Y(T15993_Y), .C(T2757_Y), .A(T5477_Y),     .B(T8271_Y));
KC_OA12B_X1 T15767 ( .Y(T15767_Y), .C(T791_Y), .A(T7644_Y),     .B(T7844_Y));
KC_OA12B_X1 T16094 ( .Y(T16094_Y), .C(T1102_Y), .A(T5025_Q),     .B(T15843_Y));
KC_AOI22B_X1 T16312 ( .A0N(T7574_Y), .B0(T16331_Y), .B1(T797_Y),     .Y(T16312_Y), .A1(T7832_Y));
KC_AOI22B_X1 T6428 ( .A0N(T7669_Y), .B0(T16329_Y), .B1(T642_Y),     .Y(T6428_Y), .A1(T7822_Y));
KC_AOI22B_X1 T15794 ( .A0N(T16390_Y), .B0(T1334_Y), .B1(T1287_Y),     .Y(T15794_Y), .A1(T8081_Y));
KC_AOI22B_X1 T15793 ( .A0N(T7910_Y), .B0(T1272_Y), .B1(T1217_Y),     .Y(T15793_Y), .A1(T8080_Y));
KC_AOI22B_X1 T704 ( .A0N(T273_Q), .B0(T281_Q), .B1(T347_Y), .Y(T704_Y),     .A1(T272_Q));
KC_AOI22B_X1 T6395 ( .A0N(T4799_Q), .B0(T9339_Q), .B1(T499_Y),     .Y(T6395_Y), .A1(T664_Q));
KC_AOI22B_X1 T15801 ( .A0N(T8127_Y), .B0(T1421_Y), .B1(T9046_S),     .Y(T15801_Y), .A1(T966_Y));
KC_AOI22B_X1 T6245 ( .A0N(T453_Q), .B0(T6272_Y), .B1(T13270_Y),     .Y(T6245_Y), .A1(T5205_Q));
KC_AOI22B_X1 T1442 ( .A0N(T276_Q), .B0(T330_Q), .B1(T391_Y),     .Y(T1442_Y), .A1(T5196_Q));
KC_AOI22B_X1 T6403 ( .A0N(T5280_Q), .B0(T181_Q), .B1(T15412_Y),     .Y(T6403_Y), .A1(T7367_Q));
KC_AOI22B_X1 T6394 ( .A0N(T695_Q), .B0(T663_Q), .B1(T6699_Y),     .Y(T6394_Y), .A1(T687_Q));
KC_AOI22B_X1 T6427 ( .A0N(T716_Q), .B0(T741_Q), .B1(T9378_Y),     .Y(T6427_Y), .A1(T713_Q));
KC_AOI22B_X1 T15785 ( .A0N(T8942_Y), .B0(T8860_Y), .B1(T905_Y),     .Y(T15785_Y), .A1(T8859_Y));
KC_AOI22B_X1 T15784 ( .A0N(T9010_Y), .B0(T8860_Y), .B1(T932_Y),     .Y(T15784_Y), .A1(T8859_Y));
KC_AOI22B_X1 T15742 ( .A0N(T9316_Y), .B0(T692_Y), .B1(T15722_Y),     .Y(T15742_Y), .A1(T16440_Y));
KC_AOI22B_X1 T15741 ( .A0N(T9318_Y), .B0(T692_Y), .B1(T7385_Y),     .Y(T15741_Y), .A1(T16440_Y));
KC_AOI22B_X1 T15738 ( .A0N(T15740_Y), .B0(T9313_Y), .B1(T7385_Y),     .Y(T15738_Y), .A1(T16440_Y));
KC_AOI22B_X1 T6798 ( .A0N(T11087_Y), .B0(T15223_Y), .B1(T1039_Y),     .Y(T6798_Y), .A1(T715_Y));
KC_AOI22B_X1 T6380 ( .A0N(T6835_Y), .B0(T9334_Y), .B1(T7385_Y),     .Y(T6380_Y), .A1(T16440_Y));
KC_AOI22B_X1 T15799 ( .A0N(T16278_Y), .B0(T9431_Y), .B1(T1157_Q),     .Y(T15799_Y), .A1(T7809_Y));
KC_AOI22B_X1 T15811 ( .A0N(T2034_Y), .B0(T5363_Q), .B1(T4935_Y),     .Y(T15811_Y), .A1(T2628_Q));
KC_AOI22B_X1 T16172 ( .A0N(T15815_Q), .B0(T10251_Y), .B1(T15552_Y),     .Y(T16172_Y), .A1(T10244_Y));
KC_AOI22B_X1 T6564 ( .A0N(T5109_Y), .B0(T10553_Y), .B1(T12106_Y),     .Y(T6564_Y), .A1(T10550_Y));
KC_AOI22B_X1 T15836 ( .A0N(T4436_Y), .B0(T11379_Y), .B1(T11322_Y),     .Y(T15836_Y), .A1(T11985_Y));
KC_AOI22B_X1 T15757 ( .A0N(T11787_Y), .B0(T4732_Y), .B1(T4700_Y),     .Y(T15757_Y), .A1(T4704_Y));
KC_AOI22B_X1 T6402 ( .A0N(T6803_Y), .B0(T9312_Y), .B1(T7385_Y),     .Y(T6402_Y), .A1(T16440_Y));
KC_AOI22B_X1 T6382 ( .A0N(T124_Q), .B0(T9313_Y), .B1(T15722_Y),     .Y(T6382_Y), .A1(T16440_Y));
KC_AOI22B_X1 T6381 ( .A0N(T6819_Y), .B0(T9312_Y), .B1(T15722_Y),     .Y(T6381_Y), .A1(T16440_Y));
KC_AOI22B_X1 T6414 ( .A0N(T4840_Q), .B0(T716_Q), .B1(T912_Y),     .Y(T6414_Y), .A1(T5346_Q));
KC_AOI22B_X1 T16383 ( .A0N(T953_Y), .B0(T1127_Q), .B1(T951_Y),     .Y(T16383_Y), .A1(T15454_Y));
KC_AOI22B_X1 T15790 ( .A0N(T9415_Y), .B0(T8860_Y), .B1(T916_Y),     .Y(T15790_Y), .A1(T8859_Y));
KC_AOI22B_X1 T15783 ( .A0N(T9407_Y), .B0(T8860_Y), .B1(T15434_Y),     .Y(T15783_Y), .A1(T8859_Y));
KC_AND2_X3 T15241 ( .B(T1431_Y), .A(T12915_Y), .Y(T15241_Y));
KC_AND2_X3 T15240 ( .B(T1431_Y), .A(T12913_Y), .Y(T15240_Y));
KC_AND2_X3 T15239 ( .B(T1431_Y), .A(T12914_Y), .Y(T15239_Y));
KC_AND2_X3 T15238 ( .B(T1431_Y), .A(T12502_Y), .Y(T15238_Y));
KC_AND2_X3 T15196 ( .B(T1431_Y), .A(T12503_Y), .Y(T15196_Y));
KC_AND2_X3 T15210 ( .B(T1431_Y), .A(T12545_Y), .Y(T15210_Y));
KC_AND2_X3 T15209 ( .B(T1431_Y), .A(T12530_Y), .Y(T15209_Y));
KC_AND2_X3 T15206 ( .B(T4885_Y), .A(T12543_Y), .Y(T15206_Y));
KC_AND2_X3 T15203 ( .B(T1431_Y), .A(T12539_Y), .Y(T15203_Y));
KC_AND2_X3 T15236 ( .B(T1418_Y), .A(T12917_Y), .Y(T15236_Y));
KC_AND2_X3 T15208 ( .B(T1431_Y), .A(T12535_Y), .Y(T15208_Y));
KC_AND2_X3 T15226 ( .B(T1491_Y), .A(T12617_Y), .Y(T15226_Y));
KC_AND2_X3 T15225 ( .B(T1491_Y), .A(T12681_Y), .Y(T15225_Y));
KC_AND2_X3 T15249 ( .B(T2452_Y), .A(T12929_Y), .Y(T15249_Y));
KC_AND2_X3 T15200 ( .B(T2452_Y), .A(T12552_Y), .Y(T15200_Y));
KC_AND2_X3 T15230 ( .B(T5745_Y), .A(T15806_Q), .Y(T15230_Y));
KC_AND2_X3 T15199 ( .B(T3025_Y), .A(T12566_Y), .Y(T15199_Y));
KC_AND2_X3 T15252 ( .B(T2651_Y), .A(T12930_Y), .Y(T15252_Y));
KC_AND2_X3 T15243 ( .B(T1431_Y), .A(T12911_Y), .Y(T15243_Y));
KC_AND2_X3 T15242 ( .B(T1431_Y), .A(T12912_Y), .Y(T15242_Y));
KC_AND2_X3 T15255 ( .B(T2525_Q), .A(T15443_Y), .Y(T15255_Y));
KC_AND2_X3 T15250 ( .B(T2452_Y), .A(T12926_Y), .Y(T15250_Y));
KC_AND2_X3 T15193 ( .B(T4885_Y), .A(T12537_Y), .Y(T15193_Y));
KC_AND2_X3 T15227 ( .B(T1491_Y), .A(T12685_Y), .Y(T15227_Y));
KC_AOI21B_X1 T121 ( .A0N(T12367_Y), .Y(T121_Y), .B(T12470_Y),     .A1(T8557_Y));
KC_AOI21B_X1 T122 ( .A0N(T5601_Y), .Y(T122_Y), .B(T12470_Y),     .A1(T126_Y));
KC_AOI21B_X1 T210 ( .A0N(T211_Q), .Y(T210_Y), .B(T7682_Y),     .A1(T16176_Y));
KC_AOI21B_X1 T220 ( .A0N(T7681_Y), .Y(T220_Y), .B(T12608_Y),     .A1(T9390_Y));
KC_AOI21B_X1 T230 ( .A0N(T9382_Y), .Y(T230_Y), .B(T9393_Y),     .A1(T9414_Y));
KC_AOI21B_X1 T899 ( .A0N(T7410_Y), .Y(T899_Y), .B(T16425_Y),     .A1(T689_Q));
KC_AOI21B_X1 T929 ( .A0N(T7645_Y), .Y(T929_Y), .B(T791_Y),     .A1(T928_Y));
KC_AOI21B_X1 T1248 ( .A0N(T7951_Y), .Y(T1248_Y), .B(T10170_Y),     .A1(T10315_Y));
KC_AOI21B_X1 T1369 ( .A0N(T10724_Y), .Y(T1369_Y), .B(T1371_Y),     .A1(T4825_Y));
KC_AOI21B_X1 T1370 ( .A0N(T1371_Y), .Y(T1370_Y), .B(T1371_Y),     .A1(T1368_Y));
KC_AOI21B_X1 T1563 ( .A0N(T9782_Y), .Y(T1563_Y), .B(T10756_Y),     .A1(T15662_Y));
KC_AOI21B_X1 T2003 ( .A0N(T6687_Y), .Y(T2003_Y), .B(T6686_S),     .A1(T2599_Y));
KC_AOI21B_X1 T2061 ( .A0N(T12734_Y), .Y(T2061_Y), .B(T12737_Y),     .A1(T2058_Y));
KC_AOI21B_X1 T2347 ( .A0N(T16129_Y), .Y(T2347_Y), .B(T6588_Y),     .A1(T2343_Y));
KC_AOI21B_X1 T2387 ( .A0N(T8432_Y), .Y(T2387_Y), .B(T6502_Y),     .A1(T8433_Y));
KC_AOI21B_X1 T2396 ( .A0N(T6492_Y), .Y(T2396_Y), .B(T2366_Y),     .A1(T8436_Y));
KC_AOI21B_X1 T2588 ( .A0N(T2572_Q), .Y(T2588_Y), .B(T15843_Y),     .A1(T2520_Y));
KC_AOI21B_X1 T2712 ( .A0N(T2703_Y), .Y(T2712_Y), .B(T8198_Y),     .A1(T15886_Y));
KC_AOI21B_X1 T2783 ( .A0N(T2791_Y), .Y(T2783_Y), .B(T6295_Y),     .A1(T5877_Y));
KC_AOI21B_X1 T2810 ( .A0N(T2811_Y), .Y(T2810_Y), .B(T16003_Y),     .A1(T16456_Y));
KC_AOI21B_X1 T2834 ( .A0N(T8469_Y), .Y(T2834_Y), .B(T11662_Y),     .A1(T8346_Y));
KC_AOI21B_X1 T2877 ( .A0N(T10594_Y), .Y(T2877_Y), .B(T16132_Y),     .A1(T5518_Y));
KC_AOI21B_X1 T2919 ( .A0N(T8515_Y), .Y(T2919_Y), .B(T6579_Y),     .A1(T11741_Y));
KC_AOI21B_X1 T3259 ( .A0N(T3262_Y), .Y(T3259_Y), .B(T3250_Y),     .A1(T15857_Y));
KC_AOI21B_X1 T3341 ( .A0N(T3328_Y), .Y(T3341_Y), .B(T5964_Y),     .A1(T3363_Y));
KC_AOI21B_X1 T3450 ( .A0N(T10975_Y), .Y(T3450_Y), .B(T12877_Y),     .A1(T3429_Y));
KC_AOI21B_X1 T3920 ( .A0N(T3913_Y), .Y(T3920_Y), .B(T11587_Y),     .A1(T5981_Y));
KC_AOI21B_X1 T3972 ( .A0N(T3883_Q), .Y(T3972_Y), .B(T3950_Y),     .A1(T6352_Y));
KC_AOI21B_X1 T4011 ( .A0N(T4042_Y), .Y(T4011_Y), .B(T5995_Y),     .A1(T15610_Y));
KC_AOI21B_X1 T4103 ( .A0N(T4071_Y), .Y(T4103_Y), .B(T6148_Y),     .A1(T4691_Y));
KC_AOI21B_X1 T4564 ( .A0N(T4563_Y), .Y(T4564_Y), .B(T4543_Y),     .A1(T15966_Y));
KC_AOI21B_X1 T4604 ( .A0N(T12017_Y), .Y(T4604_Y), .B(T2757_Y),     .A1(T10956_Y));
KC_AOI21B_X1 T4615 ( .A0N(T9486_Y), .Y(T4615_Y), .B(T3982_Y),     .A1(T9486_Y));
KC_AOI21B_X1 T4616 ( .A0N(T6326_Y), .Y(T4616_Y), .B(T4614_Y),     .A1(T5485_Y));
KC_AOI21B_X1 T4689 ( .A0N(T4687_Y), .Y(T4689_Y), .B(T4661_Y),     .A1(T4661_Y));
KC_AOI21B_X1 T5013 ( .A0N(T5999_Y), .Y(T5013_Y), .B(T2812_Y),     .A1(T12064_Y));
KC_AOI21B_X1 T5014 ( .A0N(T5009_Y), .Y(T5014_Y), .B(T2812_Y),     .A1(T12064_Y));
KC_AOI21B_X1 T5069 ( .A0N(T8345_Y), .Y(T5069_Y), .B(T11640_Y),     .A1(T5059_Y));
KC_AOI21B_X1 T5119 ( .A0N(T3918_Y), .Y(T5119_Y), .B(T11587_Y),     .A1(T5989_Y));
KC_AOI21B_X1 T5289 ( .A0N(T9786_Y), .Y(T5289_Y), .B(T16089_Y),     .A1(T7778_Y));
KC_AOI21B_X1 T5344 ( .A0N(T7916_Y), .Y(T5344_Y), .B(T7913_Y),     .A1(T7916_Y));
KC_AOI21B_X1 T5347 ( .A0N(T9400_Y), .Y(T5347_Y), .B(T8936_Y),     .A1(T5353_Q));
KC_XOR2_X5 T7914 ( .B(T15146_Y), .A(T8971_Y), .Y(T7914_Y));
KC_XOR2_X5 T7920 ( .B(T8883_Y), .A(T8881_Y), .Y(T7920_Y));
KC_XOR2_X5 T7874 ( .B(T8841_Y), .A(T8787_Y), .Y(T7874_Y));
KC_XOR2_X5 T7865 ( .B(T8823_Y), .A(T8840_Y), .Y(T7865_Y));
KC_XOR2_X5 T7864 ( .B(T8843_Y), .A(T8826_Y), .Y(T7864_Y));
KC_XOR2_X5 T8092 ( .B(T8968_Y), .A(T8959_Y), .Y(T8092_Y));
KC_XOR2_X5 T8091 ( .B(T16064_Y), .A(T8969_Y), .Y(T8091_Y));
KC_XOR2_X5 T8090 ( .B(T8970_Y), .A(T8967_Y), .Y(T8090_Y));
KC_XOR2_X5 T8089 ( .B(T8886_Y), .A(T8966_Y), .Y(T8089_Y));
KC_XOR2_X5 T8056 ( .B(T8926_Y), .A(T8927_Y), .Y(T8056_Y));
KC_XOR2_X5 T8055 ( .B(T8915_Y), .A(T8925_Y), .Y(T8055_Y));
KC_XOR2_X5 T9139 ( .B(T5336_Y), .A(T9134_Y), .Y(T9139_Y));
KC_XOR2_X5 T15084 ( .B(T9090_Y), .A(T9218_Y), .Y(T15084_Y));
KC_XOR2_X5 T9020 ( .B(T387_Y), .A(T9205_Y), .Y(T9020_Y));
KC_XOR2_X5 T9019 ( .B(T9023_Y), .A(T9209_Y), .Y(T9019_Y));
KC_XOR2_X5 T9018 ( .B(T9074_Y), .A(T9214_Y), .Y(T9018_Y));
KC_XOR2_X5 T9017 ( .B(T9022_Y), .A(T9201_Y), .Y(T9017_Y));
KC_XOR2_X5 T8136 ( .B(T8149_Y), .A(T9217_Y), .Y(T8136_Y));
KC_XOR2_X5 T8108 ( .B(T8146_Y), .A(T9208_Y), .Y(T8108_Y));
KC_XOR2_X5 T8107 ( .B(T8985_Y), .A(T9202_Y), .Y(T8107_Y));
KC_XOR2_X5 T8098 ( .B(T8988_Y), .A(T9249_Y), .Y(T8098_Y));
KC_XOR2_X5 T8087 ( .B(T8144_Y), .A(T9204_Y), .Y(T8087_Y));
KC_XOR2_X5 T8086 ( .B(T8145_Y), .A(T9215_Y), .Y(T8086_Y));
KC_XOR2_X5 T9149 ( .B(T9151_Y), .A(T9238_Y), .Y(T9149_Y));
KC_XOR2_X5 T9148 ( .B(T9152_Y), .A(T9216_Y), .Y(T9148_Y));
KC_XOR2_X5 T9068 ( .B(T9076_Y), .A(T9236_Y), .Y(T9068_Y));
KC_XOR2_X5 T9067 ( .B(T419_Y), .A(T9491_Y), .Y(T9067_Y));
KC_XOR2_X5 T9066 ( .B(T9075_Y), .A(T9179_Y), .Y(T9066_Y));
KC_XOR2_X5 T9241 ( .B(T9463_Y), .A(T16508_Y), .Y(T9241_Y));
KC_XOR2_X5 T1274 ( .B(T16171_Y), .A(T13054_Q), .Y(T1274_Y));
KC_XOR2_X5 T10032 ( .B(T1724_Y), .A(T16440_Y), .Y(T10032_Y));
KC_XOR2_X5 T2200 ( .B(T2670_Y), .A(T2249_Q), .Y(T2200_Y));
KC_XOR2_X5 T2207 ( .B(T2673_Y), .A(T2281_Q), .Y(T2207_Y));
KC_XOR2_X5 T2219 ( .B(T16069_Y), .A(T16010_Q), .Y(T2219_Y));
KC_XOR2_X5 T2220 ( .B(T2671_Y), .A(T2835_Q), .Y(T2220_Y));
KC_XOR2_X5 T2295 ( .B(T10612_Y), .A(T2311_Q), .Y(T2295_Y));
KC_XOR2_X5 T3185 ( .B(T15815_Q), .A(T4381_Q), .Y(T3185_Y));
KC_XOR2_X5 T9498 ( .B(T5284_Y), .A(T9494_Y), .Y(T9498_Y));
KC_XOR2_X5 T2714 ( .B(T11730_Y), .A(T15138_Q), .Y(T2714_Y));
KC_XOR2_X5 T10305 ( .B(T15660_Y), .A(T1471_Y), .Y(T10305_Y));
KC_XOR2_X5 T8143 ( .B(T8986_Y), .A(T9211_Y), .Y(T8143_Y));
KC_BUF_X8 T14983 ( .Y(T14983_Y), .A(T943_Y));
KC_BUF_X8 T16415 ( .Y(T16415_Y), .A(T991_Y));
KC_BUF_X8 T14964 ( .Y(T14964_Y), .A(T2083_Y));
KC_BUF_X8 T14982 ( .Y(T14982_Y), .A(T4841_Y));
KC_BUF_X8 T869 ( .Y(T869_Y), .A(T15230_Y));
KC_BUF_X8 T14998 ( .Y(T14998_Y), .A(T1598_Y));
KC_AND2_X1 T6852 ( .B(T15330_Y), .A(T13211_Y), .Y(T6852_Y));
KC_AND2_X1 T6851 ( .B(T15326_Y), .A(T13211_Y), .Y(T6851_Y));
KC_AND2_X1 T5583 ( .B(T15326_Y), .A(T13211_Y), .Y(T5583_Y));
KC_AND2_X1 T5635 ( .B(T13317_Y), .A(T13211_Y), .Y(T5635_Y));
KC_AND2_X1 T5626 ( .B(T13317_Y), .A(T13211_Y), .Y(T5626_Y));
KC_AND2_X1 T5632 ( .B(T15322_Y), .A(T13211_Y), .Y(T5632_Y));
KC_AND2_X1 T5638 ( .B(T15322_Y), .A(T13211_Y), .Y(T5638_Y));
KC_AND2_X1 T7405 ( .B(T195_Y), .A(T1283_RN), .Y(T7405_Y));
KC_AND2_X1 T7608 ( .B(T203_Y), .A(T193_Y), .Y(T7608_Y));
KC_AND2_X1 T8141 ( .B(T1339_Y), .A(T1428_Y), .Y(T8141_Y));
KC_AND2_X1 T5224 ( .B(T5274_Y), .A(T9199_Y), .Y(T5224_Y));
KC_AND2_X1 T7101 ( .B(T15370_Y), .A(T662_Y), .Y(T7101_Y));
KC_AND2_X1 T7094 ( .B(T15370_Y), .A(T662_Y), .Y(T7094_Y));
KC_AND2_X1 T8068 ( .B(T15657_Y), .A(T662_Y), .Y(T8068_Y));
KC_AND2_X1 T8043 ( .B(T15657_Y), .A(T662_Y), .Y(T8043_Y));
KC_AND2_X1 T7889 ( .B(T15485_Y), .A(T1597_Y), .Y(T7889_Y));
KC_AND2_X1 T7184 ( .B(T15672_Y), .A(T662_Y), .Y(T7184_Y));
KC_AND2_X1 T7353 ( .B(T15672_Y), .A(T662_Y), .Y(T7353_Y));
KC_AND2_X1 T7408 ( .B(T15410_Y), .A(T662_Y), .Y(T7408_Y));
KC_AND2_X1 T10755 ( .B(T15499_Y), .A(T1505_Y), .Y(T10755_Y));
KC_AND2_X1 T10722 ( .B(T15499_Y), .A(T1505_Y), .Y(T10722_Y));
KC_AND2_X1 T10659 ( .B(T16118_Y), .A(T2073_Y), .Y(T10659_Y));
KC_AND2_X1 T10740 ( .B(T1127_Q), .A(T2073_Y), .Y(T10740_Y));
KC_AND2_X1 T6873 ( .B(T15345_Y), .A(T1929_Y), .Y(T6873_Y));
KC_AND2_X1 T6871 ( .B(T15345_Y), .A(T1929_Y), .Y(T6871_Y));
KC_AND2_X1 T7539 ( .B(T15416_Y), .A(T1505_Y), .Y(T7539_Y));
KC_AND2_X1 T10739 ( .B(T16119_Y), .A(T2073_Y), .Y(T10739_Y));
KC_AND2_X1 T7129 ( .B(T15376_Y), .A(T1929_Y), .Y(T7129_Y));
KC_AND2_X1 T7128 ( .B(T15376_Y), .A(T1929_Y), .Y(T7128_Y));
KC_AND2_X1 T10756 ( .B(T15328_Y), .A(T15328_Y), .Y(T10756_Y));
KC_AND2_X1 T7985 ( .B(T15459_Y), .A(T1505_Y), .Y(T7985_Y));
KC_AND2_X1 T7925 ( .B(T15459_Y), .A(T1505_Y), .Y(T7925_Y));
KC_AND2_X1 T6716 ( .B(T12947_Y), .A(T1930_Y), .Y(T6716_Y));
KC_AND2_X1 T5836 ( .B(T15426_Y), .A(T1929_Y), .Y(T5836_Y));
KC_AND2_X1 T6212 ( .B(T11498_Y), .A(T15959_Y), .Y(T6212_Y));
KC_AND2_X1 T6342 ( .B(T2243_Y), .A(T3306_Y), .Y(T6342_Y));
KC_AND2_X1 T6563 ( .B(T12869_Y), .A(T290_Y), .Y(T6563_Y));
KC_AND2_X1 T5709 ( .B(T15346_Y), .A(T1929_Y), .Y(T5709_Y));
KC_AND2_X1 T5743 ( .B(T15380_Y), .A(T1929_Y), .Y(T5743_Y));
KC_AND2_X1 T5728 ( .B(T15380_Y), .A(T1929_Y), .Y(T5728_Y));
KC_AND2_X1 T5918 ( .B(T15508_Y), .A(T1505_Y), .Y(T5918_Y));
KC_AND2_X1 T5901 ( .B(T15508_Y), .A(T1505_Y), .Y(T5901_Y));
KC_AND2_X1 T5970 ( .B(T12769_Y), .A(T2651_Y), .Y(T5970_Y));
KC_AND2_X1 T6095 ( .B(T2706_Y), .A(T2705_Y), .Y(T6095_Y));
KC_AND2_X1 T6150 ( .B(T3283_Y), .A(T2744_Y), .Y(T6150_Y));
KC_AND2_X1 T6477 ( .B(T8401_Y), .A(T2871_Y), .Y(T6477_Y));
KC_AND2_X1 T5949 ( .B(T12760_Y), .A(T2651_Y), .Y(T5949_Y));
KC_AND2_X1 T5948 ( .B(T12743_Y), .A(T2651_Y), .Y(T5948_Y));
KC_AND2_X1 T6093 ( .B(T15561_Y), .A(T15184_Y), .Y(T6093_Y));
KC_AND2_X1 T6092 ( .B(T15561_Y), .A(T15184_Y), .Y(T6092_Y));
KC_AND2_X1 T6271 ( .B(T15707_Y), .A(T15187_Y), .Y(T6271_Y));
KC_AND2_X1 T6333 ( .B(T15599_Y), .A(T15187_Y), .Y(T6333_Y));
KC_AND2_X1 T6308 ( .B(T15599_Y), .A(T15187_Y), .Y(T6308_Y));
KC_AND2_X1 T6508 ( .B(T6551_Y), .A(T15187_Y), .Y(T6508_Y));
KC_AND2_X1 T6507 ( .B(T6551_Y), .A(T15187_Y), .Y(T6507_Y));
KC_AND2_X1 T5829 ( .B(T15423_Y), .A(T15184_Y), .Y(T5829_Y));
KC_AND2_X1 T5828 ( .B(T15423_Y), .A(T15184_Y), .Y(T5828_Y));
KC_AND2_X1 T5933 ( .B(T15510_Y), .A(T15184_Y), .Y(T5933_Y));
KC_AND2_X1 T6293 ( .B(T15707_Y), .A(T15187_Y), .Y(T6293_Y));
KC_AND2_X1 T6469 ( .B(T6137_Y), .A(T8502_Y), .Y(T6469_Y));
KC_AND2_X1 T5723 ( .B(T15362_Y), .A(T1929_Y), .Y(T5723_Y));
KC_AND2_X1 T5716 ( .B(T15362_Y), .A(T1929_Y), .Y(T5716_Y));
KC_AND2_X1 T5744 ( .B(T15678_Y), .A(T15184_Y), .Y(T5744_Y));
KC_AND2_X1 T6779 ( .B(T4564_Y), .A(T3940_Y), .Y(T6779_Y));
KC_AND2_X1 T6325 ( .B(T16020_Y), .A(T16020_Y), .Y(T6325_Y));
KC_AND2_X1 T15165 ( .B(T15330_Y), .A(T13211_Y), .Y(T15165_Y));
KC_AND2_X1 T10787 ( .B(T15416_Y), .A(T1505_Y), .Y(T10787_Y));
KC_AND2_X1 T6675 ( .B(T15426_Y), .A(T1929_Y), .Y(T6675_Y));
KC_AND2_X1 T6772 ( .B(T15162_Y), .A(T16000_Y), .Y(T6772_Y));
KC_AND2_X1 T6705 ( .B(T5737_Y), .A(T15184_Y), .Y(T6705_Y));
KC_AND2_X1 T6704 ( .B(T5737_Y), .A(T15184_Y), .Y(T6704_Y));
KC_AND2_X1 T6628 ( .B(T15678_Y), .A(T15184_Y), .Y(T6628_Y));
KC_AND2_X1 T5708 ( .B(T15346_Y), .A(T1929_Y), .Y(T5708_Y));
KC_AND2_X1 T7409 ( .B(T15410_Y), .A(T662_Y), .Y(T7409_Y));
KC_AND2_X1 T5931 ( .B(T15510_Y), .A(T15184_Y), .Y(T5931_Y));
KC_XNOR2_X8 T10031 ( .B(T15064_Y), .A(T8882_Y), .Y(T10031_Y));
KC_XNOR2_X8 T9490 ( .B(T15061_Y), .A(T8878_Y), .Y(T9490_Y));
KC_XNOR2_X8 T9489 ( .B(T9448_Y), .A(T9248_Y), .Y(T9489_Y));
KC_XNOR2_X8 T9488 ( .B(T9146_Y), .A(T9492_Y), .Y(T9488_Y));
KC_XNOR2_X8 T9143 ( .B(T9105_Y), .A(T9237_Y), .Y(T9143_Y));
KC_XNOR2_X8 T6800 ( .B(T9122_Y), .A(T9212_Y), .Y(T6800_Y));
KC_XNOR2_X8 T9116 ( .B(T9070_Y), .A(T9210_Y), .Y(T9116_Y));
KC_XNOR2_X8 T9101 ( .B(T9147_Y), .A(T9493_Y), .Y(T9101_Y));
KC_XNOR2_X8 T9058 ( .B(T9104_Y), .A(T9206_Y), .Y(T9058_Y));
KC_XNOR2_X8 T9016 ( .B(T9108_Y), .A(T9250_Y), .Y(T9016_Y));
KC_XNOR2_X8 T8871 ( .B(T9064_Y), .A(T9198_Y), .Y(T8871_Y));
KC_XNOR2_X8 T8397 ( .B(T9063_Y), .A(T9197_Y), .Y(T8397_Y));
KC_XNOR2_X8 T5587 ( .B(T8128_Y), .A(T4842_Y), .Y(T5587_Y));
KC_XNOR2_X8 T5147 ( .B(T1270_Q), .A(T4902_Y), .Y(T5147_Y));
KC_XNOR2_X8 T2103 ( .B(T5404_Q), .A(T4868_Y), .Y(T2103_Y));
KC_XNOR2_X8 T4951 ( .B(T13053_Q), .A(T4865_Y), .Y(T4951_Y));
KC_XNOR2_X8 T4702 ( .B(T7702_Y), .A(T1665_Q), .Y(T4702_Y));
KC_XNOR2_X8 T4419 ( .B(T1578_Y), .A(T1597_Y), .Y(T4419_Y));
KC_XNOR2_X8 T4412 ( .B(T1058_Y), .A(T1450_Y), .Y(T4412_Y));
KC_XNOR2_X8 T3898 ( .B(T1517_Y), .A(T16413_Q), .Y(T3898_Y));
KC_XNOR2_X8 T3786 ( .B(T15519_Y), .A(T8880_Q), .Y(T3786_Y));
KC_XNOR2_X8 T3785 ( .B(T5486_Q), .A(T4912_Y), .Y(T3785_Y));
KC_XNOR2_X8 T3784 ( .B(T5494_Q), .A(T2259_Y), .Y(T3784_Y));
KC_XNOR2_X8 T3079 ( .B(T2313_Q), .A(T2310_Y), .Y(T3079_Y));
KC_XNOR2_X8 T2687 ( .B(T2345_Q), .A(T2261_Y), .Y(T2687_Y));
KC_XNOR2_X8 T2574 ( .B(T2316_Q), .A(T2298_Y), .Y(T2574_Y));
KC_XNOR2_X8 T2398 ( .B(T2315_Q), .A(T2293_Y), .Y(T2398_Y));
KC_XNOR2_X8 T4157 ( .B(T4767_Y), .A(T5501_Q), .Y(T4157_Y));
KC_XNOR2_X8 T412 ( .B(T4777_Y), .A(T4663_Q), .Y(T412_Y));
KC_XNOR2_X8 T408 ( .B(T4769_Y), .A(T4685_Q), .Y(T408_Y));
KC_XNOR2_X8 T394 ( .B(T4772_Y), .A(T4675_Q), .Y(T394_Y));
KC_XNOR2_X8 T392 ( .B(T4766_Y), .A(T5513_Q), .Y(T392_Y));
KC_XNOR2_X8 T267 ( .B(T4774_Y), .A(T4043_Q), .Y(T267_Y));
KC_XNOR2_X8 T263 ( .B(T4776_Y), .A(T4714_Q), .Y(T263_Y));
KC_XNOR2_X8 T2642 ( .B(T4771_Y), .A(T5496_Q), .Y(T2642_Y));
KC_XNOR2_X8 T262 ( .B(T4765_Y), .A(T4056_Q), .Y(T262_Y));
KC_XNOR2_X8 T261 ( .B(T4763_Y), .A(T16049_Q), .Y(T261_Y));
KC_XNOR2_X8 T259 ( .B(T4762_Y), .A(T5502_Q), .Y(T259_Y));
KC_XNOR2_X8 T258 ( .B(T4770_Y), .A(T4693_Q), .Y(T258_Y));
KC_XNOR2_X8 T241 ( .B(T4768_Y), .A(T4686_Q), .Y(T241_Y));
KC_XNOR2_X8 T240 ( .B(T9106_Y), .A(T9499_Y), .Y(T240_Y));
KC_XNOR2_X8 T233 ( .B(T9103_Y), .A(T9213_Y), .Y(T233_Y));
KC_XNOR2_X8 T231 ( .B(T9165_Y), .A(T9183_Y), .Y(T231_Y));
KC_AOI31_X1 T9059 ( .B2(T10941_Y), .B0(T16274_Y), .Y(T9059_Y),     .A(T4895_Y), .B1(T10188_Y));
KC_NOR3_X4 T16182 ( .Y(T16182_Y), .B(T4921_Y), .C(T2539_Y),     .A(T1675_Q));
KC_NOR3_X4 T16236 ( .Y(T16236_Y), .B(T12110_Y), .C(T2067_Y),     .A(T2643_Y));
KC_OAI22_X3 T16170 ( .A1(T1352_Y), .B0(T5307_Y), .B1(T9166_Y),     .A0(T5335_Y), .Y(T16170_Y));
KC_NOR2_X4 T16006 ( .Y(T16006_Y), .A(T2839_Y), .B(T6070_Y));
KC_NOR2_X4 T16149 ( .Y(T16149_Y), .A(T6190_Y), .B(T10977_Y));
KC_NOR2_X4 T8503 ( .Y(T8503_Y), .A(T2838_Y), .B(T12322_Y));
KC_NOR2_X4 T10257 ( .Y(T10257_Y), .A(T4872_Y), .B(T2633_Y));
KC_NOR2_X4 T16168 ( .Y(T16168_Y), .A(T2076_Y), .B(T2074_Y));
KC_BUF_X13 T536 ( .Y(T536_Y), .A(T685_Y));
KC_BUF_X13 T226 ( .Y(T226_Y), .A(T685_Y));
KC_BUF_X13 T398 ( .Y(T398_Y), .A(T685_Y));
KC_BUF_X13 T16392 ( .Y(T16392_Y), .A(T1600_Y));
KC_BUF_X13 T5351 ( .Y(T5351_Y), .A(T15182_Q));
KC_BUF_X13 T5725 ( .Y(T5725_Y), .A(T15188_Y));
KC_BUF_X13 T4897 ( .Y(T4897_Y), .A(T14964_Y));
KC_BUF_X13 T16134 ( .Y(T16134_Y), .A(T2097_Y));
KC_BUF_X13 T16253 ( .Y(T16253_Y), .A(T4897_Y));
KC_BUF_X13 T943 ( .Y(T943_Y), .A(T14982_Y));
KC_BUF_X13 T5715 ( .Y(T5715_Y), .A(T4897_Y));
KC_TLAT_X2 T15179 ( .D(T12446_Y), .Q(T15179_Q), .CK(T5423_Y));
KC_TLAT_X2 T15189 ( .D(T1289_Y), .Q(T15189_Q), .CK(T15168_Q));
KC_TLAT_X2 T15183 ( .D(T6334_Y), .Q(T15183_Q), .CK(T1380_Y));
KC_TLAT_X2 T15182 ( .D(T16148_Y), .Q(T15182_Q), .CK(T1376_Y));
KC_TLAT_X2 T15181 ( .D(T1288_Y), .Q(T15181_Q), .CK(T13064_Q));
KC_TLAT_X2 T15177 ( .D(T1379_Y), .Q(T15177_Q), .CK(T13064_Q));
KC_TLAT_X2 T15191 ( .D(T15006_Y), .Q(T15191_Q), .CK(T1382_Y));
KC_TLAT_X2 T15178 ( .D(T1379_Y), .Q(T15178_Q), .CK(T1384_Y));
KC_TLAT_X2 T15168 ( .D(T15543_Y), .Q(T15168_Q), .CK(T15168_CK));
KC_BUF_X1 T130 ( .Y(T130_Y), .A(T13440_Q));
KC_BUF_X1 T662 ( .Y(T662_Y), .A(T15180_Y));
KC_BUF_X1 T774 ( .Y(T774_Y), .A(T991_Y));
KC_BUF_X1 T942 ( .Y(T942_Y), .A(T991_Y));
KC_BUF_X1 T959 ( .Y(T959_Y), .A(T14369_Q));
KC_BUF_X1 T1011 ( .Y(T1011_Y), .A(T14369_Q));
KC_BUF_X1 T1105 ( .Y(T1105_Y), .A(T991_Y));
KC_BUF_X1 T1137 ( .Y(T1137_Y), .A(T943_Y));
KC_BUF_X1 T1324 ( .Y(T1324_Y), .A(T1403_Y));
KC_BUF_X1 T1505 ( .Y(T1505_Y), .A(T15180_Y));
KC_BUF_X1 T1855 ( .Y(T1855_Y), .A(T1855_A));
KC_BUF_X1 T1929 ( .Y(T1929_Y), .A(T15180_Y));
KC_BUF_X1 T2157 ( .Y(T2157_Y), .A(T2156_Y));
KC_BUF_X1 T3217 ( .Y(T3217_Y), .A(T3215_Y));
KC_BUF_X1 T3888 ( .Y(T3888_Y), .A(T869_Y));
KC_BUF_X1 T4841 ( .Y(T4841_Y), .A(T13262_Y));
KC_BUF_X1 T4879 ( .Y(T4879_Y), .A(T15179_Q));
KC_BUF_X1 T5423 ( .Y(T5423_Y), .A(T15188_Y));
KC_OR3_X1 T14971 ( .Y(T14971_Y), .A(T107_Q), .B(T5604_Y), .C(T5605_Y));
KC_OR3_X1 T14981 ( .Y(T14981_Y), .A(T683_Q), .B(T698_Q), .C(T689_Q));
KC_OR3_X1 T15036 ( .Y(T15036_Y), .A(T1764_Y), .B(T1765_Y),     .C(T11531_Y));
KC_OR3_X1 T14966 ( .Y(T14966_Y), .A(T2072_Y), .B(T10253_Y),     .C(T2074_Y));
KC_OR3_X1 T15019 ( .Y(T15019_Y), .A(T13132_Q), .B(T2723_Y),     .C(T2152_Q));
KC_OR3_X1 T14969 ( .Y(T14969_Y), .A(T2341_Y), .B(T4962_Y),     .C(T6540_Y));
KC_OR3_X1 T15007 ( .Y(T15007_Y), .A(T3807_Y), .B(T3799_Y),     .C(T5433_Y));
KC_OR3_X1 T15012 ( .Y(T15012_Y), .A(T14494_Q), .B(T4486_Y),     .C(T3856_Y));
KC_OR3_X1 T15025 ( .Y(T15025_Y), .A(T154_Q), .B(T157_Q), .C(T151_Q));
KC_OR3_X1 T15010 ( .Y(T15010_Y), .A(T14540_Q), .B(T14543_Q),     .C(T14541_Q));
KC_NAND4B_X1 T12371 ( .C(T8545_Y), .B(T5203_Q), .A(T107_Q),     .Y(T12371_Y), .DN(T5596_Y));
KC_NAND4B_X1 T12369 ( .C(T15316_Y), .B(T8555_Y), .A(T5203_Q),     .Y(T12369_Y), .DN(T5619_Y));
KC_NAND4B_X1 T12383 ( .C(T8578_Y), .B(T136_Q), .A(T5225_Q),     .Y(T12383_Y), .DN(T8581_Y));
KC_NAND4B_X1 T12382 ( .C(T260_Y), .B(T5225_Q), .A(T131_Q),     .Y(T12382_Y), .DN(T6934_Y));
KC_NAND4B_X1 T12418 ( .C(T647_Y), .B(T212_Q), .A(T208_Q), .Y(T12418_Y),     .DN(T223_Q));
KC_NAND4B_X1 T12443 ( .C(T9397_Y), .B(T941_Y), .A(T878_Y),     .Y(T12443_Y), .DN(T9270_Y));
KC_NAND4B_X1 T12451 ( .C(T7862_Y), .B(T8873_Y), .A(T7917_Y),     .Y(T12451_Y), .DN(T7913_Y));
KC_NAND4B_X1 T4917 ( .C(T5228_Y), .B(T957_Y), .A(T9115_Y), .Y(T4917_Y),     .DN(T9174_Y));
KC_NAND4B_X1 T1327 ( .C(T1350_Y), .B(T8981_Y), .A(T572_Q), .Y(T1327_Y),     .DN(T8073_Y));
KC_NAND4B_X1 T12400 ( .C(T11171_Y), .B(T11193_Y), .A(T514_Y),     .Y(T12400_Y), .DN(T9723_Y));
KC_NAND4B_X1 T12087 ( .C(T15500_Y), .B(T927_Y), .A(T1133_Q),     .Y(T12087_Y), .DN(T980_Q));
KC_NAND4B_X1 T12093 ( .C(T9982_Y), .B(T1365_Y), .A(T1366_Y),     .Y(T12093_Y), .DN(T10159_Y));
KC_NAND4B_X1 T12110 ( .C(T12982_Y), .B(T10936_Y), .A(T1366_Y),     .Y(T12110_Y), .DN(T16040_Y));
KC_NAND4B_X1 T12111 ( .C(T16233_Y), .B(T4902_Y), .A(T10154_Y),     .Y(T12111_Y), .DN(T3966_Y));
KC_NAND4B_X1 T12160 ( .C(T6097_Co), .B(T2098_Y), .A(T6097_Co),     .Y(T12160_Y), .DN(T6097_S));
KC_NAND4B_X1 T12314 ( .C(T12869_Y), .B(T2346_Y), .A(T2317_Y),     .Y(T12314_Y), .DN(T2317_Y));
KC_NAND4B_X1 T12085 ( .C(T5318_Y), .B(T2507_Y), .A(T15447_Y),     .Y(T12085_Y), .DN(T2507_Y));
KC_NAND4B_X1 T12091 ( .C(T10517_Y), .B(T2583_Q), .A(T2570_Q),     .Y(T12091_Y), .DN(T2584_Q));
KC_NAND4B_X1 T12115 ( .C(T2666_Y), .B(T2654_Y), .A(T10276_Y),     .Y(T12115_Y), .DN(T2674_Y));
KC_NAND4B_X1 T12336 ( .C(T12789_Y), .B(T2686_Y), .A(T2678_Y),     .Y(T12336_Y), .DN(T4993_Y));
KC_NAND4B_X1 T12164 ( .C(T2702_Y), .B(T15851_Y), .A(T1743_Y),     .Y(T12164_Y), .DN(T10887_Y));
KC_NAND4B_X1 T12253 ( .C(T8351_Y), .B(T6324_Y), .A(T2263_Y),     .Y(T12253_Y), .DN(T10964_Y));
KC_NAND4B_X1 T12276 ( .C(T2862_Y), .B(T6208_Y), .A(T12275_Y),     .Y(T12276_Y), .DN(T10624_Y));
KC_NAND4B_X1 T12297 ( .C(T290_Y), .B(T8426_Y), .A(T2948_Y),     .Y(T12297_Y), .DN(T2936_Y));
KC_NAND4B_X1 T12066 ( .C(T11005_Y), .B(T6506_Y), .A(T5536_Q),     .Y(T12066_Y), .DN(T10570_Y));
KC_NAND4B_X1 T12132 ( .C(T3207_Y), .B(T3815_Y), .A(T12955_Y),     .Y(T12132_Y), .DN(T11987_Y));
KC_NAND4B_X1 T12210 ( .C(T6230_S), .B(T3315_Y), .A(T3293_Y),     .Y(T12210_Y), .DN(T3296_Y));
KC_NAND4B_X1 T12284 ( .C(T12285_Y), .B(T6144_Y), .A(T6144_Y),     .Y(T12284_Y), .DN(T8401_Y));
KC_NAND4B_X1 T12322 ( .C(T6514_Y), .B(T6489_Y), .A(T3522_Q),     .Y(T12322_Y), .DN(T11006_Y));
KC_NAND4B_X1 T12134 ( .C(T10889_Y), .B(T3790_Y), .A(T15836_Y),     .Y(T12134_Y), .DN(T11330_Y));
KC_NAND4B_X1 T12167 ( .C(T14546_Q), .B(T14544_Q), .A(T14540_Q),     .Y(T12167_Y), .DN(T3223_Y));
KC_NAND4B_X1 T12159 ( .C(T3843_Y), .B(T11980_Y), .A(T4385_Y),     .Y(T12159_Y), .DN(T11372_Y));
KC_NAND4B_X1 T12186 ( .C(T3265_Y), .B(T15939_Y), .A(T3868_Y),     .Y(T12186_Y), .DN(T6797_S));
KC_NAND4B_X1 T12182 ( .C(T12806_Y), .B(T15910_Y), .A(T5858_Y),     .Y(T12182_Y), .DN(T5130_Q));
KC_NAND4B_X1 T12195 ( .C(T15963_Y), .B(T4541_Y), .A(T4541_Y),     .Y(T12195_Y), .DN(T4541_Y));
KC_NAND4B_X1 T12348 ( .C(T10944_Y), .B(T12013_Y), .A(T5554_Y),     .Y(T12348_Y), .DN(T8271_Y));
KC_NAND4B_X1 T12243 ( .C(T3975_Y), .B(T6020_Y), .A(T15704_Y),     .Y(T12243_Y), .DN(T4588_Y));
KC_NAND4B_X1 T12281 ( .C(T4716_Y), .B(T4691_Y), .A(T12277_Y),     .Y(T12281_Y), .DN(T6151_Y));
KC_NAND4B_X1 T12071 ( .C(T4168_Q), .B(T11764_Y), .A(T11736_Y),     .Y(T12071_Y), .DN(T4119_Y));
KC_NAND4B_X1 T12150 ( .C(T5854_Y), .B(T5853_Y), .A(T4486_Y),     .Y(T12150_Y), .DN(T4441_Y));
KC_NAND4B_X1 T12356 ( .C(T4481_Y), .B(T12355_Y), .A(T11451_Y),     .Y(T12356_Y), .DN(T12208_Y));
KC_NAND4B_X1 T12355 ( .C(T5932_Y), .B(T11454_Y), .A(T4497_Y),     .Y(T12355_Y), .DN(T4506_Y));
KC_NAND4B_X1 T12181 ( .C(T15697_Y), .B(T14551_Q), .A(T14547_Q),     .Y(T12181_Y), .DN(T4478_Y));
KC_NAND4B_X1 T12199 ( .C(T15969_Y), .B(T5888_Y), .A(T8247_Y),     .Y(T12199_Y), .DN(T15971_Y));
KC_NAND4B_X1 T12196 ( .C(T4532_Y), .B(T15968_Y), .A(T4475_Y),     .Y(T12196_Y), .DN(T5879_Y));
KC_NAND4B_X1 T12212 ( .C(T12016_Y), .B(T4575_Q), .A(T4572_Q),     .Y(T12212_Y), .DN(T4556_Y));
KC_NAND4B_X1 T12238 ( .C(T6023_Y), .B(T6009_Y), .A(T6009_Y),     .Y(T12238_Y), .DN(T6009_Y));
KC_NAND4B_X1 T12277 ( .C(T6151_Y), .B(T4698_Y), .A(T4698_Y),     .Y(T12277_Y), .DN(T4716_Y));
KC_NAND4B_X1 T12308 ( .C(T4735_Y), .B(T4738_Y), .A(T11787_Y),     .Y(T12308_Y), .DN(T4732_Y));
KC_NAND4B_X1 T12449 ( .C(T927_Y), .B(T946_Y), .A(T1133_Q),     .Y(T12449_Y), .DN(T980_Q));
KC_NAND4B_X1 T4916 ( .C(T13258_Y), .B(T5224_Y), .A(T16077_Y),     .Y(T4916_Y), .DN(T10138_Y));
KC_NAND4B_X1 T12174 ( .C(T3230_Y), .B(T6068_Y), .A(T3830_Y),     .Y(T12174_Y), .DN(T5843_Y));
KC_AO222_X1 T12313 ( .A0(T10998_Y), .Y(T12313_Y), .C1(T2331_Y),     .C0(T2350_Y), .B1(T6243_Y), .B0(T6243_Y), .A1(T2323_Y));
KC_AO222_X1 T12118 ( .A0(T10241_Y), .Y(T12118_Y), .C1(T10242_Y),     .C0(T2461_Y), .B1(T2512_Y), .B0(T10270_Y), .A1(T14480_Q));
KC_AO222_X1 T12117 ( .A0(T10241_Y), .Y(T12117_Y), .C1(T10242_Y),     .C0(T2485_Y), .B1(T2513_Y), .B0(T10270_Y), .A1(T14479_Q));
KC_AO222_X1 T12179 ( .A0(T15844_Q), .Y(T12179_Y), .C1(T5791_Y),     .C0(T16098_Y), .B1(T3245_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12178 ( .A0(T5076_Q), .Y(T12178_Y), .C1(T2671_Y),     .C0(T5791_Y), .B1(T5845_Y), .B0(T15005_Y), .A1(T3872_Y));
KC_AO222_X1 T12177 ( .A0(T15796_Q), .Y(T12177_Y), .C1(T5791_Y),     .C0(T16071_Y), .B1(T3226_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12176 ( .A0(T5439_Q), .Y(T12176_Y), .C1(T2670_Y),     .C0(T5791_Y), .B1(T5845_Y), .B0(T16088_Q), .A1(T3872_Y));
KC_AO222_X1 T12175 ( .A0(T15798_Q), .Y(T12175_Y), .C1(T5791_Y),     .C0(T16096_Y), .B1(T2710_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12171 ( .A0(T15809_Q), .Y(T12171_Y), .C1(T5791_Y),     .C0(T16097_Y), .B1(T2716_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12170 ( .A0(T2711_Q), .Y(T12170_Y), .C1(T16235_Y),     .C0(T5791_Y), .B1(T5845_Y), .B0(T15807_Q), .A1(T3872_Y));
KC_AO222_X1 T12169 ( .A0(T15805_Q), .Y(T12169_Y), .C1(T5791_Y),     .C0(T16073_Y), .B1(T5441_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12163 ( .A0(T2703_Y), .Y(T12163_Y), .C1(T15886_Y),     .C0(T2712_Y), .B1(T5819_Y), .B0(T2124_Y), .A1(T5819_Y));
KC_AO222_X1 T12162 ( .A0(T16299_Q), .Y(T12162_Y), .C1(T5791_Y),     .C0(T16074_Y), .B1(T2713_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12161 ( .A0(T15808_Q), .Y(T12161_Y), .C1(T5791_Y),     .C0(T16072_Y), .B1(T2715_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12154 ( .A0(T3228_Q), .Y(T12154_Y), .C1(T16075_Y),     .C0(T5791_Y), .B1(T5845_Y), .B0(T15803_Q), .A1(T3872_Y));
KC_AO222_X1 T12153 ( .A0(T5380_Q), .Y(T12153_Y), .C1(T5791_Y),     .C0(T16069_Y), .B1(T3244_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12068 ( .A0(T15044_Y), .Y(T12068_Y), .C1(T6538_Y),     .C0(T2948_Y), .B1(T6580_Y), .B0(T6561_Y), .A1(T6196_Y));
KC_AO222_X1 T12343 ( .A0(T5041_Y), .Y(T12343_Y), .C1(T5040_Y),     .C0(T11015_Y), .B1(T15562_Y), .B0(T3210_Y), .A1(T11989_Y));
KC_AO222_X1 T12215 ( .A0(T3324_Y), .Y(T12215_Y), .C1(T12463_Y),     .C0(T3333_Y), .B1(T3344_Y), .B0(T3333_Y), .A1(T3332_Y));
KC_AO222_X1 T12244 ( .A0(T10618_Y), .Y(T12244_Y), .C1(T4097_Y),     .C0(T8392_Y), .B1(T6484_Y), .B0(T12281_Y), .A1(T4072_Y));
KC_AO222_X1 T12282 ( .A0(T8401_Y), .Y(T12282_Y), .C1(T6478_Y),     .C0(T6477_Y), .B1(T8393_Y), .B0(T5509_Y), .A1(T16502_Y));
KC_AO222_X1 T12184 ( .A0(T5140_Y), .Y(T12184_Y), .C1(T6167_S),     .C0(T5868_Y), .B1(T3903_Y), .B0(T10634_Y), .A1(T3871_Y));
KC_AO222_X1 T12235 ( .A0(T4042_Y), .Y(T12235_Y), .C1(T4042_Y),     .C0(T12957_Y), .B1(T6033_Y), .B0(T4011_Y), .A1(T15610_Y));
KC_AO222_X1 T12346 ( .A0(T4037_Y), .Y(T12346_Y), .C1(T16017_Y),     .C0(T3984_Y), .B1(T16030_Y), .B0(T4928_Y), .A1(T12246_Y));
KC_AO222_X1 T12292 ( .A0(T11735_Y), .Y(T12292_Y), .C1(T11781_Y),     .C0(T5530_Q), .B1(T4138_Y), .B0(T6547_Y), .A1(T10581_Y));
KC_AO222_X1 T12318 ( .A0(T5115_Y), .Y(T12318_Y), .C1(T4761_Y),     .C0(T4158_Y), .B1(T8166_Y), .B0(T5115_Y), .A1(T4175_Y));
KC_AO222_X1 T12242 ( .A0(T4593_Y), .Y(T12242_Y), .C1(T3308_Y),     .C0(T12834_Y), .B1(T4593_Y), .B0(T12834_Y), .A1(T8331_Y));
KC_AO222_X1 T12339 ( .A0(T3246_Q), .Y(T12339_Y), .C1(T2673_Y),     .C0(T5791_Y), .B1(T5845_Y), .B0(T15797_Q), .A1(T3872_Y));
KC_AO222_X1 T12338 ( .A0(T964_Q), .Y(T12338_Y), .C1(T5791_Y),     .C0(T16076_Y), .B1(T5075_Q), .B0(T3872_Y), .A1(T5845_Y));
KC_AO222_X1 T12119 ( .A0(T10241_Y), .Y(T12119_Y), .C1(T10242_Y),     .C0(T2455_Y), .B1(T2509_Y), .B0(T10270_Y), .A1(T14465_Q));
KC_AO222_X1 T12152 ( .A0(T3227_Q), .Y(T12152_Y), .C1(T16070_Y),     .C0(T5791_Y), .B1(T5845_Y), .B0(T16301_Q), .A1(T3872_Y));
KC_OR2_X4 T10202 ( .Y(T10202_Y), .A(T5937_Y), .B(T3904_Y));
KC_OR2_X4 T10201 ( .Y(T10201_Y), .A(T2750_Y), .B(T3283_Y));
KC_DFFSNHQ_X2 T13054 ( .Q(T13054_Q), .D(T1298_Y), .CK(T14998_Y),     .SN(T13053_SN));
KC_DFFSNHQ_X2 T16488 ( .Q(T16488_Q), .D(T2090_Y), .CK(T14554_Q),     .SN(T15034_Y));
KC_DFFSNHQ_X2 T16487 ( .Q(T16487_Q), .D(T2094_Y), .CK(T14554_Q),     .SN(T15008_Y));
KC_DFFSNHQ_X2 T16486 ( .Q(T16486_Q), .D(T2092_Y), .CK(T14554_Q),     .SN(T15008_Y));
KC_DFFSNHQ_X2 T16485 ( .Q(T16485_Q), .D(T2094_Y), .CK(T14960_Q),     .SN(T15008_Y));
KC_DFFSNHQ_X2 T16484 ( .Q(T16484_Q), .D(T2092_Y), .CK(T14960_Q),     .SN(T15008_Y));
KC_DFFSNHQ_X2 T16483 ( .Q(T16483_Q), .D(T2088_Y), .CK(T14554_Q),     .SN(T15008_Y));
KC_DFFSNHQ_X2 T1984 ( .Q(T1984_Q), .D(T15040_Y), .CK(T14960_Q),     .SN(T15008_Y));
KC_DFFSNHQ_X2 T16481 ( .Q(T16481_Q), .D(T13098_Y), .CK(T14960_Q),     .SN(T15015_Y));
KC_DFFSNHQ_X2 T4924 ( .Q(T4924_Q), .D(T15124_Y), .CK(T14554_Q),     .SN(T15011_Y));
KC_DFFSNHQ_X2 T13102 ( .Q(T13102_Q), .D(T2158_Y), .CK(T14554_Q),     .SN(T15011_Y));
KC_TIELO_X1 T15330 ( .Y(T15330_Y));
KC_TIELO_X1 T15329 ( .Y(T15329_Y));
KC_TIELO_X1 T13074 ( .Y(T13074_Y));
KC_TIELO_X1 T15326 ( .Y(T15326_Y));
KC_TIELO_X1 T15325 ( .Y(T15325_Y));
KC_TIELO_X1 T13317 ( .Y(T13317_Y));
KC_TIELO_X1 T13080 ( .Y(T13080_Y));
KC_TIELO_X1 T15323 ( .Y(T15323_Y));
KC_TIELO_X1 T15322 ( .Y(T15322_Y));
KC_TIELO_X1 T15170 ( .Y(T15170_Y));
KC_TIELO_X1 T16490 ( .Y(T16490_Y));
KC_TIELO_X1 T15337 ( .Y(T15337_Y));
KC_TIELO_X1 T6832 ( .Y(T6832_Y));
KC_TIELO_X1 T570 ( .Y(T570_Y));
KC_TIELO_X1 T15653 ( .Y(T15653_Y));
KC_TIELO_X1 T15652 ( .Y(T15652_Y));
KC_TIELO_X1 T643 ( .Y(T643_Y));
KC_TIELO_X1 T15370 ( .Y(T15370_Y));
KC_TIELO_X1 T15368 ( .Y(T15368_Y));
KC_TIELO_X1 T15657 ( .Y(T15657_Y));
KC_TIELO_X1 T15483 ( .Y(T15483_Y));
KC_TIELO_X1 T15541 ( .Y(T15541_Y));
KC_TIELO_X1 T785 ( .Y(T785_Y));
KC_TIELO_X1 T16175 ( .Y(T16175_Y));
KC_TIELO_X1 T15456 ( .Y(T15456_Y));
KC_TIELO_X1 T15482 ( .Y(T15482_Y));
KC_TIELO_X1 T15539 ( .Y(T15539_Y));
KC_TIELO_X1 T15649 ( .Y(T15649_Y));
KC_TIELO_X1 T15334 ( .Y(T15334_Y));
KC_TIELO_X1 T15333 ( .Y(T15333_Y));
KC_TIELO_X1 T15409 ( .Y(T15409_Y));
KC_TIELO_X1 T885 ( .Y(T885_Y));
KC_TIELO_X1 T16300 ( .Y(T16300_Y));
KC_TIELO_X1 T15481 ( .Y(T15481_Y));
KC_TIELO_X1 T15522 ( .Y(T15522_Y));
KC_TIELO_X1 T15672 ( .Y(T15672_Y));
KC_TIELO_X1 T15410 ( .Y(T15410_Y));
KC_TIELO_X1 T15465 ( .Y(T15465_Y));
KC_TIELO_X1 T15491 ( .Y(T15491_Y));
KC_TIELO_X1 T15521 ( .Y(T15521_Y));
KC_TIELO_X1 T15460 ( .Y(T15460_Y));
KC_TIELO_X1 T15499 ( .Y(T15499_Y));
KC_TIELO_X1 T15498 ( .Y(T15498_Y));
KC_TIELO_X1 T15528 ( .Y(T15528_Y));
KC_TIELO_X1 T15544 ( .Y(T15544_Y));
KC_TIELO_X1 T15343 ( .Y(T15343_Y));
KC_TIELO_X1 T15340 ( .Y(T15340_Y));
KC_TIELO_X1 T15394 ( .Y(T15394_Y));
KC_TIELO_X1 T588 ( .Y(T588_Y));
KC_TIELO_X1 T15418 ( .Y(T15418_Y));
KC_TIELO_X1 T15417 ( .Y(T15417_Y));
KC_TIELO_X1 T15530 ( .Y(T15530_Y));
KC_TIELO_X1 T15345 ( .Y(T15345_Y));
KC_TIELO_X1 T15344 ( .Y(T15344_Y));
KC_TIELO_X1 T15341 ( .Y(T15341_Y));
KC_TIELO_X1 T15339 ( .Y(T15339_Y));
KC_TIELO_X1 T15338 ( .Y(T15338_Y));
KC_TIELO_X1 T15361 ( .Y(T15361_Y));
KC_TIELO_X1 T15360 ( .Y(T15360_Y));
KC_TIELO_X1 T15416 ( .Y(T15416_Y));
KC_TIELO_X1 T15414 ( .Y(T15414_Y));
KC_TIELO_X1 T15438 ( .Y(T15438_Y));
KC_TIELO_X1 T15661 ( .Y(T15661_Y));
KC_TIELO_X1 T15495 ( .Y(T15495_Y));
KC_TIELO_X1 T15494 ( .Y(T15494_Y));
KC_TIELO_X1 T15493 ( .Y(T15493_Y));
KC_TIELO_X1 T15526 ( .Y(T15526_Y));
KC_TIELO_X1 T15542 ( .Y(T15542_Y));
KC_TIELO_X1 T15668 ( .Y(T15668_Y));
KC_TIELO_X1 T15669 ( .Y(T15669_Y));
KC_TIELO_X1 T15359 ( .Y(T15359_Y));
KC_TIELO_X1 T15376 ( .Y(T15376_Y));
KC_TIELO_X1 T15374 ( .Y(T15374_Y));
KC_TIELO_X1 T16180 ( .Y(T16180_Y));
KC_TIELO_X1 T849 ( .Y(T849_Y));
KC_TIELO_X1 T818 ( .Y(T818_Y));
KC_TIELO_X1 T15437 ( .Y(T15437_Y));
KC_TIELO_X1 T1051 ( .Y(T1051_Y));
KC_TIELO_X1 T15459 ( .Y(T15459_Y));
KC_TIELO_X1 T15698 ( .Y(T15698_Y));
KC_TIELO_X1 T15718 ( .Y(T15718_Y));
KC_TIELO_X1 T15717 ( .Y(T15717_Y));
KC_TIELO_X1 T15716 ( .Y(T15716_Y));
KC_TIELO_X1 T15348 ( .Y(T15348_Y));
KC_TIELO_X1 T15427 ( .Y(T15427_Y));
KC_TIELO_X1 T15426 ( .Y(T15426_Y));
KC_TIELO_X1 T15479 ( .Y(T15479_Y));
KC_TIELO_X1 T15575 ( .Y(T15575_Y));
KC_TIELO_X1 T15950 ( .Y(T15950_Y));
KC_TIELO_X1 T15583 ( .Y(T15583_Y));
KC_TIELO_X1 T15617 ( .Y(T15617_Y));
KC_TIELO_X1 T6554 ( .Y(T6554_Y));
KC_TIELO_X1 T15346 ( .Y(T15346_Y));
KC_TIELO_X1 T373 ( .Y(T373_Y));
KC_TIELO_X1 T15380 ( .Y(T15380_Y));
KC_TIELO_X1 T1139 ( .Y(T1139_Y));
KC_TIELO_X1 T15475 ( .Y(T15475_Y));
KC_TIELO_X1 T15508 ( .Y(T15508_Y));
KC_TIELO_X1 T15505 ( .Y(T15505_Y));
KC_TIELO_X1 T15504 ( .Y(T15504_Y));
KC_TIELO_X1 T15547 ( .Y(T15547_Y));
KC_TIELO_X1 T15603 ( .Y(T15603_Y));
KC_TIELO_X1 T15710 ( .Y(T15710_Y));
KC_TIELO_X1 T15614 ( .Y(T15614_Y));
KC_TIELO_X1 T15715 ( .Y(T15715_Y));
KC_TIELO_X1 T15644 ( .Y(T15644_Y));
KC_TIELO_X1 T6838 ( .Y(T6838_Y));
KC_TIELO_X1 T15449 ( .Y(T15449_Y));
KC_TIELO_X1 T15446 ( .Y(T15446_Y));
KC_TIELO_X1 T15536 ( .Y(T15536_Y));
KC_TIELO_X1 T5737 ( .Y(T5737_Y));
KC_TIELO_X1 T5757 ( .Y(T5757_Y));
KC_TIELO_X1 T15695 ( .Y(T15695_Y));
KC_TIELO_X1 T15556 ( .Y(T15556_Y));
KC_TIELO_X1 T15564 ( .Y(T15564_Y));
KC_TIELO_X1 T15561 ( .Y(T15561_Y));
KC_TIELO_X1 T15560 ( .Y(T15560_Y));
KC_TIELO_X1 T15567 ( .Y(T15567_Y));
KC_TIELO_X1 T15595 ( .Y(T15595_Y));
KC_TIELO_X1 T15602 ( .Y(T15602_Y));
KC_TIELO_X1 T15599 ( .Y(T15599_Y));
KC_TIELO_X1 T6551 ( .Y(T6551_Y));
KC_TIELO_X1 T15626 ( .Y(T15626_Y));
KC_TIELO_X1 T15719 ( .Y(T15719_Y));
KC_TIELO_X1 T15642 ( .Y(T15642_Y));
KC_TIELO_X1 T15423 ( .Y(T15423_Y));
KC_TIELO_X1 T16109 ( .Y(T16109_Y));
KC_TIELO_X1 T15476 ( .Y(T15476_Y));
KC_TIELO_X1 T15517 ( .Y(T15517_Y));
KC_TIELO_X1 T15516 ( .Y(T15516_Y));
KC_TIELO_X1 T15514 ( .Y(T15514_Y));
KC_TIELO_X1 T15510 ( .Y(T15510_Y));
KC_TIELO_X1 T15563 ( .Y(T15563_Y));
KC_TIELO_X1 T15948 ( .Y(T15948_Y));
KC_TIELO_X1 T15979 ( .Y(T15979_Y));
KC_TIELO_X1 T15680 ( .Y(T15680_Y));
KC_TIELO_X1 T15364 ( .Y(T15364_Y));
KC_TIELO_X1 T15363 ( .Y(T15363_Y));
KC_TIELO_X1 T15362 ( .Y(T15362_Y));
KC_TIELO_X1 T15386 ( .Y(T15386_Y));
KC_TIELO_X1 T15385 ( .Y(T15385_Y));
KC_TIELO_X1 T15382 ( .Y(T15382_Y));
KC_TIELO_X1 T16173 ( .Y(T16173_Y));
KC_TIELO_X1 T15450 ( .Y(T15450_Y));
KC_TIELO_X1 T15448 ( .Y(T15448_Y));
KC_TIELO_X1 T15445 ( .Y(T15445_Y));
KC_TIELO_X1 T15513 ( .Y(T15513_Y));
KC_TIELO_X1 T15509 ( .Y(T15509_Y));
KC_TIELO_X1 T4870 ( .Y(T4870_Y));
KC_TIELO_X1 T15573 ( .Y(T15573_Y));
KC_TIELO_X1 T5880 ( .Y(T5880_Y));
KC_TIELO_X1 T15593 ( .Y(T15593_Y));
KC_TIELO_X1 T15585 ( .Y(T15585_Y));
KC_TIELO_X1 T15605 ( .Y(T15605_Y));
KC_TIELO_X1 T15635 ( .Y(T15635_Y));
KC_TIELO_X1 T15651 ( .Y(T15651_Y));
KC_TIELO_X1 T15674 ( .Y(T15674_Y));
KC_TIELO_X1 T15714 ( .Y(T15714_Y));
KC_TIELO_X1 T15708 ( .Y(T15708_Y));
KC_TIELO_X1 T15690 ( .Y(T15690_Y));
KC_TIELO_X1 T15820 ( .Y(T15820_Y));
KC_TIELO_X1 T15707 ( .Y(T15707_Y));
KC_TIELO_X1 T16058 ( .Y(T16058_Y));
KC_TIELO_X1 T16054 ( .Y(T16054_Y));
KC_TIELO_X1 T15822 ( .Y(T15822_Y));
KC_TIELO_X1 T15678 ( .Y(T15678_Y));
KC_TIELO_X1 T15568 ( .Y(T15568_Y));
KC_OAI22_X2 T15038 ( .A1(T3401_Y), .B0(T5875_Y), .B1(T2168_Y),     .A0(T11025_Y), .Y(T15038_Y));
KC_BUF_X14 T6497 ( .Y(T6497_Y), .A(T1825_Y));
KC_BUF_X14 T15952 ( .Y(T15952_Y), .A(T2181_Q));
KC_AO12B_X1 T102 ( .Y(T102_Y), .B(T8596_Y), .A(T13216_Q), .C(T8563_Y));
KC_AO12B_X1 T5345 ( .Y(T5345_Y), .B(T4842_Y), .A(T16184_Y),     .C(T1599_Y));
KC_AO12B_X1 T1341 ( .Y(T1341_Y), .B(T1197_Y), .A(T16309_Y),     .C(T1196_Y));
KC_AO12B_X1 T314 ( .Y(T314_Y), .B(T3070_Y), .A(T12081_Y), .C(T1418_Y));
KC_AO12B_X1 T312 ( .Y(T312_Y), .B(T12081_Y), .A(T3070_Y), .C(T1418_Y));
KC_AO12B_X1 T595 ( .Y(T595_Y), .B(T2534_Y), .A(T3070_Y), .C(T1453_Y));
KC_AO12B_X1 T579 ( .Y(T579_Y), .B(T3070_Y), .A(T2534_Y), .C(T1453_Y));
KC_AO12B_X1 T850 ( .Y(T850_Y), .B(T12328_Y), .A(T3070_Y), .C(T1492_Y));
KC_AO12B_X1 T368 ( .Y(T368_Y), .B(T12083_Y), .A(T3070_Y), .C(T1419_Y));
KC_AO12B_X1 T830 ( .Y(T830_Y), .B(T3070_Y), .A(T12328_Y), .C(T1492_Y));
KC_AO12B_X1 T6759 ( .Y(T6759_Y), .B(T3589_Y), .A(T4937_Y),     .C(T11928_Y));
KC_AO12B_X1 T1110 ( .Y(T1110_Y), .B(T3103_Y), .A(T14994_Y),     .C(T10538_Y));
KC_AO12B_X1 T5785 ( .Y(T5785_Y), .B(T2682_Y), .A(T2691_Y),     .C(T2696_Y));
KC_AO12B_X1 T5832 ( .Y(T5832_Y), .B(T5441_Q), .A(T5141_Y),     .C(T15945_Y));
KC_AO12B_X1 T5817 ( .Y(T5817_Y), .B(T2713_Q), .A(T5141_Y),     .C(T15945_Y));
KC_AO12B_X1 T5809 ( .Y(T5809_Y), .B(T2716_Q), .A(T5141_Y),     .C(T11522_Y));
KC_AO12B_X1 T5807 ( .Y(T5807_Y), .B(T2715_Q), .A(T5141_Y),     .C(T11522_Y));
KC_AO12B_X1 T5998 ( .Y(T5998_Y), .B(T2382_Q), .A(T16156_Y),     .C(T2804_Y));
KC_AO12B_X1 T5997 ( .Y(T5997_Y), .B(T2814_Q), .A(T2804_Y),     .C(T2827_Y));
KC_AO12B_X1 T6115 ( .Y(T6115_Y), .B(T10607_Y), .A(T6193_Y),     .C(T6440_Y));
KC_AO12B_X1 T858 ( .Y(T858_Y), .B(T422_Y), .A(T2648_Y), .C(T3678_Y));
KC_AO12B_X1 T6118 ( .Y(T6118_Y), .B(T3385_Y), .A(T3515_Y),     .C(T10581_Y));
KC_AO12B_X1 T15761 ( .Y(T15761_Y), .B(T10606_Y), .A(T15616_Y),     .C(T5522_Y));
KC_AO12B_X1 T1542 ( .Y(T1542_Y), .B(T12761_Y), .A(T3070_Y),     .C(T3735_Y));
KC_AO12B_X1 T6454 ( .Y(T6454_Y), .B(T422_Y), .A(T12082_Y),     .C(T3585_Y));
KC_AO12B_X1 T877 ( .Y(T877_Y), .B(T422_Y), .A(T2530_Y), .C(T4283_Y));
KC_AO12B_X1 T876 ( .Y(T876_Y), .B(T2530_Y), .A(T422_Y), .C(T4283_Y));
KC_AO12B_X1 T1522 ( .Y(T1522_Y), .B(T3070_Y), .A(T12761_Y),     .C(T3735_Y));
KC_AO12B_X1 T6166 ( .Y(T6166_Y), .B(T10614_Y), .A(T4719_Q),     .C(T6467_Y));
KC_AO12B_X1 T15758 ( .Y(T15758_Y), .B(T13323_Q), .A(T12053_Y),     .C(T4738_Y));
KC_AO12B_X1 T16273 ( .Y(T16273_Y), .B(T9889_Y), .A(T3070_Y),     .C(T1493_Y));
KC_AO12B_X1 T16272 ( .Y(T16272_Y), .B(T3070_Y), .A(T9889_Y),     .C(T1493_Y));
KC_AO12B_X1 T16370 ( .Y(T16370_Y), .B(T4934_Y), .A(T2009_Y),     .C(T5364_Q));
KC_AO12B_X1 T15866 ( .Y(T15866_Y), .B(T11373_Y), .A(T5788_Y),     .C(T11390_Y));
KC_AO12B_X1 T15759 ( .Y(T15759_Y), .B(T13324_Q), .A(T11680_Y),     .C(T4738_Y));
KC_AO12B_X1 T6453 ( .Y(T6453_Y), .B(T12082_Y), .A(T422_Y),     .C(T3025_Y));
KC_AO12B_X1 T5844 ( .Y(T5844_Y), .B(T2711_Q), .A(T5141_Y),     .C(T6228_Y));
KC_AO12B_X1 T5818 ( .Y(T5818_Y), .B(T2710_Q), .A(T5141_Y),     .C(T11522_Y));
KC_AO12B_X1 T15926 ( .Y(T15926_Y), .B(T2150_Q), .A(T5910_Y),     .C(T2722_Y));
KC_AO12B_X1 T5876 ( .Y(T5876_Y), .B(T1760_Q), .A(T5910_Y),     .C(T2145_Y));
KC_AO12B_X1 T5872 ( .Y(T5872_Y), .B(T5452_Q), .A(T5910_Y),     .C(T2165_Y));
KC_AO12B_X1 T5900 ( .Y(T5900_Y), .B(T2186_Q), .A(T5910_Y),     .C(T2140_Y));
KC_NAND3_X2 T69 ( .Y(T69_Y), .B(T15316_Y), .C(T15315_Y), .A(T8553_Y));
KC_NAND3_X2 T955 ( .Y(T955_Y), .B(T11230_Y), .C(T12885_Y),     .A(T7845_Y));
KC_NAND3_X2 T886 ( .Y(T886_Y), .B(T7848_Y), .C(T12449_Y), .A(T908_Y));
KC_NAND3_X2 T6121 ( .Y(T6121_Y), .B(T6237_Y), .C(T6556_Y),     .A(T6561_Y));
KC_NAND3_X2 T6208 ( .Y(T6208_Y), .B(T6214_Y), .C(T3478_Y),     .A(T15255_Y));
KC_NAND3_X2 T5879 ( .Y(T5879_Y), .B(T5914_Y), .C(T4515_Y),     .A(T10937_Y));
KC_AOI112B_X1 T100 ( .Y(T100_Y), .B(T15841_Y), .C1N(T132_Q),     .A(T12384_Y), .C0(T8596_Y));
KC_AOI112B_X1 T123 ( .Y(T123_Y), .B(T8608_Y), .C1N(T6932_Y),     .A(T8576_Y), .C0(T5192_Q));
KC_AOI112B_X1 T129 ( .Y(T129_Y), .B(T1144_Y), .C1N(T8974_Y),     .A(T8057_Y), .C0(T8938_Y));
KC_AOI112B_X1 T128 ( .Y(T128_Y), .B(T1144_Y), .C1N(T1127_Q),     .A(T1246_Y), .C0(T951_Y));
KC_AOI112B_X1 T140 ( .Y(T140_Y), .B(T10159_Y), .C1N(T13049_Y),     .A(T12446_Y), .C0(T10152_Y));
KC_AOI112B_X1 T86 ( .Y(T86_Y), .B(T13125_Y), .C1N(T11305_Y),     .A(T4902_Y), .C0(T12751_Y));
KC_AOI112B_X1 T148 ( .Y(T148_Y), .B(T11531_Y), .C1N(T5904_Y),     .A(T1765_Y), .C0(T11493_Y));
KC_AOI112B_X1 T94 ( .Y(T94_Y), .B(T6303_Y), .C1N(T10207_Y),     .A(T1778_Q), .C0(T10225_Y));
KC_AOI112B_X1 T142 ( .Y(T142_Y), .B(T10244_Y), .C1N(T2652_Y),     .A(T10252_Y), .C0(T5710_Y));
KC_AOI112B_X1 T15257 ( .Y(T15257_Y), .B(T13319_Y), .C1N(T10968_Y),     .A(T11801_Y), .C0(T16149_Y));
KC_AOI112B_X1 T147 ( .Y(T147_Y), .B(T3902_Y), .C1N(T12355_Y),     .A(T3903_Y), .C0(T16466_Q));
KC_AOI112B_X1 T143 ( .Y(T143_Y), .B(T5838_Y), .C1N(T4461_Y),     .A(T11976_Y), .C0(T5788_Y));
KC_AOI112B_X1 T146 ( .Y(T146_Y), .B(T13118_Y), .C1N(T10228_Y),     .A(T4494_Y), .C0(T4523_Y));
KC_AOI112B_X1 T159 ( .Y(T159_Y), .B(T11533_Y), .C1N(T3870_Y),     .A(T5969_Y), .C0(T6283_Y));
KC_AOI112B_X1 T149 ( .Y(T149_Y), .B(T11535_Y), .C1N(T11574_Y),     .A(T11533_Y), .C0(T4561_Y));
KC_AOI112B_X1 T15762 ( .Y(T15762_Y), .B(T10556_Y), .C1N(T2893_Y),     .A(T6222_Y), .C0(T8281_Y));
KC_AOI112B_X1 T15873 ( .Y(T15873_Y), .B(T11387_Y), .C1N(T4448_Y),     .A(T12954_Y), .C0(T11348_Y));
KC_AOI112B_X1 T53 ( .Y(T53_Y), .B(T15841_Y), .C1N(T6355_Q),     .A(T8546_Y), .C0(T119_Y));
KC_AOI112B_X1 T89 ( .Y(T89_Y), .B(T4494_Y), .C1N(T3880_Y),     .A(T10931_Y), .C0(T6219_Y));
KC_OAI21B_X1 T16158 ( .A0N(T9137_Y), .B(T9138_Y), .A1(T9156_Y),     .Y(T16158_Y));
KC_OAI21B_X1 T12379 ( .A0N(T69_Y), .B(T11262_Y), .A1(T16420_Y),     .Y(T12379_Y));
KC_OAI21B_X1 T12459 ( .A0N(T8109_Y), .B(T400_Y), .A1(T8088_Y),     .Y(T12459_Y));
KC_OAI21B_X1 T12390 ( .A0N(T836_Y), .B(T4853_Y), .A1(T8629_Y),     .Y(T12390_Y));
KC_OAI21B_X1 T12432 ( .A0N(T8719_Y), .B(T730_Y), .A1(T5360_Q),     .Y(T12432_Y));
KC_OAI21B_X1 T12079 ( .A0N(T7357_Y), .B(T1048_Q), .A1(T7630_Y),     .Y(T12079_Y));
KC_OAI21B_X1 T12430 ( .A0N(T9504_Y), .B(T8717_Y), .A1(T5343_Q),     .Y(T12430_Y));
KC_OAI21B_X1 T12326 ( .A0N(T7533_Y), .B(T11923_Y), .A1(T15398_Y),     .Y(T12326_Y));
KC_OAI21B_X1 T12330 ( .A0N(T16406_Y), .B(T16406_Y), .A1(T2007_Y),     .Y(T12330_Y));
KC_OAI21B_X1 T12092 ( .A0N(T9968_Y), .B(T12097_Y), .A1(T5369_Y),     .Y(T12092_Y));
KC_OAI21B_X1 T12165 ( .A0N(T11562_Y), .B(T12160_Y), .A1(T6097_S),     .Y(T12165_Y));
KC_OAI21B_X1 T12316 ( .A0N(T2321_Y), .B(T16129_Y), .A1(T2321_Y),     .Y(T12316_Y));
KC_OAI21B_X1 T12315 ( .A0N(T6570_Y), .B(T12314_Y), .A1(T6563_Y),     .Y(T12315_Y));
KC_OAI21B_X1 T12321 ( .A0N(T11824_Y), .B(T2960_Y), .A1(T11840_Y),     .Y(T12321_Y));
KC_OAI21B_X1 T12320 ( .A0N(T7836_Y), .B(T2386_Y), .A1(T6539_Y),     .Y(T12320_Y));
KC_OAI21B_X1 T12083 ( .A0N(T10493_Y), .B(T5979_Y), .A1(T4984_Y),     .Y(T12083_Y));
KC_OAI21B_X1 T12082 ( .A0N(T9779_Y), .B(T5979_Y), .A1(T4984_Y),     .Y(T12082_Y));
KC_OAI21B_X1 T12081 ( .A0N(T9874_Y), .B(T5979_Y), .A1(T4984_Y),     .Y(T12081_Y));
KC_OAI21B_X1 T12124 ( .A0N(T13062_Y), .B(T12123_Y), .A1(T2658_Y),     .Y(T12124_Y));
KC_OAI21B_X1 T12123 ( .A0N(T4381_Q), .B(T10537_Y), .A1(T16181_Y),     .Y(T12123_Y));
KC_OAI21B_X1 T12149 ( .A0N(T14957_Q), .B(T2698_Y), .A1(T15849_Y),     .Y(T12149_Y));
KC_OAI21B_X1 T12241 ( .A0N(T2811_Y), .B(T2810_Y), .A1(T2782_Y),     .Y(T12241_Y));
KC_OAI21B_X1 T12252 ( .A0N(T16055_Y), .B(T6072_Y), .A1(T2830_Y),     .Y(T12252_Y));
KC_OAI21B_X1 T12206 ( .A0N(T5921_Y), .B(T3289_Y), .A1(T3286_Y),     .Y(T12206_Y));
KC_OAI21B_X1 T12202 ( .A0N(T9227_Y), .B(T3268_Y), .A1(T11487_Y),     .Y(T12202_Y));
KC_OAI21B_X1 T12216 ( .A0N(T3324_Y), .B(T15162_Y), .A1(T3333_Y),     .Y(T12216_Y));
KC_OAI21B_X1 T12249 ( .A0N(T5492_Y), .B(T12251_Y), .A1(T3382_Y),     .Y(T12249_Y));
KC_OAI21B_X1 T12309 ( .A0N(T6575_Y), .B(T6586_Y), .A1(T11721_Y),     .Y(T12309_Y));
KC_OAI21B_X1 T12151 ( .A0N(T3851_Y), .B(T16211_Y), .A1(T3852_Y),     .Y(T12151_Y));
KC_OAI21B_X1 T12236 ( .A0N(T13145_Q), .B(T15622_Y), .A1(T3373_Y),     .Y(T12236_Y));
KC_OAI21B_X1 T12290 ( .A0N(T4058_Y), .B(T15619_Y), .A1(T10581_Y),     .Y(T12290_Y));
KC_OAI21B_X1 T12144 ( .A0N(T11349_Y), .B(T11346_Y), .A1(T3833_Y),     .Y(T12144_Y));
KC_OAI21B_X1 T12209 ( .A0N(T4601_Y), .B(T5934_Y), .A1(T4524_Y),     .Y(T12209_Y));
KC_OAI21B_X1 T12197 ( .A0N(T4524_Y), .B(T12810_Y), .A1(T5884_Y),     .Y(T12197_Y));
KC_OAI21B_X1 T12352 ( .A0N(T3940_Y), .B(T15965_Y), .A1(T4563_Y),     .Y(T12352_Y));
KC_OAI21B_X1 T12237 ( .A0N(T5485_Y), .B(T4615_Y), .A1(T3982_Y),     .Y(T12237_Y));
KC_OAI21B_X1 T12328 ( .A0N(T9747_Y), .B(T5979_Y), .A1(T4984_Y),     .Y(T12328_Y));
KC_OAI21B_X1 T12070 ( .A0N(T1_Y), .B(T6845_Y), .A1(T287_Y),     .Y(T12070_Y));
KC_OAI21B_X1 T12349 ( .A0N(T6025_Y), .B(T6340_Y), .A1(T15996_Y),     .Y(T12349_Y));
KC_OAI21B_X1 T12142 ( .A0N(T14526_Q), .B(T10904_Y), .A1(T5427_Y),     .Y(T12142_Y));
KC_OAI21B_X1 T12204 ( .A0N(T5458_Y), .B(T13115_Y), .A1(T3936_Q),     .Y(T12204_Y));
KC_OAI21B_X1 T12194 ( .A0N(T4539_Y), .B(T3939_Y), .A1(T9487_Y),     .Y(T12194_Y));
KC_MXI2_X2 T10884 ( .Y(T10884_Y), .A(T5480_Q), .S0(T15014_Y),     .B(T11446_Y));
KC_MXI2_X2 T10883 ( .Y(T10883_Y), .A(T2809_Q), .S0(T15014_Y),     .B(T5042_Y));
KC_MXI2_X2 T10942 ( .Y(T10942_Y), .A(T6555_Q), .S0(T3294_Y),     .B(T3909_Y));
KC_MXI2_X2 T10941 ( .Y(T10941_Y), .A(T6549_Q), .S0(T3294_Y),     .B(T3908_Y));
KC_MXI2_X2 T10880 ( .Y(T10880_Y), .A(T6526_Q), .S0(T3294_Y),     .B(T3910_Y));
KC_MXI2_X2 T10918 ( .Y(T10918_Y), .A(T8306_Y), .S0(T15014_Y),     .B(T5844_Y));
KC_MXI2_X2 T10916 ( .Y(T10916_Y), .A(T16018_Q), .S0(T15014_Y),     .B(T3251_Y));
KC_MXI2_X2 T10912 ( .Y(T10912_Y), .A(T5481_Q), .S0(T15014_Y),     .B(T5818_Y));
KC_MXI2_X2 T10906 ( .Y(T10906_Y), .A(T5987_Q), .S0(T15014_Y),     .B(T11445_Y));
KC_MXI2_X2 T10934 ( .Y(T10934_Y), .A(T5530_Q), .S0(T3294_Y),     .B(T5484_Y));
KC_MXI2_X2 T11016 ( .Y(T11016_Y), .A(T15990_Q), .S0(T15014_Y),     .B(T5807_Y));
KC_MXI2_X2 T11011 ( .Y(T11011_Y), .A(T16010_Q), .S0(T15014_Y),     .B(T11434_Y));
KC_MXI2_X2 T11010 ( .Y(T11010_Y), .A(T16007_Q), .S0(T15014_Y),     .B(T3865_Y));
KC_MXI2_X2 T10917 ( .Y(T10917_Y), .A(T16025_Y), .S0(T15014_Y),     .B(T5832_Y));
KC_MXI2_X2 T10907 ( .Y(T10907_Y), .A(T16023_Q), .S0(T15014_Y),     .B(T5809_Y));
KC_MXI2_X2 T10905 ( .Y(T10905_Y), .A(T2237_Q), .S0(T15014_Y),     .B(T5817_Y));
KC_MXI2_X2 T10936 ( .Y(T10936_Y), .A(T15760_Q), .S0(T3294_Y),     .B(T5459_Y));
KC_OR2_X1 T5588 ( .Y(T5588_Y), .A(T45_Q), .B(T5586_Q));
KC_OR2_X1 T116 ( .Y(T116_Y), .A(T5630_Y), .B(T14971_Y));
KC_OR2_X1 T119 ( .Y(T119_Y), .A(T33_Y), .B(T15312_Y));
KC_OR2_X1 T126 ( .Y(T126_Y), .A(T33_Y), .B(T5614_Y));
KC_OR2_X1 T137 ( .Y(T137_Y), .A(T9272_Y), .B(T12382_Y));
KC_OR2_X1 T229 ( .Y(T229_Y), .A(T9270_Y), .B(T9395_Y));
KC_OR2_X1 T482 ( .Y(T482_Y), .A(T9282_Y), .B(T7056_Y));
KC_OR2_X1 T538 ( .Y(T538_Y), .A(T11230_Y), .B(T15841_Y));
KC_OR2_X1 T560 ( .Y(T560_Y), .A(T8130_Y), .B(T1350_Y));
KC_OR2_X1 T590 ( .Y(T590_Y), .A(T1839_Y), .B(T16183_Y));
KC_OR2_X1 T655 ( .Y(T655_Y), .A(T7050_Y), .B(T7112_Y));
KC_OR2_X1 T661 ( .Y(T661_Y), .A(T9275_Y), .B(T7051_Y));
KC_OR2_X1 T678 ( .Y(T678_Y), .A(T7241_Y), .B(T7299_Y));
KC_OR2_X1 T745 ( .Y(T745_Y), .A(T10738_Y), .B(T757_Y));
KC_OR2_X1 T840 ( .Y(T840_Y), .A(T836_Y), .B(T833_Y));
KC_OR2_X1 T961 ( .Y(T961_Y), .A(T9438_Y), .B(T10142_Y));
KC_OR2_X1 T1149 ( .Y(T1149_Y), .A(T15014_Y), .B(T16040_Y));
KC_OR2_X1 T1288 ( .Y(T1288_Y), .A(T13198_Q), .B(T15544_Y));
KC_OR2_X1 T1368 ( .Y(T1368_Y), .A(T1363_Y), .B(T4819_Y));
KC_OR2_X1 T1379 ( .Y(T1379_Y), .A(T8395_Y), .B(T16120_Y));
KC_OR2_X1 T1555 ( .Y(T1555_Y), .A(T7780_Y), .B(T10756_Y));
KC_OR2_X1 T1773 ( .Y(T1773_Y), .A(T11530_Y), .B(T11502_Y));
KC_OR2_X1 T2014 ( .Y(T2014_Y), .A(T1162_Y), .B(T2024_Y));
KC_OR2_X1 T2055 ( .Y(T2055_Y), .A(T16295_Y), .B(T10085_Y));
KC_OR2_X1 T2060 ( .Y(T2060_Y), .A(T12736_Y), .B(T1509_Y));
KC_OR2_X1 T2188 ( .Y(T2188_Y), .A(T8242_Y), .B(T2167_Y));
KC_OR2_X1 T2243 ( .Y(T2243_Y), .A(T13152_Y), .B(T6013_Y));
KC_OR2_X1 T2244 ( .Y(T2244_Y), .A(T13152_Y), .B(T3306_Y));
KC_OR2_X1 T2274 ( .Y(T2274_Y), .A(T11665_Y), .B(T5878_Y));
KC_OR2_X1 T2309 ( .Y(T2309_Y), .A(T3214_Y), .B(T2276_Q));
KC_OR2_X1 T2346 ( .Y(T2346_Y), .A(T2824_Y), .B(T6566_Y));
KC_OR2_X1 T2394 ( .Y(T2394_Y), .A(T2396_Y), .B(T2396_Y));
KC_OR2_X1 T2573 ( .Y(T2573_Y), .A(T16363_Y), .B(T16412_Y));
KC_OR2_X1 T10239 ( .Y(T10239_Y), .A(T10243_Y), .B(T2665_Y));
KC_OR2_X1 T2668 ( .Y(T2668_Y), .A(T10271_Y), .B(T10244_Y));
KC_OR2_X1 T2758 ( .Y(T2758_Y), .A(T2762_Y), .B(T3284_Y));
KC_OR2_X1 T2837 ( .Y(T2837_Y), .A(T5512_Q), .B(T4048_Q));
KC_OR2_X1 T2872 ( .Y(T2872_Y), .A(T12276_Y), .B(T5053_Y));
KC_OR2_X1 T2961 ( .Y(T2961_Y), .A(T11000_Y), .B(T4055_Y));
KC_OR2_X1 T3062 ( .Y(T3062_Y), .A(T5270_Y), .B(T2496_Y));
KC_OR2_X1 T3230 ( .Y(T3230_Y), .A(T11357_Y), .B(T15896_Y));
KC_OR2_X1 T3309 ( .Y(T3309_Y), .A(T3345_Y), .B(T6230_Co));
KC_OR2_X1 T3337 ( .Y(T3337_Y), .A(T11557_Y), .B(T3325_Y));
KC_OR2_X1 T3361 ( .Y(T3361_Y), .A(T8325_Y), .B(T15607_Y));
KC_OR2_X1 T3498 ( .Y(T3498_Y), .A(T10990_Y), .B(T10544_Y));
KC_OR2_X1 T3922 ( .Y(T3922_Y), .A(T3924_Y), .B(T6797_Co));
KC_OR2_X1 T3923 ( .Y(T3923_Y), .A(T15932_Y), .B(T3904_Y));
KC_OR2_X1 T3924 ( .Y(T3924_Y), .A(T3265_Y), .B(T11495_Y));
KC_OR2_X1 T4010 ( .Y(T4010_Y), .A(T16455_Q), .B(T4622_Y));
KC_OR2_X1 T4105 ( .Y(T4105_Y), .A(T3368_Y), .B(T4062_Y));
KC_OR2_X1 T4499 ( .Y(T4499_Y), .A(T11442_Y), .B(T5854_Y));
KC_OR2_X1 T4522 ( .Y(T4522_Y), .A(T5156_Y), .B(T12197_Y));
KC_OR2_X1 T4525 ( .Y(T4525_Y), .A(T4526_Q), .B(T4528_Q));
KC_OR2_X1 T4533 ( .Y(T4533_Y), .A(T5885_Y), .B(T8244_Y));
KC_OR2_X1 T4563 ( .Y(T4563_Y), .A(T15970_Y), .B(T4411_Y));
KC_OR2_X1 T4688 ( .Y(T4688_Y), .A(T16112_Y), .B(T4692_Y));
KC_OR2_X1 T4709 ( .Y(T4709_Y), .A(T16122_Y), .B(T4724_Y));
KC_OR2_X1 T4710 ( .Y(T4710_Y), .A(T6169_Y), .B(T8390_Y));
KC_OR2_X1 T4744 ( .Y(T4744_Y), .A(T12307_Y), .B(T4729_Y));
KC_OR2_X1 T4752 ( .Y(T4752_Y), .A(T4731_Y), .B(T4734_Y));
KC_OR2_X1 T4820 ( .Y(T4820_Y), .A(T9450_Y), .B(T9071_Y));
KC_OR2_X1 T4821 ( .Y(T4821_Y), .A(T1427_Y), .B(T15097_Y));
KC_OR2_X1 T4829 ( .Y(T4829_Y), .A(T390_Y), .B(T4821_Y));
KC_OR2_X1 T4833 ( .Y(T4833_Y), .A(T9280_Y), .B(T7060_Y));
KC_OR2_X1 T15733 ( .Y(T15733_Y), .A(T7443_Y), .B(T9336_Y));
KC_OR2_X1 T4839 ( .Y(T4839_Y), .A(T9509_Y), .B(T9315_Y));
KC_OR2_X1 T5061 ( .Y(T5061_Y), .A(T11591_Y), .B(T3319_Y));
KC_OR2_X1 T5080 ( .Y(T5080_Y), .A(T2676_Y), .B(T2467_Y));
KC_OR2_X1 T5123 ( .Y(T5123_Y), .A(T12349_Y), .B(T6340_Y));
KC_OR2_X1 T5152 ( .Y(T5152_Y), .A(T4717_Q), .B(T6171_Y));
KC_OR2_X1 T5157 ( .Y(T5157_Y), .A(T4573_Q), .B(T15703_Y));
KC_OR2_X1 T5244 ( .Y(T5244_Y), .A(T9285_Y), .B(T7068_Y));
KC_OR2_X1 T601 ( .Y(T601_Y), .A(T9337_Y), .B(T9335_Y));
KC_OR2_X1 T5460 ( .Y(T5460_Y), .A(T1760_Q), .B(T2186_Q));
KC_MXI2B_X4 T9115 ( .Y(T9115_Y), .A(T9127_Y), .BN(T427_Y),     .S0(T957_Y));
KC_MXI2B_X4 T139 ( .Y(T139_Y), .A(T7877_Y), .BN(T9393_Y), .S0(T980_Q));
KC_MXI2B_X4 T16113 ( .Y(T16113_Y), .A(T864_Y), .BN(T5825_S),     .S0(T881_Y));
KC_MXI2B_X4 T15702 ( .Y(T15702_Y), .A(T16294_Y), .BN(T2618_Q),     .S0(T12738_Y));
KC_MXI2B_X4 T15444 ( .Y(T15444_Y), .A(T8230_Y), .BN(T11468_Y),     .S0(T3259_Y));
KC_MXI2B_X4 T9227 ( .Y(T9227_Y), .A(T12201_Y), .BN(T13120_Y),     .S0(T8246_Y));
KC_MXI2B_X4 T7915 ( .Y(T7915_Y), .A(T16015_Y), .BN(T6024_Y),     .S0(T3351_Y));
KC_MXI2B_X4 T9163 ( .Y(T9163_Y), .A(T4151_Y), .BN(T4173_Y),     .S0(T4156_Y));
KC_MXI2B_X4 T5044 ( .Y(T5044_Y), .A(T15160_Y), .BN(T4447_Y),     .S0(T15874_Y));
KC_MXI2B_X4 T4708 ( .Y(T4708_Y), .A(T15572_Y), .BN(T11466_Y),     .S0(T5873_Y));
KC_MXI2B_X4 T9100 ( .Y(T9100_Y), .A(T4738_Y), .BN(T13167_Q),     .S0(T5151_Y));
KC_MXI2B_X4 T5469 ( .Y(T5469_Y), .A(T15694_Y), .BN(T14530_Q),     .S0(T16160_Y));
KC_MXI2B_X4 T88 ( .Y(T88_Y), .A(T12451_Y), .BN(T7916_Y), .S0(T8080_Y));
KC_MXI2B_X4 T4411 ( .Y(T4411_Y), .A(T15987_Y), .BN(T4552_Y),     .S0(T15986_Y));
KC_XOR2_X3 T13215 ( .A(T6853_Y), .B(T13068_Y), .Y(T13215_Y));
KC_XOR2_X3 T13214 ( .A(T6854_Y), .B(T13068_Y), .Y(T13214_Y));
KC_XOR2_X3 T13213 ( .A(T5646_Y), .B(T13075_Y), .Y(T13213_Y));
KC_XOR2_X3 T13212 ( .A(T5645_Y), .B(T13075_Y), .Y(T13212_Y));
KC_XOR2_X3 T13231 ( .A(T5621_Y), .B(T15321_Y), .Y(T13231_Y));
KC_XOR2_X3 T13230 ( .A(T5610_Y), .B(T70_Y), .Y(T13230_Y));
KC_XOR2_X3 T13225 ( .A(T72_Y), .B(T70_Y), .Y(T13225_Y));
KC_XOR2_X3 T13224 ( .A(T5620_Y), .B(T15321_Y), .Y(T13224_Y));
KC_XOR2_X3 T13236 ( .A(T7459_Y), .B(T15407_Y), .Y(T13236_Y));
KC_XOR2_X3 T13235 ( .A(T7433_Y), .B(T15407_Y), .Y(T13235_Y));
KC_XOR2_X3 T13223 ( .A(T7116_Y), .B(T15369_Y), .Y(T13223_Y));
KC_XOR2_X3 T13222 ( .A(T7117_Y), .B(T15369_Y), .Y(T13222_Y));
KC_XOR2_X3 T13259 ( .A(T16282_Y), .B(T16282_Y), .Y(T13259_Y));
KC_XOR2_X3 T13252 ( .A(T8040_Y), .B(T15484_Y), .Y(T13252_Y));
KC_XOR2_X3 T13251 ( .A(T8039_Y), .B(T15484_Y), .Y(T13251_Y));
KC_XOR2_X3 T13228 ( .A(T6857_Y), .B(T15335_Y), .Y(T13228_Y));
KC_XOR2_X3 T13227 ( .A(T6858_Y), .B(T15335_Y), .Y(T13227_Y));
KC_XOR2_X3 T13234 ( .A(T7406_Y), .B(T15411_Y), .Y(T13234_Y));
KC_XOR2_X3 T12989 ( .A(T7183_Y), .B(T15673_Y), .Y(T12989_Y));
KC_XOR2_X3 T13199 ( .A(T10039_Y), .B(T15496_Y), .Y(T13199_Y));
KC_XOR2_X3 T13034 ( .A(T10020_Y), .B(T15496_Y), .Y(T13034_Y));
KC_XOR2_X3 T12987 ( .A(T6891_Y), .B(T15342_Y), .Y(T12987_Y));
KC_XOR2_X3 T12986 ( .A(T6870_Y), .B(T15342_Y), .Y(T12986_Y));
KC_XOR2_X3 T13204 ( .A(T10336_Y), .B(T15415_Y), .Y(T13204_Y));
KC_XOR2_X3 T13004 ( .A(T7534_Y), .B(T15415_Y), .Y(T13004_Y));
KC_XOR2_X3 T12990 ( .A(T7186_Y), .B(T8671_Y), .Y(T12990_Y));
KC_XOR2_X3 T12988 ( .A(T10400_Y), .B(T8671_Y), .Y(T12988_Y));
KC_XOR2_X3 T12996 ( .A(T5705_Y), .B(T15347_Y), .Y(T12996_Y));
KC_XOR2_X3 T13302 ( .A(T4354_Y), .B(T10643_Y), .Y(T13302_Y));
KC_XOR2_X3 T13301 ( .A(T10900_Y), .B(T8448_Y), .Y(T13301_Y));
KC_XOR2_X3 T13152 ( .A(T3306_Y), .B(T6013_Y), .Y(T13152_Y));
KC_XOR2_X3 T13197 ( .A(T12879_Y), .B(T2369_Y), .Y(T13197_Y));
KC_XOR2_X3 T12995 ( .A(T5742_Y), .B(T15381_Y), .Y(T12995_Y));
KC_XOR2_X3 T12992 ( .A(T5727_Y), .B(T15381_Y), .Y(T12992_Y));
KC_XOR2_X3 T13044 ( .A(T5916_Y), .B(T16303_Y), .Y(T13044_Y));
KC_XOR2_X3 T13142 ( .A(T11491_Y), .B(T11478_Y), .Y(T13142_Y));
KC_XOR2_X3 T13137 ( .A(T2784_Y), .B(T5978_Y), .Y(T13137_Y));
KC_XOR2_X3 T13061 ( .A(T6002_Y), .B(T15551_Y), .Y(T13061_Y));
KC_XOR2_X3 T13069 ( .A(T15826_Y), .B(T12776_Y), .Y(T13069_Y));
KC_XOR2_X3 T13095 ( .A(T6110_Y), .B(T15565_Y), .Y(T13095_Y));
KC_XOR2_X3 T13094 ( .A(T6122_Y), .B(T15565_Y), .Y(T13094_Y));
KC_XOR2_X3 T13120 ( .A(T5893_Y), .B(T8267_Y), .Y(T13120_Y));
KC_XOR2_X3 T13139 ( .A(T11548_Y), .B(T15962_Y), .Y(T13139_Y));
KC_XOR2_X3 T13147 ( .A(T6306_Y), .B(T4352_Y), .Y(T13147_Y));
KC_XOR2_X3 T13181 ( .A(T6843_Y), .B(T15639_Y), .Y(T13181_Y));
KC_XOR2_X3 T13192 ( .A(T6596_Y), .B(T15639_Y), .Y(T13192_Y));
KC_XOR2_X3 T13206 ( .A(T6669_Y), .B(T3290_Y), .Y(T13206_Y));
KC_XOR2_X3 T13011 ( .A(T3707_Y), .B(T857_Y), .Y(T13011_Y));
KC_XOR2_X3 T13138 ( .A(T6287_Y), .B(T15594_Y), .Y(T13138_Y));
KC_XOR2_X3 T13153 ( .A(T4594_Y), .B(T4605_Y), .Y(T13153_Y));
KC_XOR2_X3 T13146 ( .A(T6307_Y), .B(T4352_Y), .Y(T13146_Y));
KC_XOR2_X3 T12985 ( .A(T5711_Y), .B(T15366_Y), .Y(T12985_Y));
KC_XOR2_X3 T12984 ( .A(T5722_Y), .B(T15366_Y), .Y(T12984_Y));
KC_XOR2_X3 T12993 ( .A(T6627_Y), .B(T6455_Y), .Y(T12993_Y));
KC_XOR2_X3 T12991 ( .A(T6626_Y), .B(T6455_Y), .Y(T12991_Y));
KC_XOR2_X3 T13045 ( .A(T5396_Y), .B(T2724_Y), .Y(T13045_Y));
KC_XOR2_X3 T13043 ( .A(T5912_Y), .B(T2724_Y), .Y(T13043_Y));
KC_XOR2_X3 T13208 ( .A(T6677_Y), .B(T6848_Y), .Y(T13208_Y));
KC_XOR2_X3 T13290 ( .A(T6001_Y), .B(T15551_Y), .Y(T13290_Y));
KC_XOR2_X3 T13207 ( .A(T5831_Y), .B(T3290_Y), .Y(T13207_Y));
KC_XOR2_X3 T13315 ( .A(T12353_Y), .B(T15938_Y), .Y(T13315_Y));
KC_XOR2_X3 T12994 ( .A(T5707_Y), .B(T15347_Y), .Y(T12994_Y));
KC_XOR2_X3 T12997 ( .A(T10405_Y), .B(T15673_Y), .Y(T12997_Y));
KC_XOR2_X3 T13271 ( .A(T7390_Y), .B(T15411_Y), .Y(T13271_Y));
KC_XOR2_X3 T13005 ( .A(T5796_Y), .B(T6848_Y), .Y(T13005_Y));
KC_XOR2_X3 T13024 ( .A(T7979_Y), .B(T984_Y), .Y(T13024_Y));
KC_XOR2_X3 T13021 ( .A(T10304_Y), .B(T984_Y), .Y(T13021_Y));
KC_XOR2_X3 T13258 ( .A(T427_Y), .B(T957_Y), .Y(T13258_Y));
KC_XOR2_X3 T13041 ( .A(T5915_Y), .B(T16303_Y), .Y(T13041_Y));
KC_XOR2_X3 T12979 ( .A(T6788_Y), .B(T15594_Y), .Y(T12979_Y));
KC_OR4_X1 T8550 ( .Y(T8550_Y), .C(T52_Y), .B(T13294_Y), .D(T5184_Q),     .A(T5588_Y));
KC_OR4_X1 T8561 ( .Y(T8561_Y), .C(T12371_Y), .B(T79_Y), .D(T5629_Y),     .A(T5184_Q));
KC_OR4_X1 T9024 ( .Y(T9024_Y), .C(T9080_Co), .B(T15077_Y), .D(T9080_S),     .A(T9080_Co));
KC_OR4_X1 T8869 ( .Y(T8869_Y), .C(T7917_Y), .B(T12451_Y), .D(T7862_Y),     .A(T12451_Y));
KC_OR4_X1 T8629 ( .Y(T8629_Y), .C(T6250_Y), .B(T11085_Y), .D(T16510_Y),     .A(T833_Y));
KC_OR4_X1 T10228 ( .Y(T10228_Y), .C(T1165_Y), .B(T1277_Y), .D(T9223_Y),     .A(T1166_Y));
KC_OR4_X1 T10315 ( .Y(T10315_Y), .C(T5341_Q), .B(T5337_Q), .D(T1210_Q),     .A(T5340_Q));
KC_OR4_X1 T10313 ( .Y(T10313_Y), .C(T1195_Q), .B(T1221_Q), .D(T1224_Q),     .A(T1231_Q));
KC_OR4_X1 T9925 ( .Y(T9925_Y), .C(T1188_Q), .B(T1203_Q), .D(T4869_Q),     .A(T1215_Q));
KC_OR4_X1 T9914 ( .Y(T9914_Y), .C(T1211_Q), .B(T1207_Q), .D(T1212_Q),     .A(T1208_Q));
KC_OR4_X1 T9895 ( .Y(T9895_Y), .C(T1216_Q), .B(T1209_Q), .D(T1202_Q),     .A(T1190_Q));
KC_OR4_X1 T10021 ( .Y(T10021_Y), .C(T1223_Q), .B(T1232_Q), .D(T1222_Q),     .A(T1220_Q));
KC_OR4_X1 T8342 ( .Y(T8342_Y), .C(T1781_Y), .B(T1771_Y), .D(T4911_Y),     .A(T1780_Y));
KC_OR4_X1 T10183 ( .Y(T10183_Y), .C(T2070_Y), .B(T10185_Y),     .D(T6593_Y), .A(T2069_Y));
KC_OR4_X1 T10253 ( .Y(T10253_Y), .C(T4010_Y), .B(T2082_Q), .D(T2768_Y),     .A(T2006_Y));
KC_OR4_X1 T8326 ( .Y(T8326_Y), .C(T8315_Y), .B(T8339_Y), .D(T8341_Y),     .A(T8327_Y));
KC_OR4_X1 T8318 ( .Y(T8318_Y), .C(T8310_Y), .B(T8282_Y), .D(T8309_Y),     .A(T8319_Y));
KC_OR4_X1 T8317 ( .Y(T8317_Y), .C(T8473_Y), .B(T8328_Y), .D(T8240_Y),     .A(T8343_Y));
KC_OR4_X1 T8157 ( .Y(T8157_Y), .C(T2367_Y), .B(T6492_Y), .D(T6492_Y),     .A(T6492_Y));
KC_OR4_X1 T8453 ( .Y(T8453_Y), .C(T2837_Y), .B(T10895_Y), .D(T11530_Y),     .A(T5015_Q));
KC_OR4_X1 T8198 ( .Y(T8198_Y), .C(T2706_Y), .B(T2124_Y), .D(T2124_Y),     .A(T16152_Y));
KC_OR4_X1 T8378 ( .Y(T8378_Y), .C(T10986_Y), .B(T10556_Y), .D(T2885_Y),     .A(T10594_Y));
KC_OR4_X1 T8246 ( .Y(T8246_Y), .C(T5890_Y), .B(T3312_Y), .D(T6231_Co),     .A(T3295_Y));
KC_OR4_X1 T8332 ( .Y(T8332_Y), .C(T3979_Y), .B(T5123_Y), .D(T10953_Y),     .A(T5124_Y));
KC_OR4_X1 T8467 ( .Y(T8467_Y), .C(T12064_Y), .B(T5009_Y), .D(T2812_Y),     .A(T3423_Y));
KC_OR4_X1 T8163 ( .Y(T8163_Y), .C(T4180_Y), .B(T4761_Y), .D(T4761_Y),     .A(T4662_Y));
KC_OR4_X1 T8455 ( .Y(T8455_Y), .C(T5150_Y), .B(T4692_Y), .D(T4638_Y),     .A(T12345_Y));
KC_OR4_X1 T9322 ( .Y(T9322_Y), .C(T164_Q), .B(T165_Q), .D(T163_Q),     .A(T4837_Q));
KC_OR4_X1 T10536 ( .Y(T10536_Y), .C(T15689_Y), .B(T15689_Y),     .D(T15689_Y), .A(T15689_Y));
KC_OR4_X1 T9094 ( .Y(T9094_Y), .C(T9460_Q), .B(T5407_Q), .D(T9461_Q),     .A(T998_Q));
KC_OR4_X1 T8281 ( .Y(T8281_Y), .C(T13127_Q), .B(T13136_Q),     .D(T13129_Q), .A(T13133_Q));
KC_AO21_X1 T1448 ( .A0(T9080_Co), .B(T9024_Y), .Y(T1448_Y),     .A1(T9451_Y));
KC_AO21_X1 T1446 ( .A0(T1602_Y), .B(T1367_Y), .Y(T1446_Y),     .A1(T15091_Y));
KC_AO21_X1 T1445 ( .A0(T16284_Y), .B(T16087_Y), .Y(T1445_Y),     .A1(T9025_Y));
KC_AO21_X1 T7647 ( .A0(T722_Q), .B(T8895_Y), .Y(T7647_Y), .A1(T714_Q));
KC_AO21_X1 T8041 ( .A0(T8059_Y), .B(T8070_Y), .Y(T8041_Y),     .A1(T9007_Y));
KC_AO21_X1 T16188 ( .A0(T4842_Y), .B(T16186_Y), .Y(T16188_Y),     .A1(T9474_Y));
KC_AO21_X1 T4805 ( .A0(T9442_Y), .B(T9098_Y), .Y(T4805_Y),     .A1(T231_Y));
KC_AO21_X1 T1739 ( .A0(T9442_Y), .B(T9040_Y), .Y(T1739_Y),     .A1(T240_Y));
KC_AO21_X1 T1732 ( .A0(T9442_Y), .B(T9036_Y), .Y(T1732_Y),     .A1(T6800_Y));
KC_AO21_X1 T1697 ( .A0(T9442_Y), .B(T9035_Y), .Y(T1697_Y),     .A1(T9488_Y));
KC_AO21_X1 T1634 ( .A0(T9442_Y), .B(T9095_Y), .Y(T1634_Y),     .A1(T9101_Y));
KC_AO21_X1 T1567 ( .A0(T9442_Y), .B(T9049_Y), .Y(T1567_Y),     .A1(T9066_Y));
KC_AO21_X1 T10738 ( .A0(T15014_Y), .B(T1013_Q), .Y(T10738_Y),     .A1(T5879_Y));
KC_AO21_X1 T10724 ( .A0(T1738_Y), .B(T1357_Y), .Y(T10724_Y),     .A1(T1368_Y));
KC_AO21_X1 T5968 ( .A0(T16237_Y), .B(T10183_Y), .Y(T5968_Y),     .A1(T2070_Y));
KC_AO21_X1 T6605 ( .A0(T4978_Y), .B(T2374_Y), .Y(T6605_Y),     .A1(T2393_Y));
KC_AO21_X1 T5849 ( .A0(T2507_Y), .B(T12085_Y), .Y(T5849_Y),     .A1(T5314_Y));
KC_AO21_X1 T5994 ( .A0(T14495_Q), .B(T15827_Y), .Y(T5994_Y),     .A1(T16172_Y));
KC_AO21_X1 T5993 ( .A0(T14494_Q), .B(T15827_Y), .Y(T5993_Y),     .A1(T2659_Y));
KC_AO21_X1 T5988 ( .A0(T16160_Y), .B(T12115_Y), .Y(T5988_Y),     .A1(T16079_Q));
KC_AO21_X1 T6154 ( .A0(T2738_Q), .B(T11471_Y), .Y(T6154_Y),     .A1(T4991_Y));
KC_AO21_X1 T6153 ( .A0(T2737_Q), .B(T11470_Y), .Y(T6153_Y),     .A1(T4991_Y));
KC_AO21_X1 T6152 ( .A0(T2748_Q), .B(T11471_Y), .Y(T6152_Y),     .A1(T4991_Y));
KC_AO21_X1 T6279 ( .A0(T5978_Y), .B(T2786_Y), .Y(T6279_Y),     .A1(T2789_Y));
KC_AO21_X1 T6367 ( .A0(T11632_Y), .B(T2846_Y), .Y(T6367_Y),     .A1(T2831_Y));
KC_AO21_X1 T2930 ( .A0(T2931_Y), .B(T5535_Y), .Y(T2930_Y),     .A1(T11844_Y));
KC_AO21_X1 T6278 ( .A0(T3363_Y), .B(T3316_Y), .Y(T6278_Y),     .A1(T15591_Y));
KC_AO21_X1 T6574 ( .A0(T11804_Y), .B(T11795_Y), .Y(T6574_Y),     .A1(T3394_Y));
KC_AO21_X1 T6645 ( .A0(T10457_Y), .B(T15365_Y), .Y(T6645_Y),     .A1(T6438_Y));
KC_AO21_X1 T5712 ( .A0(T6438_Y), .B(T5713_Y), .Y(T5712_Y),     .A1(T10457_Y));
KC_AO21_X1 T6136 ( .A0(T4501_Y), .B(T6127_Y), .Y(T6136_Y),     .A1(T4502_Y));
KC_AO21_X1 T6283 ( .A0(T11539_Y), .B(T12015_Y), .Y(T6283_Y),     .A1(T5155_Y));
KC_AO21_X1 T6360 ( .A0(T4690_Y), .B(T8366_Y), .Y(T6360_Y),     .A1(T4687_Y));
KC_AO21_X1 T6421 ( .A0(T13165_Q), .B(T6090_Y), .Y(T6421_Y),     .A1(T5144_Y));
KC_AO21_X1 T16282 ( .A0(T4821_Y), .B(T4829_Y), .Y(T16282_Y),     .A1(T390_Y));
KC_AO21_X1 T6844 ( .A0(T6545_Y), .B(T5029_Y), .Y(T6844_Y),     .A1(T6545_Y));
KC_AO21_X1 T6736 ( .A0(T2749_Q), .B(T11470_Y), .Y(T6736_Y),     .A1(T4991_Y));
KC_AO21_X1 T6707 ( .A0(T2669_Q), .B(T10256_Y), .Y(T6707_Y),     .A1(T10204_Y));
KC_AO21_X1 T6241 ( .A0(T6251_Y), .B(T3975_Y), .Y(T6241_Y),     .A1(T4569_Y));
KC_SDFFRNHQ_X1 T15286 ( .Q(T15286_Q), .SI(T13214_Y), .D(T15286_Q),     .SE(T15329_Y), .RN(T14970_Y), .CK(T15165_Y));
KC_SDFFRNHQ_X1 T15284 ( .Q(T15284_Q), .SI(T13215_Y), .D(T15284_Q),     .SE(T15329_Y), .RN(T14970_Y), .CK(T6852_Y));
KC_SDFFRNHQ_X1 T15285 ( .Q(T15285_Q), .SI(T13213_Y), .D(T15285_Q),     .SE(T13074_Y), .RN(T14970_Y), .CK(T6851_Y));
KC_SDFFRNHQ_X1 T15288 ( .Q(T15288_Q), .SI(T13230_Y), .D(T15288_Q),     .SE(T13080_Y), .RN(T14970_Y), .CK(T5626_Y));
KC_SDFFRNHQ_X1 T15287 ( .Q(T15287_Q), .SI(T13225_Y), .D(T15287_Q),     .SE(T13080_Y), .RN(T14970_Y), .CK(T5635_Y));
KC_SDFFRNHQ_X1 T5594 ( .Q(T5594_Q), .SI(T13224_Y), .D(T5594_Q),     .SE(T15170_Y), .RN(T15024_Y), .CK(T5638_Y));
KC_SDFFRNHQ_X1 T28 ( .Q(T28_Q), .SI(T13231_Y), .D(T28_Q),     .SE(T15170_Y), .RN(T15024_Y), .CK(T5632_Y));
KC_SDFFRNHQ_X1 T15307 ( .Q(T15307_Q), .SI(T13236_Y), .D(T15307_Q),     .SE(T15653_Y), .RN(T7609_Y), .CK(T7608_Y));
KC_SDFFRNHQ_X1 T15299 ( .Q(T15299_Q), .SI(T13235_Y), .D(T15299_Q),     .SE(T570_Y), .RN(T7609_Y), .CK(T7405_Y));
KC_SDFFRNHQ_X1 T15292 ( .Q(T15292_Q), .SI(T13222_Y), .D(T15292_Q),     .SE(T15368_Y), .RN(T7242_Y), .CK(T7101_Y));
KC_SDFFRNHQ_X1 T15291 ( .Q(T15291_Q), .SI(T13223_Y), .D(T15291_Q),     .SE(T15368_Y), .RN(T7242_Y), .CK(T7094_Y));
KC_SDFFRNHQ_X1 T15305 ( .Q(T15305_Q), .SI(T13251_Y), .D(T15305_Q),     .SE(T15483_Y), .RN(T14997_Y), .CK(T8043_Y));
KC_SDFFRNHQ_X1 T15304 ( .Q(T15304_Q), .SI(T13252_Y), .D(T15304_Q),     .SE(T15483_Y), .RN(T14997_Y), .CK(T8068_Y));
KC_SDFFRNHQ_X1 T115 ( .Q(T115_Q), .SI(T13227_Y), .D(T115_Q),     .SE(T15334_Y), .RN(T837_Y), .CK(T118_Y));
KC_SDFFRNHQ_X1 T15289 ( .Q(T15289_Q), .SI(T13228_Y), .D(T15289_Q),     .SE(T15649_Y), .RN(T837_Y), .CK(T225_Y));
KC_SDFFRNHQ_X1 T15302 ( .Q(T15302_Q), .SI(T13199_Y), .D(T15302_Q),     .SE(T15460_Y), .RN(T1112_Y), .CK(T10755_Y));
KC_SDFFRNHQ_X1 T15306 ( .Q(T15306_Q), .SI(T13034_Y), .D(T15306_Q),     .SE(T15498_Y), .RN(T10661_Y), .CK(T10722_Y));
KC_SDFFRNHQ_X1 T15309 ( .Q(T15309_Q), .SI(T12986_Y), .D(T15309_Q),     .SE(T15338_Y), .RN(T837_Y), .CK(T6873_Y));
KC_SDFFRNHQ_X1 T15300 ( .Q(T15300_Q), .SI(T13004_Y), .D(T15300_Q),     .SE(T15414_Y), .RN(T7740_Y), .CK(T7539_Y));
KC_SDFFRNHQ_X1 T15295 ( .Q(T15295_Q), .SI(T12988_Y), .D(T15295_Q),     .SE(T15374_Y), .RN(T5023_Y), .CK(T7128_Y));
KC_SDFFRNHQ_X1 T15293 ( .Q(T15293_Q), .SI(T12990_Y), .D(T15293_Q),     .SE(T15374_Y), .RN(T5023_Y), .CK(T7129_Y));
KC_SDFFRNHQ_X1 T15303 ( .Q(T15303_Q), .SI(T13024_Y), .D(T15303_Q),     .SE(T1051_Y), .RN(T14999_Y), .CK(T7985_Y));
KC_SDFFRNHQ_X1 T15301 ( .Q(T15301_Q), .SI(T13021_Y), .D(T15301_Q),     .SE(T1051_Y), .RN(T14999_Y), .CK(T7925_Y));
KC_SDFFRNHQ_X1 T5595 ( .Q(T5595_Q), .SI(T12994_Y), .D(T5595_Q),     .SE(T15348_Y), .RN(T5023_Y), .CK(T5708_Y));
KC_SDFFRNHQ_X1 T15263 ( .Q(T15263_Q), .SI(T12995_Y), .D(T15263_Q),     .SE(T373_Y), .RN(T5023_Y), .CK(T5743_Y));
KC_SDFFRNHQ_X1 T15269 ( .Q(T15269_Q), .SI(T13041_Y), .D(T15269_Q),     .SE(T15504_Y), .RN(T2522_Y), .CK(T5901_Y));
KC_SDFFRNHQ_X1 T15268 ( .Q(T15268_Q), .SI(T13044_Y), .D(T15268_Q),     .SE(T15504_Y), .RN(T2522_Y), .CK(T5918_Y));
KC_SDFFRNHQ_X1 T15282 ( .Q(T15282_Q), .SI(T13290_Y), .D(T15282_Q),     .SE(T15536_Y), .RN(T2063_Y), .CK(T6705_Y));
KC_SDFFRNHQ_X1 T15273 ( .Q(T15273_Q), .SI(T13095_Y), .D(T15273_Q),     .SE(T15560_Y), .RN(T15009_Y), .CK(T6092_Y));
KC_SDFFRNHQ_X1 T15272 ( .Q(T15272_Q), .SI(T13094_Y), .D(T15272_Q),     .SE(T15560_Y), .RN(T15009_Y), .CK(T6093_Y));
KC_SDFFRNHQ_X1 T15279 ( .Q(T15279_Q), .SI(T13192_Y), .D(T15279_Q),     .SE(T15626_Y), .RN(T837_Y), .CK(T6507_Y));
KC_SDFFRNHQ_X1 T15278 ( .Q(T15278_Q), .SI(T13181_Y), .D(T15278_Q),     .SE(T15626_Y), .RN(T837_Y), .CK(T6508_Y));
KC_SDFFRNHQ_X1 T15265 ( .Q(T15265_Q), .SI(T13206_Y), .D(T15265_Q),     .SE(T16054_Y), .RN(T2522_Y), .CK(T5829_Y));
KC_SDFFRNHQ_X1 T15264 ( .Q(T15264_Q), .SI(T13207_Y), .D(T15264_Q),     .SE(T16109_Y), .RN(T2522_Y), .CK(T5828_Y));
KC_SDFFRNHQ_X1 T15274 ( .Q(T15274_Q), .SI(T13138_Y), .D(T15274_Q),     .SE(T15979_Y), .RN(T837_Y), .CK(T6293_Y));
KC_SDFFRNHQ_X1 T15259 ( .Q(T15259_Q), .SI(T12985_Y), .D(T15259_Q),     .SE(T15364_Y), .RN(T5023_Y), .CK(T5723_Y));
KC_SDFFRNHQ_X1 T15258 ( .Q(T15258_Q), .SI(T12984_Y), .D(T15258_Q),     .SE(T15364_Y), .RN(T5023_Y), .CK(T5716_Y));
KC_SDFFRNHQ_X1 T15261 ( .Q(T15261_Q), .SI(T12991_Y), .D(T15261_Q),     .SE(T15386_Y), .RN(T5023_Y), .CK(T5744_Y));
KC_SDFFRNHQ_X1 T15260 ( .Q(T15260_Q), .SI(T12993_Y), .D(T15260_Q),     .SE(T15386_Y), .RN(T5023_Y), .CK(T6628_Y));
KC_SDFFRNHQ_X1 T15271 ( .Q(T15271_Q), .SI(T13045_Y), .D(T15271_Q),     .SE(T15509_Y), .RN(T4402_Y), .CK(T5931_Y));
KC_SDFFRNHQ_X1 T15270 ( .Q(T15270_Q), .SI(T13043_Y), .D(T15270_Q),     .SE(T15509_Y), .RN(T4402_Y), .CK(T5933_Y));
KC_SDFFRNHQ_X1 T15281 ( .Q(T15281_Q), .SI(T13061_Y), .D(T15281_Q),     .SE(T15536_Y), .RN(T2063_Y), .CK(T6704_Y));
KC_SDFFRNHQ_X1 T15290 ( .Q(T15290_Q), .SI(T12987_Y), .D(T15290_Q),     .SE(T15338_Y), .RN(T837_Y), .CK(T6871_Y));
KC_SDFFRNHQ_X1 T15283 ( .Q(T15283_Q), .SI(T13212_Y), .D(T15283_Q),     .SE(T15325_Y), .RN(T14970_Y), .CK(T5583_Y));
KC_SDFFRNHQ_X1 T15280 ( .Q(T15280_Q), .SI(T12996_Y), .D(T15280_Q),     .SE(T15348_Y), .RN(T5023_Y), .CK(T5709_Y));
KC_SDFFRNHQ_X1 T15294 ( .Q(T15294_Q), .SI(T12989_Y), .D(T15294_Q),     .SE(T15674_Y), .RN(T837_Y), .CK(T7184_Y));
KC_SDFFRNHQ_X1 T15262 ( .Q(T15262_Q), .SI(T12992_Y), .D(T15262_Q),     .SE(T373_Y), .RN(T5023_Y), .CK(T5728_Y));
KC_SDFFRNHQ_X1 T15296 ( .Q(T15296_Q), .SI(T12997_Y), .D(T15296_Q),     .SE(T15674_Y), .RN(T837_Y), .CK(T7353_Y));
KC_SDFFRNHQ_X1 T15308 ( .Q(T15308_Q), .SI(T13204_Y), .D(T15308_Q),     .SE(T15414_Y), .RN(T7740_Y), .CK(T10787_Y));
KC_SDFFRNHQ_X1 T15298 ( .Q(T15298_Q), .SI(T13271_Y), .D(T15298_Q),     .SE(T15409_Y), .RN(T837_Y), .CK(T7408_Y));
KC_SDFFRNHQ_X1 T15297 ( .Q(T15297_Q), .SI(T13234_Y), .D(T15297_Q),     .SE(T15409_Y), .RN(T837_Y), .CK(T7409_Y));
KC_SDFFRNHQ_X1 T15267 ( .Q(T15267_Q), .SI(T13208_Y), .D(T15267_Q),     .SE(T15427_Y), .RN(T2522_Y), .CK(T6675_Y));
KC_SDFFRNHQ_X1 T15266 ( .Q(T15266_Q), .SI(T13005_Y), .D(T15266_Q),     .SE(T15427_Y), .RN(T2522_Y), .CK(T5836_Y));
KC_SDFFRNHQ_X1 T15275 ( .Q(T15275_Q), .SI(T12979_Y), .D(T15275_Q),     .SE(T15595_Y), .RN(T837_Y), .CK(T6271_Y));
KC_SDFFRNHQ_X1 T15277 ( .Q(T15277_Q), .SI(T13147_Y), .D(T15277_Q),     .SE(T15602_Y), .RN(T15035_Y), .CK(T6333_Y));
KC_SDFFRNHQ_X1 T15276 ( .Q(T15276_Q), .SI(T13146_Y), .D(T15276_Q),     .SE(T15602_Y), .RN(T15035_Y), .CK(T6308_Y));
KC_BUF_X9 T14970 ( .Y(T14970_Y), .A(T7668_Y));
KC_BUF_X9 T15024 ( .Y(T15024_Y), .A(T7668_Y));
KC_BUF_X9 T14972 ( .Y(T14972_Y), .A(T135_Q));
KC_BUF_X9 T14976 ( .Y(T14976_Y), .A(T869_Y));
KC_BUF_X9 T14975 ( .Y(T14975_Y), .A(T869_Y));
KC_BUF_X9 T14978 ( .Y(T14978_Y), .A(T869_Y));
KC_BUF_X9 T14974 ( .Y(T14974_Y), .A(T14976_Y));
KC_BUF_X9 T15030 ( .Y(T15030_Y), .A(T7668_Y));
KC_BUF_X9 T14985 ( .Y(T14985_Y), .A(T7668_Y));
KC_BUF_X9 T15031 ( .Y(T15031_Y), .A(T8807_Y));
KC_BUF_X9 T15027 ( .Y(T15027_Y), .A(T7668_Y));
KC_BUF_X9 T14973 ( .Y(T14973_Y), .A(T7668_Y));
KC_BUF_X9 T14979 ( .Y(T14979_Y), .A(T7668_Y));
KC_BUF_X9 T14986 ( .Y(T14986_Y), .A(T15732_Y));
KC_BUF_X9 T15004 ( .Y(T15004_Y), .A(T15004_A));
KC_BUF_X9 T15026 ( .Y(T15026_Y), .A(T7668_Y));
KC_BUF_X9 T14977 ( .Y(T14977_Y), .A(T7668_Y));
KC_BUF_X9 T14991 ( .Y(T14991_Y), .A(T12095_Y));
KC_BUF_X9 T14997 ( .Y(T14997_Y), .A(T1244_Y));
KC_BUF_X9 T14996 ( .Y(T14996_Y), .A(T8030_Y));
KC_BUF_X9 T15001 ( .Y(T15001_Y), .A(T1244_Y));
KC_BUF_X9 T15005 ( .Y(T15005_Y), .A(T9456_Q));
KC_BUF_X9 T14993 ( .Y(T14993_Y), .A(T1244_Y));
KC_BUF_X9 T15002 ( .Y(T15002_Y), .A(T1244_Y));
KC_BUF_X9 T14992 ( .Y(T14992_Y), .A(T15000_Y));
KC_BUF_X9 T14980 ( .Y(T14980_Y), .A(T2027_Y));
KC_BUF_X9 T15000 ( .Y(T15000_Y), .A(T1244_Y));
KC_BUF_X9 T14999 ( .Y(T14999_Y), .A(T1244_Y));
KC_BUF_X9 T14988 ( .Y(T14988_Y), .A(T2000_Y));
KC_BUF_X9 T14987 ( .Y(T14987_Y), .A(T13097_Y));
KC_BUF_X9 T14968 ( .Y(T14968_Y), .A(T1751_Q));
KC_BUF_X9 T14990 ( .Y(T14990_Y), .A(T13113_Y));
KC_BUF_X9 T15003 ( .Y(T15003_Y), .A(T14999_Y));
KC_BUF_X9 T15011 ( .Y(T15011_Y), .A(T2081_Y));
KC_BUF_X9 T15015 ( .Y(T15015_Y), .A(T2081_Y));
KC_BUF_X9 T15021 ( .Y(T15021_Y), .A(T2081_Y));
KC_BUF_X9 T15037 ( .Y(T15037_Y), .A(T2081_Y));
KC_BUF_X9 T14984 ( .Y(T14984_Y), .A(T10263_Y));
KC_BUF_X9 T14989 ( .Y(T14989_Y), .A(T13082_Y));
KC_BUF_X9 T14995 ( .Y(T14995_Y), .A(T16164_Y));
KC_BUF_X9 T15034 ( .Y(T15034_Y), .A(T2709_Y));
KC_BUF_X9 T15008 ( .Y(T15008_Y), .A(T15034_Y));
KC_BUF_X9 T15013 ( .Y(T15013_Y), .A(T2709_Y));
KC_BUF_X9 T15009 ( .Y(T15009_Y), .A(T2709_Y));
KC_BUF_X9 T14994 ( .Y(T14994_Y), .A(T9957_Y));
KC_BUF_X9 T15014 ( .Y(T15014_Y), .A(T4532_Y));
KC_BUF_X9 T15023 ( .Y(T15023_Y), .A(T2709_Y));
KC_BUF_X9 T15016 ( .Y(T15016_Y), .A(T2709_Y));
KC_BUF_X9 T15017 ( .Y(T15017_Y), .A(T5023_Y));
KC_BUF_X9 T15020 ( .Y(T15020_Y), .A(T2081_Y));
KC_BUF_X9 T15033 ( .Y(T15033_Y), .A(T2709_Y));
KC_BUF_X9 T15022 ( .Y(T15022_Y), .A(T15020_Y));
KC_BUF_X9 T15029 ( .Y(T15029_Y), .A(T15721_Y));
KC_BUF_X9 T15028 ( .Y(T15028_Y), .A(T11208_Y));
KC_BUF_X9 T15035 ( .Y(T15035_Y), .A(T2709_Y));
KC_BUF_X9 T15032 ( .Y(T15032_Y), .A(T13300_Y));
KC_BUF_X9 T15018 ( .Y(T15018_Y), .A(T2081_Y));
KC_MX2_X1 T6854 ( .Y(T6854_Y), .A(T25_Y), .S0(T13068_Y), .B(T15330_Y));
KC_MX2_X1 T6853 ( .Y(T6853_Y), .A(T23_Y), .S0(T13068_Y), .B(T15330_Y));
KC_MX2_X1 T5646 ( .Y(T5646_Y), .A(T38_Y), .S0(T13075_Y), .B(T15326_Y));
KC_MX2_X1 T5645 ( .Y(T5645_Y), .A(T5191_Y), .S0(T13075_Y),     .B(T15326_Y));
KC_MX2_X1 T5610 ( .Y(T5610_Y), .A(T64_Y), .S0(T70_Y), .B(T13317_Y));
KC_MX2_X1 T72 ( .Y(T72_Y), .A(T76_Y), .S0(T70_Y), .B(T13317_Y));
KC_MX2_X1 T5621 ( .Y(T5621_Y), .A(T113_Y), .S0(T15321_Y),     .B(T15322_Y));
KC_MX2_X1 T5620 ( .Y(T5620_Y), .A(T5188_Y), .S0(T15321_Y),     .B(T15322_Y));
KC_MX2_X1 T7459 ( .Y(T7459_Y), .A(T195_Y), .S0(T15407_Y), .B(T6832_Y));
KC_MX2_X1 T7433 ( .Y(T7433_Y), .A(T194_Y), .S0(T15407_Y), .B(T6832_Y));
KC_MX2_X1 T7117 ( .Y(T7117_Y), .A(T471_Y), .S0(T15369_Y),     .B(T15370_Y));
KC_MX2_X1 T7116 ( .Y(T7116_Y), .A(T463_Y), .S0(T15369_Y),     .B(T15370_Y));
KC_MX2_X1 T8040 ( .Y(T8040_Y), .A(T581_Y), .S0(T15484_Y),     .B(T15657_Y));
KC_MX2_X1 T8039 ( .Y(T8039_Y), .A(T574_Y), .S0(T15484_Y),     .B(T15657_Y));
KC_MX2_X1 T6858 ( .Y(T6858_Y), .A(T806_Y), .S0(T15335_Y),     .B(T15333_Y));
KC_MX2_X1 T6857 ( .Y(T6857_Y), .A(T805_Y), .S0(T15335_Y),     .B(T15333_Y));
KC_MX2_X1 T7406 ( .Y(T7406_Y), .A(T888_Y), .S0(T15411_Y),     .B(T15410_Y));
KC_MX2_X1 T7390 ( .Y(T7390_Y), .A(T873_Y), .S0(T15411_Y),     .B(T15410_Y));
KC_MX2_X1 T10039 ( .Y(T10039_Y), .A(T1227_Y), .S0(T15496_Y),     .B(T15499_Y));
KC_MX2_X1 T10020 ( .Y(T10020_Y), .A(T1236_Y), .S0(T15496_Y),     .B(T15499_Y));
KC_MX2_X1 T10128 ( .Y(T10128_Y), .A(T15527_Y), .S0(T1738_Y),     .B(T1368_Y));
KC_MX2_X1 T10226 ( .Y(T10226_Y), .A(T1383_Y), .S0(T15544_Y),     .B(T1505_Y));
KC_MX2_X1 T6870 ( .Y(T6870_Y), .A(T1389_Y), .S0(T15342_Y),     .B(T15345_Y));
KC_MX2_X1 T7534 ( .Y(T7534_Y), .A(T1455_Y), .S0(T15415_Y),     .B(T15416_Y));
KC_MX2_X1 T10400 ( .Y(T10400_Y), .A(T1537_Y), .S0(T8671_Y),     .B(T15376_Y));
KC_MX2_X1 T7186 ( .Y(T7186_Y), .A(T1539_Y), .S0(T8671_Y),     .B(T15376_Y));
KC_MX2_X1 T10304 ( .Y(T10304_Y), .A(T1596_Y), .S0(T984_Y),     .B(T15459_Y));
KC_MX2_X1 T7979 ( .Y(T7979_Y), .A(T1564_Y), .S0(T984_Y), .B(T15459_Y));
KC_MX2_X1 T5705 ( .Y(T5705_Y), .A(T1869_Y), .S0(T15347_Y),     .B(T15346_Y));
KC_MX2_X1 T6604 ( .Y(T6604_Y), .A(T2375_Y), .S0(T2365_Y),     .B(T15645_Y));
KC_MX2_X1 T5742 ( .Y(T5742_Y), .A(T2439_Y), .S0(T15381_Y),     .B(T15380_Y));
KC_MX2_X1 T5727 ( .Y(T5727_Y), .A(T3010_Y), .S0(T15381_Y),     .B(T15380_Y));
KC_MX2_X1 T6297 ( .Y(T6297_Y), .A(T6295_Y), .S0(T2791_Y),     .B(T15596_Y));
KC_MX2_X1 T5915 ( .Y(T5915_Y), .A(T3150_Y), .S0(T16303_Y),     .B(T15508_Y));
KC_MX2_X1 T6002 ( .Y(T6002_Y), .A(T5078_Y), .S0(T15551_Y),     .B(T5737_Y));
KC_MX2_X1 T6001 ( .Y(T6001_Y), .A(T3187_Y), .S0(T15551_Y),     .B(T5737_Y));
KC_MX2_X1 T6122 ( .Y(T6122_Y), .A(T3231_Y), .S0(T15565_Y),     .B(T15561_Y));
KC_MX2_X1 T6110 ( .Y(T6110_Y), .A(T3238_Y), .S0(T15565_Y),     .B(T15561_Y));
KC_MX2_X1 T6149 ( .Y(T6149_Y), .A(T15911_Y), .S0(T8215_Y),     .B(T15911_Y));
KC_MX2_X1 T6306 ( .Y(T6306_Y), .A(T16026_Y), .S0(T4352_Y),     .B(T15599_Y));
KC_MX2_X1 T6843 ( .Y(T6843_Y), .A(T3503_Y), .S0(T15639_Y),     .B(T6551_Y));
KC_MX2_X1 T6596 ( .Y(T6596_Y), .A(T3531_Y), .S0(T15639_Y),     .B(T6551_Y));
KC_MX2_X1 T6669 ( .Y(T6669_Y), .A(T3647_Y), .S0(T3290_Y),     .B(T15423_Y));
KC_MX2_X1 T5831 ( .Y(T5831_Y), .A(T5132_Y), .S0(T3290_Y),     .B(T15423_Y));
KC_MX2_X1 T6287 ( .Y(T6287_Y), .A(T3956_Y), .S0(T15594_Y),     .B(T15707_Y));
KC_MX2_X1 T5722 ( .Y(T5722_Y), .A(T4188_Y), .S0(T15366_Y),     .B(T15362_Y));
KC_MX2_X1 T5721 ( .Y(T5721_Y), .A(T10457_Y), .S0(T6438_Y),     .B(T9564_Y));
KC_MX2_X1 T5711 ( .Y(T5711_Y), .A(T4195_Y), .S0(T15366_Y),     .B(T15362_Y));
KC_MX2_X1 T6626 ( .Y(T6626_Y), .A(T4207_Y), .S0(T6455_Y),     .B(T15678_Y));
KC_MX2_X1 T5396 ( .Y(T5396_Y), .A(T4328_Y), .S0(T2724_Y),     .B(T15510_Y));
KC_MX2_X1 T5912 ( .Y(T5912_Y), .A(T4329_Y), .S0(T2724_Y),     .B(T15510_Y));
KC_MX2_X1 T6127 ( .Y(T6127_Y), .A(T4502_Y), .S0(T4479_Y), .B(T4501_Y));
KC_MX2_X1 T6484 ( .Y(T6484_Y), .A(T6151_Y), .S0(T4715_Y), .B(T4071_Y));
KC_MX2_X1 T10405 ( .Y(T10405_Y), .A(T4866_Y), .S0(T15673_Y),     .B(T15672_Y));
KC_MX2_X1 T10336 ( .Y(T10336_Y), .A(T1462_Y), .S0(T15415_Y),     .B(T15416_Y));
KC_MX2_X1 T6687 ( .Y(T6687_Y), .A(T4973_Y), .S0(T12941_Y), .B(T635_Y));
KC_MX2_X1 T6788 ( .Y(T6788_Y), .A(T5118_Y), .S0(T15594_Y),     .B(T15707_Y));
KC_MX2_X1 T6627 ( .Y(T6627_Y), .A(T4225_Y), .S0(T6455_Y),     .B(T15678_Y));
KC_MX2_X1 T6891 ( .Y(T6891_Y), .A(T1396_Y), .S0(T15342_Y),     .B(T15345_Y));
KC_MX2_X1 T5707 ( .Y(T5707_Y), .A(T2408_Y), .S0(T15347_Y),     .B(T15346_Y));
KC_MX2_X1 T7183 ( .Y(T7183_Y), .A(T1180_Y), .S0(T15673_Y),     .B(T15672_Y));
KC_MX2_X1 T6677 ( .Y(T6677_Y), .A(T1960_Y), .S0(T6848_Y),     .B(T15426_Y));
KC_MX2_X1 T5796 ( .Y(T5796_Y), .A(T2498_Y), .S0(T6848_Y),     .B(T15426_Y));
KC_MX2_X1 T5916 ( .Y(T5916_Y), .A(T3151_Y), .S0(T16303_Y),     .B(T15508_Y));
KC_MX2_X1 T10129 ( .Y(T10129_Y), .A(T4825_Y), .S0(T1372_Y),     .B(T1372_Y));
KC_MX2_X1 T6068 ( .Y(T6068_Y), .A(T3830_Y), .S0(T5843_Y), .B(T3230_Y));
KC_MX2_X1 T6307 ( .Y(T6307_Y), .A(T5572_Y), .S0(T4352_Y),     .B(T15599_Y));
KC_NOR2B_X3 T15922 ( .B(T15989_Y), .AN(T1790_Q), .Y(T15922_Y));
KC_NOR2B_X3 T16281 ( .B(T10297_Y), .AN(T9437_Y), .Y(T16281_Y));
KC_NOR2B_X3 T16040 ( .B(T2276_Q), .AN(T5567_Q), .Y(T16040_Y));
KC_ADD_C_B_X1 T15927 ( .B(T1555_Y), .A(T7780_Y), .Y(T15927_Y),     .C(T9782_Y));
KC_ADD_C_B_X1 T16067 ( .B(T1734_Q), .A(T16296_Q), .Y(T16067_Y),     .C(T16297_Q));
KC_ADD_C_B_X1 T16066 ( .B(T1729_Q), .A(T1726_Q), .Y(T16066_Y),     .C(T1730_Q));
KC_ADD_C_B_X1 T16065 ( .B(T1723_Q), .A(T1725_Q), .Y(T16065_Y),     .C(T5374_Q));
KC_ADD_C_B_X1 T15915 ( .B(T15039_Y), .A(T15125_Y), .Y(T15915_Y),     .C(T2718_Y));
KC_ADD_C_B_X1 T16472 ( .B(T15646_Y), .A(T15646_Y), .Y(T16472_Y),     .C(T15645_Y));
KC_ADD_C_B_X1 T15992 ( .B(T5057_Y), .A(T16000_Y), .Y(T15992_Y),     .C(T11544_Y));
KC_ADD_C_B_X1 T16084 ( .B(T2871_Y), .A(T2871_Y), .Y(T16084_Y),     .C(T15624_Y));
KC_ADD_C_B_X1 T15874 ( .B(T5799_Y), .A(T4462_Y), .Y(T15874_Y),     .C(T4426_Y));
KC_ADD_C_B_X1 T16022 ( .B(T8325_Y), .A(T16015_Y), .Y(T16022_Y),     .C(T8325_Y));
KC_ADD_C_B_X1 T16080 ( .B(T16124_Y), .A(T8380_Y), .Y(T16080_Y),     .C(T8382_Y));
KC_NOR2_X3 T12440 ( .Y(T12440_Y), .A(T567_Q), .B(T561_Q));
KC_NOR2_X3 T12417 ( .Y(T12417_Y), .A(T561_Q), .B(T1599_Y));
KC_NOR2_X3 T12416 ( .Y(T12416_Y), .A(T1599_Y), .B(T1352_Y));
KC_NOR2_X3 T12415 ( .Y(T12415_Y), .A(T567_Q), .B(T1352_Y));
KC_NOR2_X3 T12414 ( .Y(T12414_Y), .A(T567_Q), .B(T561_Q));
KC_NOR2_X3 T12413 ( .Y(T12413_Y), .A(T561_Q), .B(T1599_Y));
KC_NOR2_X3 T12412 ( .Y(T12412_Y), .A(T1599_Y), .B(T1352_Y));
KC_NOR2_X3 T12411 ( .Y(T12411_Y), .A(T567_Q), .B(T1352_Y));
KC_NOR2_X3 T12457 ( .Y(T12457_Y), .A(T8073_Y), .B(T560_Y));
KC_NOR2_X3 T15735 ( .Y(T15735_Y), .A(T16352_Y), .B(T7684_Y));
KC_NOR2_X3 T600 ( .Y(T600_Y), .A(T16347_Y), .B(T8774_Y));
KC_NOR2_X3 T6805 ( .Y(T6805_Y), .A(T7685_Y), .B(T7644_Y));
KC_NOR2_X3 T6804 ( .Y(T6804_Y), .A(T7563_Y), .B(T7685_Y));
KC_NOR2_X3 T12409 ( .Y(T12409_Y), .A(T7803_Y), .B(T8774_Y));
KC_NOR2_X3 T12408 ( .Y(T12408_Y), .A(T16349_Y), .B(T8774_Y));
KC_NOR2_X3 T12407 ( .Y(T12407_Y), .A(T16349_Y), .B(T7684_Y));
KC_NOR2_X3 T12406 ( .Y(T12406_Y), .A(T16352_Y), .B(T8774_Y));
KC_NOR2_X3 T12405 ( .Y(T12405_Y), .A(T16347_Y), .B(T7684_Y));
KC_NOR2_X3 T12401 ( .Y(T12401_Y), .A(T7685_Y), .B(T7646_Y));
KC_NOR2_X3 T12399 ( .Y(T12399_Y), .A(T7803_Y), .B(T7684_Y));
KC_NOR2_X3 T12398 ( .Y(T12398_Y), .A(T7685_Y), .B(T7645_Y));
KC_NOR2_X3 T12435 ( .Y(T12435_Y), .A(T16350_Y), .B(T7684_Y));
KC_NOR2_X3 T12429 ( .Y(T12429_Y), .A(T16351_Y), .B(T8774_Y));
KC_NOR2_X3 T12427 ( .Y(T12427_Y), .A(T16350_Y), .B(T8774_Y));
KC_NOR2_X3 T12426 ( .Y(T12426_Y), .A(T16348_Y), .B(T8774_Y));
KC_NOR2_X3 T12425 ( .Y(T12425_Y), .A(T16353_Y), .B(T7684_Y));
KC_NOR2_X3 T12424 ( .Y(T12424_Y), .A(T16353_Y), .B(T8774_Y));
KC_NOR2_X3 T10069 ( .Y(T10069_Y), .A(T16006_Y), .B(T8934_Y));
KC_NOR2_X3 T12073 ( .Y(T12073_Y), .A(T7351_Y), .B(T9632_Y));
KC_NOR2_X3 T12327 ( .Y(T12327_Y), .A(T6748_Y), .B(T10372_Y));
KC_NOR2_X3 T12078 ( .Y(T12078_Y), .A(T7320_Y), .B(T9607_Y));
KC_NOR2_X3 T12077 ( .Y(T12077_Y), .A(T7320_Y), .B(T9614_Y));
KC_NOR2_X3 T12076 ( .Y(T12076_Y), .A(T15392_Y), .B(T9607_Y));
KC_NOR2_X3 T12075 ( .Y(T12075_Y), .A(T15392_Y), .B(T9614_Y));
KC_NOR2_X3 T12074 ( .Y(T12074_Y), .A(T7320_Y), .B(T9610_Y));
KC_NOR2_X3 T12088 ( .Y(T12088_Y), .A(T1054_Y), .B(T9920_Y));
KC_NOR2_X3 T12094 ( .Y(T12094_Y), .A(T1479_Y), .B(T9924_Y));
KC_NOR2_X3 T12325 ( .Y(T12325_Y), .A(T6462_Y), .B(T9613_Y));
KC_NOR2_X3 T12332 ( .Y(T12332_Y), .A(T15904_Y), .B(T2279_Y));
KC_NOR2_X3 T12323 ( .Y(T12323_Y), .A(T15904_Y), .B(T1788_Y));
KC_NOR2_X3 T12112 ( .Y(T12112_Y), .A(T15904_Y), .B(T1786_Y));
KC_NOR2_X3 T5732 ( .Y(T5732_Y), .A(T15904_Y), .B(T16042_Y));
KC_NOR2_X3 T12125 ( .Y(T12125_Y), .A(T15904_Y), .B(T2245_Y));
KC_NOR2_X3 T12122 ( .Y(T12122_Y), .A(T15904_Y), .B(T2247_Y));
KC_NOR2_X3 T12121 ( .Y(T12121_Y), .A(T15904_Y), .B(T2344_Y));
KC_NOR2_X3 T12120 ( .Y(T12120_Y), .A(T15904_Y), .B(T4926_Y));
KC_NOR2_X3 T12113 ( .Y(T12113_Y), .A(T15904_Y), .B(T6005_Y));
KC_NOR2_X3 T12344 ( .Y(T12344_Y), .A(T15904_Y), .B(T6028_Y));
KC_NOR2_X3 T12133 ( .Y(T12133_Y), .A(T15904_Y), .B(T2250_Y));
KC_NOR2_X3 T12166 ( .Y(T12166_Y), .A(T15904_Y), .B(T2280_Y));
KC_NOR2_X3 T12192 ( .Y(T12192_Y), .A(T15989_Y), .B(T16041_Y));
KC_NOR2_X3 T12191 ( .Y(T12191_Y), .A(T15989_Y), .B(T6125_Y));
KC_NOR2_X3 T12190 ( .Y(T12190_Y), .A(T15989_Y), .B(T5927_Y));
KC_NOR2_X3 T12188 ( .Y(T12188_Y), .A(T15989_Y), .B(T1804_Y));
KC_NOR2_X3 T12187 ( .Y(T12187_Y), .A(T15989_Y), .B(T15611_Y));
KC_NOR2_X3 T16305 ( .Y(T16305_Y), .A(T1506_Y), .B(T13048_Q));
KC_NOR2_X3 T12108 ( .Y(T12108_Y), .A(T1532_Y), .B(T2031_Y));
KC_NOR2_X3 T12107 ( .Y(T12107_Y), .A(T16269_Y), .B(T2031_Y));
KC_NOR2_X3 T12106 ( .Y(T12106_Y), .A(T15511_Y), .B(T2031_Y));
KC_NOR2_X3 T12105 ( .Y(T12105_Y), .A(T15519_Y), .B(T2031_Y));
KC_NOR2_X3 T12104 ( .Y(T12104_Y), .A(T1548_Y), .B(T2031_Y));
KC_NOR2_X3 T12103 ( .Y(T12103_Y), .A(T15512_Y), .B(T2031_Y));
KC_NOR2_X3 T12102 ( .Y(T12102_Y), .A(T1533_Y), .B(T2031_Y));
KC_NOR2_X3 T12101 ( .Y(T12101_Y), .A(T1519_Y), .B(T2031_Y));
KC_NOR2_X3 T12270 ( .Y(T12270_Y), .A(T2838_Y), .B(T6208_Y));
KC_NOR2_X3 T12269 ( .Y(T12269_Y), .A(T2838_Y), .B(T2862_Y));
KC_NOR2_X3 T12086 ( .Y(T12086_Y), .A(T883_Y), .B(T2505_Y));
KC_NOR2_X3 T12268 ( .Y(T12268_Y), .A(T3526_Y), .B(T2865_Y));
KC_NOR2_X3 T12065 ( .Y(T12065_Y), .A(T3506_Y), .B(T3513_Y));
KC_NOR2_X3 T12148 ( .Y(T12148_Y), .A(T5101_Y), .B(T3797_Y));
KC_NOR2_X3 T12248 ( .Y(T12248_Y), .A(T6555_Q), .B(T3394_Y));
KC_NOR2_X3 T12317 ( .Y(T12317_Y), .A(T11006_Y), .B(T3510_Y));
KC_NOR2_X3 T12084 ( .Y(T12084_Y), .A(T856_Y), .B(T9829_Y));
KC_NOR2_X3 T12208 ( .Y(T12208_Y), .A(T10939_Y), .B(T10925_Y));
KC_NOR2_X3 T15734 ( .Y(T15734_Y), .A(T16351_Y), .B(T7684_Y));
KC_NOR2_X3 T12331 ( .Y(T12331_Y), .A(T15904_Y), .B(T2246_Y));
KC_NOR2_X3 T12324 ( .Y(T12324_Y), .A(T7334_Y), .B(T9612_Y));
KC_NOR2_X3 T16270 ( .Y(T16270_Y), .A(T1517_Y), .B(T2031_Y));
KC_NOR2_X3 T12423 ( .Y(T12423_Y), .A(T16348_Y), .B(T7684_Y));
KC_NOR2_X3 T12329 ( .Y(T12329_Y), .A(T3712_Y), .B(T10505_Y));
KC_NOR2_X3 T12263 ( .Y(T12263_Y), .A(T10617_Y), .B(T3443_Y));
KC_XNOR2_X2 T9430 ( .Y(T9430_Y), .A(T8925_Y), .B(T8826_Y));
KC_XNOR2_X2 T9428 ( .Y(T9428_Y), .A(T8958_Y), .B(T8879_Y));
KC_XNOR2_X2 T9427 ( .Y(T9427_Y), .A(T8922_Y), .B(T7865_Y));
KC_XNOR2_X2 T9426 ( .Y(T9426_Y), .A(T10031_Y), .B(T7874_Y));
KC_XNOR2_X2 T8885 ( .Y(T8885_Y), .A(T8886_Y), .B(T8788_Y));
KC_XNOR2_X2 T8876 ( .Y(T8876_Y), .A(T15082_Y), .B(T8883_Y));
KC_XNOR2_X2 T8875 ( .Y(T8875_Y), .A(T15147_Y), .B(T8090_Y));
KC_XNOR2_X2 T8839 ( .Y(T8839_Y), .A(T15060_Y), .B(T8841_Y));
KC_XNOR2_X2 T8822 ( .Y(T8822_Y), .A(T9490_Y), .B(T2277_Y));
KC_XNOR2_X2 T8820 ( .Y(T8820_Y), .A(T15058_Y), .B(T8929_Y));
KC_XNOR2_X2 T8819 ( .Y(T8819_Y), .A(T15083_Y), .B(T7864_Y));
KC_XNOR2_X2 T8818 ( .Y(T8818_Y), .A(T15079_Y), .B(T7864_Y));
KC_XNOR2_X2 T8817 ( .Y(T8817_Y), .A(T15057_Y), .B(T8823_Y));
KC_XNOR2_X2 T8816 ( .Y(T8816_Y), .A(T8787_Y), .B(T8843_Y));
KC_XNOR2_X2 T8961 ( .Y(T8961_Y), .A(T232_Y), .B(T8959_Y));
KC_XNOR2_X2 T8955 ( .Y(T8955_Y), .A(T8966_Y), .B(T8967_Y));
KC_XNOR2_X2 T8954 ( .Y(T8954_Y), .A(T8970_Y), .B(T8056_Y));
KC_XNOR2_X2 T8953 ( .Y(T8953_Y), .A(T15075_Y), .B(T8089_Y));
KC_XNOR2_X2 T8952 ( .Y(T8952_Y), .A(T8091_Y), .B(T8056_Y));
KC_XNOR2_X2 T8931 ( .Y(T8931_Y), .A(T15144_Y), .B(T8924_Y));
KC_XNOR2_X2 T8930 ( .Y(T8930_Y), .A(T8956_Y), .B(T8089_Y));
KC_XNOR2_X2 T8921 ( .Y(T8921_Y), .A(T15077_Y), .B(T2312_Y));
KC_XNOR2_X2 T8920 ( .Y(T8920_Y), .A(T15078_Y), .B(T232_Y));
KC_XNOR2_X2 T9177 ( .Y(T9177_Y), .A(T1167_Y), .B(T620_Y));
KC_XNOR2_X2 T9176 ( .Y(T9176_Y), .A(T9238_Y), .B(T9499_Y));
KC_XNOR2_X2 T9175 ( .Y(T9175_Y), .A(T15114_Y), .B(T1252_Y));
KC_XNOR2_X2 T9155 ( .Y(T9155_Y), .A(T9179_Y), .B(T9212_Y));
KC_XNOR2_X2 T9154 ( .Y(T9154_Y), .A(T1523_Y), .B(T9179_Y));
KC_XNOR2_X2 T9153 ( .Y(T9153_Y), .A(T15099_Y), .B(T9183_Y));
KC_XNOR2_X2 T9131 ( .Y(T9131_Y), .A(T15094_Y), .B(T2049_Y));
KC_XNOR2_X2 T9130 ( .Y(T9130_Y), .A(T15096_Y), .B(T9139_Y));
KC_XNOR2_X2 T9081 ( .Y(T9081_Y), .A(T9451_Y), .B(T1538_Y));
KC_XNOR2_X2 T9247 ( .Y(T9247_Y), .A(T15119_Y), .B(T9495_Y));
KC_XNOR2_X2 T9245 ( .Y(T9245_Y), .A(T1252_Y), .B(T9213_Y));
KC_XNOR2_X2 T9235 ( .Y(T9235_Y), .A(T9209_Y), .B(T9238_Y));
KC_XNOR2_X2 T9233 ( .Y(T9233_Y), .A(T15111_Y), .B(T15117_Y));
KC_XNOR2_X2 T9232 ( .Y(T9232_Y), .A(T9211_Y), .B(T9208_Y));
KC_XNOR2_X2 T9231 ( .Y(T9231_Y), .A(T15108_Y), .B(T15115_Y));
KC_XNOR2_X2 T8821 ( .Y(T8821_Y), .A(T8825_Y), .B(T88_Y));
KC_XNOR2_X2 T9480 ( .Y(T9480_Y), .A(T15148_Y), .B(T9483_Y));
KC_XNOR2_X2 T9479 ( .Y(T9479_Y), .A(T15116_Y), .B(T620_Y));
KC_XNOR2_X2 T9167 ( .Y(T9167_Y), .A(T654_Y), .B(T9249_Y));
KC_XNOR2_X2 T9244 ( .Y(T9244_Y), .A(T15151_Y), .B(T608_Y));
KC_XNOR2_X2 T9230 ( .Y(T9230_Y), .A(T15106_Y), .B(T9497_Y));
KC_XNOR2_X2 T9229 ( .Y(T9229_Y), .A(T15105_Y), .B(T16516_Y));
KC_XNOR2_X2 T9228 ( .Y(T9228_Y), .A(T426_Y), .B(T16516_Y));
KC_XNOR2_X2 T9196 ( .Y(T9196_Y), .A(T15107_Y), .B(T15149_Y));
KC_XNOR2_X2 T9195 ( .Y(T9195_Y), .A(T9218_Y), .B(T9202_Y));
KC_XNOR2_X2 T9192 ( .Y(T9192_Y), .A(T605_Q), .B(T15860_Q));
KC_XNOR2_X2 T9190 ( .Y(T9190_Y), .A(T567_Q), .B(T15879_Q));
KC_XNOR2_X2 T9189 ( .Y(T9189_Y), .A(T605_Q), .B(T15860_Q));
KC_XNOR2_X2 T9191 ( .Y(T9191_Y), .A(T567_Q), .B(T15879_Q));
KC_XNOR2_X2 T10229 ( .Y(T10229_Y), .A(T15891_Q), .B(T15879_Q));
KC_XNOR2_X2 T9975 ( .Y(T9975_Y), .A(T10529_Y), .B(T9977_Y));
KC_XNOR2_X2 T9942 ( .Y(T9942_Y), .A(T15168_Q), .B(T2021_Y));
KC_XNOR2_X2 T9901 ( .Y(T9901_Y), .A(T15067_Y), .B(T1059_Y));
KC_XNOR2_X2 T10030 ( .Y(T10030_Y), .A(T4412_Y), .B(T1472_Y));
KC_XNOR2_X2 T10029 ( .Y(T10029_Y), .A(T15086_Y), .B(T1456_Y));
KC_XNOR2_X2 T9842 ( .Y(T9842_Y), .A(T15053_Y), .B(T1981_Q));
KC_XNOR2_X2 T9841 ( .Y(T9841_Y), .A(T1970_Q), .B(T13009_Q));
KC_XNOR2_X2 T9840 ( .Y(T9840_Y), .A(T15051_Y), .B(T13017_Q));
KC_XNOR2_X2 T10081 ( .Y(T10081_Y), .A(T10092_Y), .B(T10086_Y));
KC_XNOR2_X2 T8191 ( .Y(T8191_Y), .A(T3339_Y), .B(T2105_Y));
KC_XNOR2_X2 T8210 ( .Y(T8210_Y), .A(T2148_Y), .B(T2106_Y));
KC_XNOR2_X2 T8483 ( .Y(T8483_Y), .A(T2244_Y), .B(T16008_Y));
KC_XNOR2_X2 T8419 ( .Y(T8419_Y), .A(T8410_Y), .B(T2331_Y));
KC_XNOR2_X2 T8158 ( .Y(T8158_Y), .A(T12879_Y), .B(T2393_Y));
KC_XNOR2_X2 T9872 ( .Y(T9872_Y), .A(T9873_Y), .B(T2529_Y));
KC_XNOR2_X2 T9835 ( .Y(T9835_Y), .A(T14093_Q), .B(T2557_Y));
KC_XNOR2_X2 T10514 ( .Y(T10514_Y), .A(T3093_Y), .B(T14893_Q));
KC_XNOR2_X2 T10119 ( .Y(T10119_Y), .A(T16262_Y), .B(T11176_Y));
KC_XNOR2_X2 T10054 ( .Y(T10054_Y), .A(T2614_Y), .B(T11946_Y));
KC_XNOR2_X2 T8214 ( .Y(T8214_Y), .A(T6149_Y), .B(T3249_Y));
KC_XNOR2_X2 T8479 ( .Y(T8479_Y), .A(T3324_Y), .B(T3333_Y));
KC_XNOR2_X2 T8292 ( .Y(T8292_Y), .A(T3321_Y), .B(T8487_Y));
KC_XNOR2_X2 T8336 ( .Y(T8336_Y), .A(T16014_Y), .B(T5478_Y));
KC_XNOR2_X2 T8314 ( .Y(T8314_Y), .A(T8325_Y), .B(T15607_Y));
KC_XNOR2_X2 T9871 ( .Y(T9871_Y), .A(T9861_Y), .B(T6429_Y));
KC_XNOR2_X2 T8221 ( .Y(T8221_Y), .A(T3922_Y), .B(T3886_Y));
KC_XNOR2_X2 T8212 ( .Y(T8212_Y), .A(T2077_Y), .B(T11444_Y));
KC_XNOR2_X2 T8245 ( .Y(T8245_Y), .A(T3934_Y), .B(T5937_Y));
KC_XNOR2_X2 T8476 ( .Y(T8476_Y), .A(T8265_Y), .B(T13119_Q));
KC_XNOR2_X2 T8439 ( .Y(T8439_Y), .A(T15158_Y), .B(T15824_Y));
KC_XNOR2_X2 T8438 ( .Y(T8438_Y), .A(T6031_S), .B(T5746_Y));
KC_XNOR2_X2 T8177 ( .Y(T8177_Y), .A(T12786_Y), .B(T15823_Y));
KC_XNOR2_X2 T8299 ( .Y(T8299_Y), .A(T4623_Y), .B(T4638_Y));
KC_XNOR2_X2 T8365 ( .Y(T8365_Y), .A(T4641_Y), .B(T8370_Y));
KC_XNOR2_X2 T9481 ( .Y(T9481_Y), .A(T9217_Y), .B(T9238_Y));
KC_XNOR2_X2 T10321 ( .Y(T10321_Y), .A(T10322_Y), .B(T11172_Y));
KC_XNOR2_X2 T10511 ( .Y(T10511_Y), .A(T16095_Y), .B(T9843_Y));
KC_XNOR2_X2 T10510 ( .Y(T10510_Y), .A(T4983_Y), .B(T15052_Y));
KC_XNOR2_X2 T8454 ( .Y(T8454_Y), .A(T2689_Q), .B(T5574_Q));
KC_XNOR2_X2 T8169 ( .Y(T8169_Y), .A(T12070_Y), .B(T6545_Y));
KC_XNOR2_X2 T8168 ( .Y(T8168_Y), .A(T6546_Y), .B(T15042_Y));
KC_XNOR2_X2 T8443 ( .Y(T8443_Y), .A(T15163_Y), .B(T15831_Y));
KC_XNOR2_X2 T8449 ( .Y(T8449_Y), .A(T5799_Y), .B(T4462_Y));
KC_XNOR2_X2 T8437 ( .Y(T8437_Y), .A(T15555_Y), .B(T15553_Y));
KC_XNOR2_X2 T8615 ( .Y(T8615_Y), .A(T832_Y), .B(T12390_Y));
KC_XNOR2_X2 T9881 ( .Y(T9881_Y), .A(T4419_Y), .B(T975_Y));
KC_XNOR2_X2 T9429 ( .Y(T9429_Y), .A(T15145_Y), .B(T15080_Y));
KC_XNOR2_X2 T8919 ( .Y(T8919_Y), .A(T8055_Y), .B(T8928_Y));
KC_XNOR2_X2 T8918 ( .Y(T8918_Y), .A(T15076_Y), .B(T8927_Y));
KC_XNOR2_X2 T9473 ( .Y(T9473_Y), .A(T9198_Y), .B(T9206_Y));
KC_XNOR2_X2 T9246 ( .Y(T9246_Y), .A(T15112_Y), .B(T608_Y));
KC_XNOR2_X2 T9234 ( .Y(T9234_Y), .A(T9237_Y), .B(T9210_Y));
KC_XNOR2_X2 T9200 ( .Y(T9200_Y), .A(T15113_Y), .B(T9498_Y));
KC_XNOR2_X2 T8231 ( .Y(T8231_Y), .A(T15857_Y), .B(T3266_Y));
KC_XNOR2_X2 T8383 ( .Y(T8383_Y), .A(T16080_Y), .B(T10603_Y));
KC_BUF_X4 T16477 ( .Y(T16477_Y), .A(T13332_Q));
KC_BUF_X4 T16476 ( .Y(T16476_Y), .A(T991_Y));
KC_BUF_X4 T15175 ( .Y(T15175_Y), .A(T991_Y));
KC_BUF_X4 T837 ( .Y(T837_Y), .A(T7668_Y));
KC_BUF_X4 T15173 ( .Y(T15173_Y), .A(T991_Y));
KC_BUF_X4 T15185 ( .Y(T15185_Y), .A(T991_Y));
KC_BUF_X4 T15184 ( .Y(T15184_Y), .A(T15183_Q));
KC_BUF_X4 T15180 ( .Y(T15180_Y), .A(T13064_Q));
KC_BUF_X4 T15167 ( .Y(T15167_Y), .A(T15167_A));
KC_BUF_X4 T15190 ( .Y(T15190_Y), .A(T15190_A));
KC_BUF_X4 T15176 ( .Y(T15176_Y), .A(T1515_Y));
KC_BUF_X4 T15188 ( .Y(T15188_Y), .A(T1374_Y));
KC_BUF_X4 T16475 ( .Y(T16475_Y), .A(T1855_Y));
KC_BUF_X4 T1851 ( .Y(T1851_Y), .A(T2401_Y));
KC_BUF_X4 T1852 ( .Y(T1852_Y), .A(T15957_Y));
KC_BUF_X4 T1853 ( .Y(T1853_Y), .A(T8420_Y));
KC_BUF_X4 T1854 ( .Y(T1854_Y), .A(T5547_Y));
KC_BUF_X4 T15174 ( .Y(T15174_Y), .A(T14964_Y));
KC_BUF_X4 T2125 ( .Y(T2125_Y), .A(T2128_Q));
KC_BUF_X4 T15187 ( .Y(T15187_Y), .A(T15180_Y));
KC_BUF_X4 T15186 ( .Y(T15186_Y), .A(T14545_Q));
KC_BUF_X4 T15192 ( .Y(T15192_Y), .A(T16134_Y));
KC_BUF_X4 T5023 ( .Y(T5023_Y), .A(T15230_Y));
KC_BUF_X4 T15172 ( .Y(T15172_Y), .A(T991_Y));
KC_BUF_X4 T5508 ( .Y(T5508_Y), .A(T2309_Y));
KC_NAND3_X1 T8560 ( .Y(T8560_Y), .B(T5203_Q), .C(T8559_Y), .A(T107_Q));
KC_NAND3_X1 T8554 ( .Y(T8554_Y), .B(T107_Q), .C(T5202_Q), .A(T8553_Y));
KC_NAND3_X1 T8542 ( .Y(T8542_Y), .B(T8545_Y), .C(T16479_Y),     .A(T8543_Y));
KC_NAND3_X1 T8541 ( .Y(T8541_Y), .B(T8546_Y), .C(T16310_Y),     .A(T1201_Y));
KC_NAND3_X1 T8540 ( .Y(T8540_Y), .B(T15318_Y), .C(T5614_Y),     .A(T12368_Y));
KC_NAND3_X1 T8539 ( .Y(T8539_Y), .B(T12470_Y), .C(T5616_Y),     .A(T878_Y));
KC_NAND3_X1 T8603 ( .Y(T8603_Y), .B(T8601_Y), .C(T236_Y), .A(T5222_Q));
KC_NAND3_X1 T8582 ( .Y(T8582_Y), .B(T255_Y), .C(T257_Y), .A(T8579_Y));
KC_NAND3_X1 T8581 ( .Y(T8581_Y), .B(T133_Q), .C(T15358_Y), .A(T150_Q));
KC_NAND3_X1 T8568 ( .Y(T8568_Y), .B(T878_Y), .C(T12475_Y), .A(T228_Y));
KC_NAND3_X1 T8628 ( .Y(T8628_Y), .B(T8746_Y), .C(T7845_Y),     .A(T7122_Y));
KC_NAND3_X1 T8747 ( .Y(T8747_Y), .B(T15765_Y), .C(T15430_Y),     .A(T208_Q));
KC_NAND3_X1 T8746 ( .Y(T8746_Y), .B(T215_Q), .C(T650_Y), .A(T15769_Y));
KC_NAND3_X1 T9029 ( .Y(T9029_Y), .B(T16289_Y), .C(T1430_Y),     .A(T9086_Y));
KC_NAND3_X1 T9157 ( .Y(T9157_Y), .B(T4800_Y), .C(T15118_Y),     .A(T15100_Y));
KC_NAND3_X1 T9156 ( .Y(T9156_Y), .B(T15100_Y), .C(T4800_Y),     .A(T4818_Y));
KC_NAND3_X1 T8704 ( .Y(T8704_Y), .B(T16323_Y), .C(T16312_Y),     .A(T7694_Y));
KC_NAND3_X1 T8703 ( .Y(T8703_Y), .B(T7692_Y), .C(T16322_Y),     .A(T7691_Y));
KC_NAND3_X1 T8874 ( .Y(T8874_Y), .B(T8950_Y), .C(T9066_Y),     .A(T8865_Y));
KC_NAND3_X1 T8815 ( .Y(T8815_Y), .B(T9259_Y), .C(T9110_Y), .A(T371_Y));
KC_NAND3_X1 T8785 ( .Y(T8785_Y), .B(T9381_Y), .C(T9149_Y),     .A(T8777_Y));
KC_NAND3_X1 T9023 ( .Y(T9023_Y), .B(T1438_Y), .C(T16286_Y),     .A(T1429_Y));
KC_NAND3_X1 T9022 ( .Y(T9022_Y), .B(T1438_Y), .C(T16286_Y),     .A(T1439_Y));
KC_NAND3_X1 T8988 ( .Y(T8988_Y), .B(T1440_Y), .C(T16286_Y),     .A(T1439_Y));
KC_NAND3_X1 T8987 ( .Y(T8987_Y), .B(T1440_Y), .C(T16286_Y),     .A(T1429_Y));
KC_NAND3_X1 T8986 ( .Y(T8986_Y), .B(T1440_Y), .C(T16286_Y),     .A(T9071_Y));
KC_NAND3_X1 T8985 ( .Y(T8985_Y), .B(T1438_Y), .C(T16286_Y),     .A(T9071_Y));
KC_NAND3_X1 T8984 ( .Y(T8984_Y), .B(T1594_Y), .C(T8779_Y),     .A(T5354_Q));
KC_NAND3_X1 T8951 ( .Y(T8951_Y), .B(T8085_Y), .C(T15794_Y),     .A(T8054_Y));
KC_NAND3_X1 T8917 ( .Y(T8917_Y), .B(T8047_Y), .C(T8084_Y),     .A(T8074_Y));
KC_NAND3_X1 T8907 ( .Y(T8907_Y), .B(T16361_Y), .C(T15793_Y),     .A(T8051_Y));
KC_NAND3_X1 T9076 ( .Y(T9076_Y), .B(T9119_Y), .C(T9447_Y),     .A(T9072_Y));
KC_NAND3_X1 T9075 ( .Y(T9075_Y), .B(T9069_Y), .C(T9447_Y),     .A(T9119_Y));
KC_NAND3_X1 T9074 ( .Y(T9074_Y), .B(T9123_Y), .C(T9447_Y),     .A(T9120_Y));
KC_NAND3_X1 T8573 ( .Y(T8573_Y), .B(T8852_Y), .C(T6247_Y), .A(T311_Y));
KC_NAND3_X1 T8624 ( .Y(T8624_Y), .B(T8894_Y), .C(T1096_Y),     .A(T6348_Y));
KC_NAND3_X1 T9514 ( .Y(T9514_Y), .B(T8895_Y), .C(T6601_Y),     .A(T6613_Y));
KC_NAND3_X1 T8653 ( .Y(T8653_Y), .B(T7252_Y), .C(T7301_Y),     .A(T8652_Y));
KC_NAND3_X1 T8645 ( .Y(T8645_Y), .B(T7270_Y), .C(T7265_Y),     .A(T8644_Y));
KC_NAND3_X1 T8642 ( .Y(T8642_Y), .B(T7100_Y), .C(T6349_Y),     .A(T9258_Y));
KC_NAND3_X1 T9348 ( .Y(T9348_Y), .B(T9411_Y), .C(T15726_Y),     .A(T6671_Y));
KC_NAND3_X1 T9347 ( .Y(T9347_Y), .B(T6664_Y), .C(T7447_Y),     .A(T9345_Y));
KC_NAND3_X1 T9324 ( .Y(T9324_Y), .B(T5252_Q), .C(T6808_Y), .A(T905_Y));
KC_NAND3_X1 T9323 ( .Y(T9323_Y), .B(T6606_Y), .C(T6710_Y),     .A(T8668_Y));
KC_NAND3_X1 T8681 ( .Y(T8681_Y), .B(T7377_Y), .C(T7445_Y),     .A(T8680_Y));
KC_NAND3_X1 T8674 ( .Y(T8674_Y), .B(T7401_Y), .C(T7370_Y),     .A(T8672_Y));
KC_NAND3_X1 T8664 ( .Y(T8664_Y), .B(T6397_Y), .C(T535_Y), .A(T562_Y));
KC_NAND3_X1 T8750 ( .Y(T8750_Y), .B(T512_Q), .C(T916_Y), .A(T5357_Q));
KC_NAND3_X1 T8712 ( .Y(T8712_Y), .B(T9001_Y), .C(T15727_Y),     .A(T6662_Y));
KC_NAND3_X1 T8947 ( .Y(T8947_Y), .B(T1350_Y), .C(T1328_Y),     .A(T5377_Q));
KC_NAND3_X1 T8946 ( .Y(T8946_Y), .B(T16311_Y), .C(T1323_Y),     .A(T8977_Y));
KC_NAND3_X1 T8909 ( .Y(T8909_Y), .B(T8059_Y), .C(T16310_Y),     .A(T1201_Y));
KC_NAND3_X1 T8908 ( .Y(T8908_Y), .B(T1201_Y), .C(T8059_Y),     .A(T1205_Y));
KC_NAND3_X1 T9166 ( .Y(T9166_Y), .B(T9469_Q), .C(T9164_Y),     .A(T5406_Q));
KC_NAND3_X1 T9160 ( .Y(T9160_Y), .B(T8123_Y), .C(T9107_Y),     .A(T5406_Q));
KC_NAND3_X1 T9111 ( .Y(T9111_Y), .B(T9469_Q), .C(T9145_Y),     .A(T5406_Q));
KC_NAND3_X1 T9110 ( .Y(T9110_Y), .B(T9469_Q), .C(T9144_Y),     .A(T5406_Q));
KC_NAND3_X1 T8622 ( .Y(T8622_Y), .B(T9408_Y), .C(T6248_Y),     .A(T6332_Y));
KC_NAND3_X1 T8621 ( .Y(T8621_Y), .B(T9409_Y), .C(T6249_Y), .A(T333_Y));
KC_NAND3_X1 T8620 ( .Y(T8620_Y), .B(T8802_Y), .C(T6246_Y), .A(T339_Y));
KC_NAND3_X1 T8643 ( .Y(T8643_Y), .B(T12526_Y), .C(T675_Y),     .A(T6485_Y));
KC_NAND3_X1 T8721 ( .Y(T8721_Y), .B(T8854_Y), .C(T15766_Y),     .A(T737_Y));
KC_NAND3_X1 T8693 ( .Y(T8693_Y), .B(T701_Q), .C(T932_Y), .A(T724_Q));
KC_NAND3_X1 T8688 ( .Y(T8688_Y), .B(T8767_Y), .C(T7646_Y),     .A(T8831_Y));
KC_NAND3_X1 T15842 ( .Y(T15842_Y), .B(T8946_Y), .C(T16388_Y),     .A(T758_Y));
KC_NAND3_X1 T8773 ( .Y(T8773_Y), .B(T8767_Y), .C(T7563_Y), .A(T786_Y));
KC_NAND3_X1 T9006 ( .Y(T9006_Y), .B(T9028_Y), .C(T972_Y), .A(T9440_Y));
KC_NAND3_X1 T8905 ( .Y(T8905_Y), .B(T8064_Y), .C(T8117_Y),     .A(T16420_Y));
KC_NAND3_X1 T8904 ( .Y(T8904_Y), .B(T8117_Y), .C(T8038_Y),     .A(T8072_Y));
KC_NAND3_X1 T9278 ( .Y(T9278_Y), .B(T6919_Y), .C(T6290_Y), .A(T822_Q));
KC_NAND3_X1 T8619 ( .Y(T8619_Y), .B(T8893_Y), .C(T6252_Y), .A(T334_Y));
KC_NAND3_X1 T8641 ( .Y(T8641_Y), .B(T9410_Y), .C(T6480_Y),     .A(T15647_Y));
KC_NAND3_X1 T9328 ( .Y(T9328_Y), .B(T8676_Y), .C(T11877_Y),     .A(T8732_Y));
KC_NAND3_X1 T9305 ( .Y(T9305_Y), .B(T6694_Y), .C(T9373_Y),     .A(T8670_Y));
KC_NAND3_X1 T9304 ( .Y(T9304_Y), .B(T6694_Y), .C(T9374_Y),     .A(T8670_Y));
KC_NAND3_X1 T8676 ( .Y(T8676_Y), .B(T9340_Q), .C(T10345_Y),     .A(T6825_Y));
KC_NAND3_X1 T8732 ( .Y(T8732_Y), .B(T8728_Y), .C(T15454_Y),     .A(T15431_Y));
KC_NAND3_X1 T8731 ( .Y(T8731_Y), .B(T8729_Y), .C(T11180_Y),     .A(T8732_Y));
KC_NAND3_X1 T8730 ( .Y(T8730_Y), .B(T5300_Q), .C(T639_Y), .A(T6825_Y));
KC_NAND3_X1 T8729 ( .Y(T8729_Y), .B(T6825_Y), .C(T7635_Y), .A(T711_Q));
KC_NAND3_X1 T8709 ( .Y(T8709_Y), .B(T8708_Y), .C(T11195_Y),     .A(T8732_Y));
KC_NAND3_X1 T8708 ( .Y(T8708_Y), .B(T710_Q), .C(T15428_Y),     .A(T6825_Y));
KC_NAND3_X1 T8687 ( .Y(T8687_Y), .B(T8730_Y), .C(T11179_Y),     .A(T8732_Y));
KC_NAND3_X1 T9414 ( .Y(T9414_Y), .B(T129_Y), .C(T7876_Y),     .A(T16386_Y));
KC_NAND3_X1 T8849 ( .Y(T8849_Y), .B(T938_Q), .C(T8845_Y), .A(T925_Y));
KC_NAND3_X1 T8800 ( .Y(T8800_Y), .B(T8791_Y), .C(T15458_Y),     .A(T949_Q));
KC_NAND3_X1 T8799 ( .Y(T8799_Y), .B(T938_Q), .C(T8796_Y), .A(T940_Q));
KC_NAND3_X1 T8892 ( .Y(T8892_Y), .B(T12884_Y), .C(T7835_Y),     .A(T1196_Y));
KC_NAND3_X1 T9187 ( .Y(T9187_Y), .B(T9222_Y), .C(T9186_Y),     .A(T9184_Y));
KC_NAND3_X1 T8677 ( .Y(T8677_Y), .B(T8678_Y), .C(T11875_Y),     .A(T8732_Y));
KC_NAND3_X1 T8659 ( .Y(T8659_Y), .B(T8658_Y), .C(T11876_Y),     .A(T8732_Y));
KC_NAND3_X1 T9404 ( .Y(T9404_Y), .B(T8032_Y), .C(T16384_Y),     .A(T980_Q));
KC_NAND3_X1 T8850 ( .Y(T8850_Y), .B(T7840_Y), .C(T9404_Y),     .A(T1095_Q));
KC_NAND3_X1 T8798 ( .Y(T8798_Y), .B(T980_Q), .C(T946_Y), .A(T1131_Q));
KC_NAND3_X1 T10007 ( .Y(T10007_Y), .B(T1130_Q), .C(T1131_Q),     .A(T980_Q));
KC_NAND3_X1 T8938 ( .Y(T8938_Y), .B(T8032_Y), .C(T8935_Y),     .A(T1469_Y));
KC_NAND3_X1 T9983 ( .Y(T9983_Y), .B(T1362_Y), .C(T10155_Y),     .A(T1366_Y));
KC_NAND3_X1 T10172 ( .Y(T10172_Y), .B(T12093_Y), .C(T9986_Y),     .A(T10162_Y));
KC_NAND3_X1 T10403 ( .Y(T10403_Y), .B(T3072_Y), .C(T361_Y),     .A(T3071_Y));
KC_NAND3_X1 T9582 ( .Y(T9582_Y), .B(T361_Y), .C(T1633_Y), .A(T3071_Y));
KC_NAND3_X1 T9581 ( .Y(T9581_Y), .B(T361_Y), .C(T6595_Y), .A(T3072_Y));
KC_NAND3_X1 T10428 ( .Y(T10428_Y), .B(T6747_Y), .C(T6595_Y),     .A(T3072_Y));
KC_NAND3_X1 T10427 ( .Y(T10427_Y), .B(T6747_Y), .C(T1633_Y),     .A(T3071_Y));
KC_NAND3_X1 T10426 ( .Y(T10426_Y), .B(T3072_Y), .C(T6747_Y),     .A(T3071_Y));
KC_NAND3_X1 T10424 ( .Y(T10424_Y), .B(T403_Y), .C(T6839_Y),     .A(T3650_Y));
KC_NAND3_X1 T9633 ( .Y(T9633_Y), .B(T3650_Y), .C(T403_Y), .A(T3653_Y));
KC_NAND3_X1 T9632 ( .Y(T9632_Y), .B(T403_Y), .C(T6839_Y), .A(T3650_Y));
KC_NAND3_X1 T9631 ( .Y(T9631_Y), .B(T403_Y), .C(T6802_Y), .A(T3653_Y));
KC_NAND3_X1 T9543 ( .Y(T9543_Y), .B(T12081_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T9542 ( .Y(T9542_Y), .B(T12081_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T9541 ( .Y(T9541_Y), .B(T12083_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T9540 ( .Y(T9540_Y), .B(T12083_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T9721 ( .Y(T9721_Y), .B(T2534_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T9720 ( .Y(T9720_Y), .B(T2534_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T9810 ( .Y(T9810_Y), .B(T12328_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T10015 ( .Y(T10015_Y), .B(T9889_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T10014 ( .Y(T10014_Y), .B(T9889_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T10415 ( .Y(T10415_Y), .B(T403_Y), .C(T6802_Y),     .A(T3653_Y));
KC_NAND3_X1 T10414 ( .Y(T10414_Y), .B(T403_Y), .C(T6839_Y),     .A(T3650_Y));
KC_NAND3_X1 T10411 ( .Y(T10411_Y), .B(T2451_Y), .C(T1633_Y),     .A(T3071_Y));
KC_NAND3_X1 T10410 ( .Y(T10410_Y), .B(T2451_Y), .C(T6595_Y),     .A(T3072_Y));
KC_NAND3_X1 T9614 ( .Y(T9614_Y), .B(T403_Y), .C(T6802_Y), .A(T3653_Y));
KC_NAND3_X1 T9610 ( .Y(T9610_Y), .B(T403_Y), .C(T6839_Y), .A(T3650_Y));
KC_NAND3_X1 T9607 ( .Y(T9607_Y), .B(T3650_Y), .C(T403_Y), .A(T3653_Y));
KC_NAND3_X1 T10356 ( .Y(T10356_Y), .B(T3650_Y), .C(T403_Y),     .A(T3653_Y));
KC_NAND3_X1 T9787 ( .Y(T9787_Y), .B(T12328_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T10319 ( .Y(T10319_Y), .B(T3650_Y), .C(T16397_Y),     .A(T3653_Y));
KC_NAND3_X1 T9924 ( .Y(T9924_Y), .B(T3683_Y), .C(T1633_Y),     .A(T3071_Y));
KC_NAND3_X1 T9922 ( .Y(T9922_Y), .B(T3683_Y), .C(T6595_Y),     .A(T3072_Y));
KC_NAND3_X1 T9921 ( .Y(T9921_Y), .B(T16397_Y), .C(T6839_Y),     .A(T3650_Y));
KC_NAND3_X1 T9920 ( .Y(T9920_Y), .B(T16397_Y), .C(T6802_Y),     .A(T3653_Y));
KC_NAND3_X1 T9894 ( .Y(T9894_Y), .B(T3072_Y), .C(T3683_Y),     .A(T3071_Y));
KC_NAND3_X1 T10412 ( .Y(T10412_Y), .B(T416_Y), .C(T6751_Y),     .A(T7533_Y));
KC_NAND3_X1 T9688 ( .Y(T9688_Y), .B(T6989_Y), .C(T494_Y), .A(T416_Y));
KC_NAND3_X1 T9659 ( .Y(T9659_Y), .B(T7347_Y), .C(T458_Y), .A(T416_Y));
KC_NAND3_X1 T9658 ( .Y(T9658_Y), .B(T7185_Y), .C(T461_Y), .A(T416_Y));
KC_NAND3_X1 T9613 ( .Y(T9613_Y), .B(T3072_Y), .C(T2451_Y),     .A(T3071_Y));
KC_NAND3_X1 T9612 ( .Y(T9612_Y), .B(T2451_Y), .C(T6595_Y),     .A(T3072_Y));
KC_NAND3_X1 T9611 ( .Y(T9611_Y), .B(T2451_Y), .C(T1633_Y),     .A(T3071_Y));
KC_NAND3_X1 T10887 ( .Y(T10887_Y), .B(T15855_Y), .C(T15857_Y),     .A(T15858_Y));
KC_NAND3_X1 T10947 ( .Y(T10947_Y), .B(T15942_Y), .C(T15590_Y),     .A(T1778_Q));
KC_NAND3_X1 T9685 ( .Y(T9685_Y), .B(T10386_Y), .C(T15399_Y),     .A(T416_Y));
KC_NAND3_X1 T9684 ( .Y(T9684_Y), .B(T1628_Y), .C(T491_Y), .A(T416_Y));
KC_NAND3_X1 T9683 ( .Y(T9683_Y), .B(T1899_Y), .C(T15400_Y),     .A(T414_Y));
KC_NAND3_X1 T9682 ( .Y(T9682_Y), .B(T6980_Y), .C(T490_Y), .A(T414_Y));
KC_NAND3_X1 T9674 ( .Y(T9674_Y), .B(T1885_Y), .C(T409_Y), .A(T414_Y));
KC_NAND3_X1 T9673 ( .Y(T9673_Y), .B(T1913_Y), .C(T485_Y), .A(T414_Y));
KC_NAND3_X1 T9643 ( .Y(T9643_Y), .B(T1892_Y), .C(T407_Y), .A(T414_Y));
KC_NAND3_X1 T10482 ( .Y(T10482_Y), .B(T1941_Y), .C(T6778_Y),     .A(T416_Y));
KC_NAND3_X1 T10481 ( .Y(T10481_Y), .B(T7481_Y), .C(T6777_Y),     .A(T416_Y));
KC_NAND3_X1 T10480 ( .Y(T10480_Y), .B(T10334_Y), .C(T15692_Y),     .A(T416_Y));
KC_NAND3_X1 T10479 ( .Y(T10479_Y), .B(T1939_Y), .C(T6756_Y),     .A(T416_Y));
KC_NAND3_X1 T9755 ( .Y(T9755_Y), .B(T1648_Y), .C(T6775_Y), .A(T416_Y));
KC_NAND3_X1 T10527 ( .Y(T10527_Y), .B(T10522_Y), .C(T9882_Y),     .A(T1496_Y));
KC_NAND3_X1 T9974 ( .Y(T9974_Y), .B(T12719_Y), .C(T15478_Y),     .A(T2008_Q));
KC_NAND3_X1 T9973 ( .Y(T9973_Y), .B(T16378_Y), .C(T1116_Y),     .A(T1117_Y));
KC_NAND3_X1 T9972 ( .Y(T9972_Y), .B(T10525_Y), .C(T16368_Y),     .A(T1719_Q));
KC_NAND3_X1 T9971 ( .Y(T9971_Y), .B(T2016_Q), .C(T16369_Y),     .A(T1997_Y));
KC_NAND3_X1 T9967 ( .Y(T9967_Y), .B(T9969_Y), .C(T15478_Y),     .A(T2008_Q));
KC_NAND3_X1 T9951 ( .Y(T9951_Y), .B(T9949_Y), .C(T11949_Y),     .A(T2023_Q));
KC_NAND3_X1 T10104 ( .Y(T10104_Y), .B(T10099_Y), .C(T1518_Y),     .A(T2033_Y));
KC_NAND3_X1 T10085 ( .Y(T10085_Y), .B(T12737_Y), .C(T12737_Y),     .A(T1495_Y));
KC_NAND3_X1 T10084 ( .Y(T10084_Y), .B(T2048_Y), .C(T4936_Y),     .A(T1509_Y));
KC_NAND3_X1 T11017 ( .Y(T11017_Y), .B(T11993_Y), .C(T11384_Y),     .A(T4943_Y));
KC_NAND3_X1 T10886 ( .Y(T10886_Y), .B(T11992_Y), .C(T11994_Y),     .A(T2132_Y));
KC_NAND3_X1 T10919 ( .Y(T10919_Y), .B(T11417_Y), .C(T11429_Y),     .A(T2104_Y));
KC_NAND3_X1 T10908 ( .Y(T10908_Y), .B(T11386_Y), .C(T11385_Y),     .A(T2145_Y));
KC_NAND3_X1 T10900 ( .Y(T10900_Y), .B(T8448_Y), .C(T4931_Y),     .A(T5444_Y));
KC_NAND3_X1 T10998 ( .Y(T10998_Y), .B(T13105_Y), .C(T8410_Y),     .A(T2350_Y));
KC_NAND3_X1 T10997 ( .Y(T10997_Y), .B(T12105_Y), .C(T12102_Y),     .A(T12108_Y));
KC_NAND3_X1 T10992 ( .Y(T10992_Y), .B(T16270_Y), .C(T11774_Y),     .A(T12101_Y));
KC_NAND3_X1 T10561 ( .Y(T10561_Y), .B(T12103_Y), .C(T15633_Y),     .A(T12105_Y));
KC_NAND3_X1 T10440 ( .Y(T10440_Y), .B(T1620_Y), .C(T6457_Y),     .A(T414_Y));
KC_NAND3_X1 T10439 ( .Y(T10439_Y), .B(T1914_Y), .C(T406_Y),     .A(T414_Y));
KC_NAND3_X1 T9676 ( .Y(T9676_Y), .B(T5208_Y), .C(T444_Y), .A(T414_Y));
KC_NAND3_X1 T9675 ( .Y(T9675_Y), .B(T1886_Y), .C(T437_Y), .A(T414_Y));
KC_NAND3_X1 T8529 ( .Y(T8529_Y), .B(T3039_Y), .C(T6758_Y), .A(T414_Y));
KC_NAND3_X1 T8528 ( .Y(T8528_Y), .B(T1949_Y), .C(T6757_Y), .A(T416_Y));
KC_NAND3_X1 T9849 ( .Y(T9849_Y), .B(T1132_Y), .C(T10942_Y),     .A(T4872_Y));
KC_NAND3_X1 T10509 ( .Y(T10509_Y), .B(T2522_Y), .C(T15443_Y),     .A(T8453_Y));
KC_NAND3_X1 T10105 ( .Y(T10105_Y), .B(T11662_Y), .C(T2717_Y),     .A(T10100_Y));
KC_NAND3_X1 T10080 ( .Y(T10080_Y), .B(T2612_Y), .C(T10105_Y),     .A(T4982_Y));
KC_NAND3_X1 T10204 ( .Y(T10204_Y), .B(T13051_Q), .C(T2633_Y),     .A(T4898_Y));
KC_NAND3_X1 T10282 ( .Y(T10282_Y), .B(T10276_Y), .C(T142_Y),     .A(T10279_Y));
KC_NAND3_X1 T10281 ( .Y(T10281_Y), .B(T5751_Y), .C(T5754_Y),     .A(T5018_Q));
KC_NAND3_X1 T11009 ( .Y(T11009_Y), .B(T5576_Q), .C(T11961_Y),     .A(T5018_Q));
KC_NAND3_X1 T10897 ( .Y(T10897_Y), .B(T2696_Y), .C(T11361_Y),     .A(T16161_Y));
KC_NAND3_X1 T10896 ( .Y(T10896_Y), .B(T11360_Y), .C(T5019_Y),     .A(T2696_Y));
KC_NAND3_X1 T10891 ( .Y(T10891_Y), .B(T15830_Y), .C(T12149_Y),     .A(T10890_Y));
KC_NAND3_X1 T10890 ( .Y(T10890_Y), .B(T14954_Q), .C(T11009_Y),     .A(T2656_Y));
KC_NAND3_X1 T10913 ( .Y(T10913_Y), .B(T15892_Y), .C(T15041_Y),     .A(T5436_Y));
KC_NAND3_X1 T10909 ( .Y(T10909_Y), .B(T11396_Y), .C(T11383_Y),     .A(T2722_Y));
KC_NAND3_X1 T10899 ( .Y(T10899_Y), .B(T11430_Y), .C(T11368_Y),     .A(T2140_Y));
KC_NAND3_X1 T10930 ( .Y(T10930_Y), .B(T2165_Y), .C(T2171_Y),     .A(T2733_Y));
KC_NAND3_X1 T10929 ( .Y(T10929_Y), .B(T2722_Y), .C(T2171_Y),     .A(T2756_Y));
KC_NAND3_X1 T10928 ( .Y(T10928_Y), .B(T16474_Y), .C(T15881_Y),     .A(T16088_Q));
KC_NAND3_X1 T10933 ( .Y(T10933_Y), .B(T6555_Q), .C(T6526_Q),     .A(T5072_Y));
KC_NAND3_X1 T10932 ( .Y(T10932_Y), .B(T6555_Q), .C(T6549_Q),     .A(T5070_Y));
KC_NAND3_X1 T11030 ( .Y(T11030_Y), .B(T5005_Y), .C(T16105_Y),     .A(T2857_Y));
KC_NAND3_X1 T10971 ( .Y(T10971_Y), .B(T11666_Y), .C(T16057_Y),     .A(T15802_Q));
KC_NAND3_X1 T10967 ( .Y(T10967_Y), .B(T6066_Y), .C(T2842_Q),     .A(T10971_Y));
KC_NAND3_X1 T10959 ( .Y(T10959_Y), .B(T15234_Y), .C(T6086_Y),     .A(T6067_Y));
KC_NAND3_X1 T10976 ( .Y(T10976_Y), .B(T16167_Y), .C(T6085_Y),     .A(T10581_Y));
KC_NAND3_X1 T10611 ( .Y(T10611_Y), .B(T12104_Y), .C(T2874_Q),     .A(T10553_Y));
KC_NAND3_X1 T10610 ( .Y(T10610_Y), .B(T10553_Y), .C(T6183_Y),     .A(T12104_Y));
KC_NAND3_X1 T10596 ( .Y(T10596_Y), .B(T5512_Q), .C(T2866_Y),     .A(T15622_Y));
KC_NAND3_X1 T6581 ( .Y(T6581_Y), .B(T10573_Y), .C(T16131_Y),     .A(T11741_Y));
KC_NAND3_X1 T10988 ( .Y(T10988_Y), .B(T6225_Y), .C(T10573_Y),     .A(T6240_Y));
KC_NAND3_X1 T10987 ( .Y(T10987_Y), .B(T6576_Y), .C(T2893_Y),     .A(T15632_Y));
KC_NAND3_X1 T10986 ( .Y(T10986_Y), .B(T2901_Y), .C(T5518_Y),     .A(T15632_Y));
KC_NAND3_X1 T10985 ( .Y(T10985_Y), .B(T2359_Q), .C(T6559_Y),     .A(T6214_Y));
KC_NAND3_X1 T10978 ( .Y(T10978_Y), .B(T11744_Y), .C(T11746_Y),     .A(T11043_Y));
KC_NAND3_X1 T10977 ( .Y(T10977_Y), .B(T2948_Y), .C(T4054_Y),     .A(T11043_Y));
KC_NAND3_X1 T10881 ( .Y(T10881_Y), .B(T4096_Y), .C(T6531_Y),     .A(T4055_Y));
KC_NAND3_X1 T11005 ( .Y(T11005_Y), .B(T5536_Q), .C(T6162_Y),     .A(T11846_Y));
KC_NAND3_X1 T11000 ( .Y(T11000_Y), .B(T11041_Y), .C(T6531_Y),     .A(T4096_Y));
KC_NAND3_X1 T10999 ( .Y(T10999_Y), .B(T11815_Y), .C(T6537_Y),     .A(T5540_Y));
KC_NAND3_X1 T8151 ( .Y(T8151_Y), .B(T2943_Q), .C(T2944_Q),     .A(T5536_Q));
KC_NAND3_X1 T9651 ( .Y(T9651_Y), .B(T2451_Y), .C(T1633_Y),     .A(T3071_Y));
KC_NAND3_X1 T9650 ( .Y(T9650_Y), .B(T3072_Y), .C(T2451_Y),     .A(T3071_Y));
KC_NAND3_X1 T9649 ( .Y(T9649_Y), .B(T2451_Y), .C(T6595_Y),     .A(T3072_Y));
KC_NAND3_X1 T9737 ( .Y(T9737_Y), .B(T3081_Y), .C(T2451_Y),     .A(T3080_Y));
KC_NAND3_X1 T9736 ( .Y(T9736_Y), .B(T2451_Y), .C(T6595_Y),     .A(T3081_Y));
KC_NAND3_X1 T9834 ( .Y(T9834_Y), .B(T3081_Y), .C(T3683_Y),     .A(T3080_Y));
KC_NAND3_X1 T10895 ( .Y(T10895_Y), .B(T12131_Y), .C(T3204_Y),     .A(T3819_Y));
KC_NAND3_X1 T11022 ( .Y(T11022_Y), .B(T12817_Y), .C(T12817_Y),     .A(T16001_Y));
KC_NAND3_X1 T11029 ( .Y(T11029_Y), .B(T6158_Y), .C(T11028_Y),     .A(T11818_Y));
KC_NAND3_X1 T11028 ( .Y(T11028_Y), .B(T12044_Y), .C(T6177_Y),     .A(T3370_Y));
KC_NAND3_X1 T11019 ( .Y(T11019_Y), .B(T6044_Y), .C(T16036_Y),     .A(T11626_Y));
KC_NAND3_X1 T10973 ( .Y(T10973_Y), .B(T11746_Y), .C(T11029_Y),     .A(T8385_Y));
KC_NAND3_X1 T10970 ( .Y(T10970_Y), .B(T6045_Y), .C(T15612_Y),     .A(T6047_Y));
KC_NAND3_X1 T10966 ( .Y(T10966_Y), .B(T6069_Y), .C(T6051_Y),     .A(T3516_Y));
KC_NAND3_X1 T10965 ( .Y(T10965_Y), .B(T6045_Y), .C(T12829_Y),     .A(T11664_Y));
KC_NAND3_X1 T10964 ( .Y(T10964_Y), .B(T15612_Y), .C(T5072_Y),     .A(T6526_Q));
KC_NAND3_X1 T10962 ( .Y(T10962_Y), .B(T16035_Y), .C(T6048_Y),     .A(T11627_Y));
KC_NAND3_X1 T10961 ( .Y(T10961_Y), .B(T3382_Y), .C(T12829_Y),     .A(T12251_Y));
KC_NAND3_X1 T10975 ( .Y(T10975_Y), .B(T3420_Y), .C(T5522_Y),     .A(T6177_Y));
KC_NAND3_X1 T10974 ( .Y(T10974_Y), .B(T12044_Y), .C(T5522_Y),     .A(T3419_Y));
KC_NAND3_X1 T10625 ( .Y(T10625_Y), .B(T2855_Y), .C(T3425_Y),     .A(T6144_Y));
KC_NAND3_X1 T10621 ( .Y(T10621_Y), .B(T6139_Y), .C(T3454_Y),     .A(T6585_Y));
KC_NAND3_X1 T10609 ( .Y(T10609_Y), .B(T3426_Y), .C(T3424_Y),     .A(T11727_Y));
KC_NAND3_X1 T10588 ( .Y(T10588_Y), .B(T3490_Y), .C(T16141_Y),     .A(T3515_Y));
KC_NAND3_X1 T10995 ( .Y(T10995_Y), .B(T3444_Y), .C(T3448_Y),     .A(T5049_Y));
KC_NAND3_X1 T10991 ( .Y(T10991_Y), .B(T3466_Y), .C(T3465_Y),     .A(T10548_Y));
KC_NAND3_X1 T10990 ( .Y(T10990_Y), .B(T3466_Y), .C(T3465_Y),     .A(T6515_Y));
KC_NAND3_X1 T10984 ( .Y(T10984_Y), .B(T6561_Y), .C(T11763_Y),     .A(T12870_Y));
KC_NAND3_X1 T10979 ( .Y(T10979_Y), .B(T11037_Y), .C(T11746_Y),     .A(T11043_Y));
KC_NAND3_X1 T10882 ( .Y(T10882_Y), .B(T11042_Y), .C(T11822_Y),     .A(T6529_Y));
KC_NAND3_X1 T11007 ( .Y(T11007_Y), .B(T3523_Q), .C(T6514_Y),     .A(T3519_Q));
KC_NAND3_X1 T11006 ( .Y(T11006_Y), .B(T6512_Y), .C(T6490_Y),     .A(T3523_Q));
KC_NAND3_X1 T11004 ( .Y(T11004_Y), .B(T8150_Y), .C(T6512_Y),     .A(T3525_Q));
KC_NAND3_X1 T11003 ( .Y(T11003_Y), .B(T10993_Y), .C(T11829_Y),     .A(T4154_Y));
KC_NAND3_X1 T11002 ( .Y(T11002_Y), .B(T6512_Y), .C(T11832_Y),     .A(T11835_Y));
KC_NAND3_X1 T8521 ( .Y(T8521_Y), .B(T622_Y), .C(T6839_Y), .A(T3677_Y));
KC_NAND3_X1 T8520 ( .Y(T8520_Y), .B(T622_Y), .C(T6802_Y), .A(T3676_Y));
KC_NAND3_X1 T9771 ( .Y(T9771_Y), .B(T622_Y), .C(T6839_Y), .A(T3650_Y));
KC_NAND3_X1 T9770 ( .Y(T9770_Y), .B(T622_Y), .C(T6802_Y), .A(T3653_Y));
KC_NAND3_X1 T9769 ( .Y(T9769_Y), .B(T3650_Y), .C(T622_Y), .A(T3653_Y));
KC_NAND3_X1 T9870 ( .Y(T9870_Y), .B(T622_Y), .C(T6802_Y), .A(T3676_Y));
KC_NAND3_X1 T9833 ( .Y(T9833_Y), .B(T3683_Y), .C(T1633_Y),     .A(T3080_Y));
KC_NAND3_X1 T9832 ( .Y(T9832_Y), .B(T3683_Y), .C(T6595_Y),     .A(T3081_Y));
KC_NAND3_X1 T9830 ( .Y(T9830_Y), .B(T3677_Y), .C(T622_Y), .A(T3676_Y));
KC_NAND3_X1 T9829 ( .Y(T9829_Y), .B(T3683_Y), .C(T6595_Y),     .A(T3081_Y));
KC_NAND3_X1 T9828 ( .Y(T9828_Y), .B(T3081_Y), .C(T3683_Y),     .A(T3080_Y));
KC_NAND3_X1 T9827 ( .Y(T9827_Y), .B(T622_Y), .C(T6839_Y), .A(T3677_Y));
KC_NAND3_X1 T10506 ( .Y(T10506_Y), .B(T3677_Y), .C(T622_Y),     .A(T3676_Y));
KC_NAND3_X1 T10894 ( .Y(T10894_Y), .B(T145_Q), .C(T11410_Y),     .A(T4465_Q));
KC_NAND3_X1 T10893 ( .Y(T10893_Y), .B(T11379_Y), .C(T11365_Y),     .A(T5830_Y));
KC_NAND3_X1 T10892 ( .Y(T10892_Y), .B(T11381_Y), .C(T5802_Y),     .A(T11378_Y));
KC_NAND3_X1 T10889 ( .Y(T10889_Y), .B(T15868_Y), .C(T4486_Y),     .A(T11379_Y));
KC_NAND3_X1 T10885 ( .Y(T10885_Y), .B(T5767_Y), .C(T11984_Y),     .A(T144_Q));
KC_NAND3_X1 T10921 ( .Y(T10921_Y), .B(T5788_Y), .C(T4440_Y),     .A(T14494_Q));
KC_NAND3_X1 T10920 ( .Y(T10920_Y), .B(T14495_Q), .C(T11427_Y),     .A(T145_Q));
KC_NAND3_X1 T10915 ( .Y(T10915_Y), .B(T11408_Y), .C(T5823_Y),     .A(T144_Q));
KC_NAND3_X1 T10911 ( .Y(T10911_Y), .B(T5815_Y), .C(T5789_Y),     .A(T5767_Y));
KC_NAND3_X1 T10903 ( .Y(T10903_Y), .B(T11408_Y), .C(T15845_Y),     .A(T14544_Q));
KC_NAND3_X1 T10898 ( .Y(T10898_Y), .B(T11969_Y), .C(T5763_Y),     .A(T145_Q));
KC_NAND3_X1 T10927 ( .Y(T10927_Y), .B(T15940_Y), .C(T3265_Y),     .A(T12186_Y));
KC_NAND3_X1 T10926 ( .Y(T10926_Y), .B(T3890_Q), .C(T3872_Y),     .A(T3873_Q));
KC_NAND3_X1 T10923 ( .Y(T10923_Y), .B(T5859_Y), .C(T3897_Y),     .A(T3891_Y));
KC_NAND3_X1 T10636 ( .Y(T10636_Y), .B(T3860_Y), .C(T10945_Y),     .A(T10943_Y));
KC_NAND3_X1 T10940 ( .Y(T10940_Y), .B(T3934_Y), .C(T3923_Y),     .A(T3925_Y));
KC_NAND3_X1 T10935 ( .Y(T10935_Y), .B(T15971_Y), .C(T5986_Y),     .A(T11476_Y));
KC_NAND3_X1 T11021 ( .Y(T11021_Y), .B(T16454_Q), .C(T15994_Y),     .A(T15997_Y));
KC_NAND3_X1 T10945 ( .Y(T10945_Y), .B(T11535_Y), .C(T16167_Y),     .A(T3988_Y));
KC_NAND3_X1 T10944 ( .Y(T10944_Y), .B(T4517_Y), .C(T5957_Y),     .A(T5955_Y));
KC_NAND3_X1 T10958 ( .Y(T10958_Y), .B(T5158_Q), .C(T5476_Y),     .A(T4606_Q));
KC_NAND3_X1 T10955 ( .Y(T10955_Y), .B(T4584_Y), .C(T15995_Y),     .A(T10958_Y));
KC_NAND3_X1 T10954 ( .Y(T10954_Y), .B(T10956_Y), .C(T15995_Y),     .A(T10958_Y));
KC_NAND3_X1 T10953 ( .Y(T10953_Y), .B(T15705_Y), .C(T6025_Y),     .A(T6340_Y));
KC_NAND3_X1 T10969 ( .Y(T10969_Y), .B(T6175_Y), .C(T5525_Q),     .A(T5070_Y));
KC_NAND3_X1 T10968 ( .Y(T10968_Y), .B(T5530_Q), .C(T4029_Y),     .A(T11641_Y));
KC_NAND3_X1 T10960 ( .Y(T10960_Y), .B(T3397_Y), .C(T10621_Y),     .A(T15622_Y));
KC_NAND3_X1 T10603 ( .Y(T10603_Y), .B(T6105_Y), .C(T16124_Y),     .A(T8380_Y));
KC_NAND3_X1 T10580 ( .Y(T10580_Y), .B(T6107_Y), .C(T3458_Y),     .A(T11745_Y));
KC_NAND3_X1 T10563 ( .Y(T10563_Y), .B(T2924_Y), .C(T8382_Y),     .A(T16124_Y));
KC_NAND3_X1 T10994 ( .Y(T10994_Y), .B(T4110_Y), .C(T3467_Y),     .A(T4126_Y));
KC_NAND3_X1 T10993 ( .Y(T10993_Y), .B(T11804_Y), .C(T6547_Y),     .A(T6158_Y));
KC_NAND3_X1 T10983 ( .Y(T10983_Y), .B(T4131_Y), .C(T3467_Y),     .A(T4125_Y));
KC_NAND3_X1 T10982 ( .Y(T10982_Y), .B(T4135_Y), .C(T3467_Y),     .A(T4121_Y));
KC_NAND3_X1 T11001 ( .Y(T11001_Y), .B(T6527_Y), .C(T15640_Y),     .A(T11813_Y));
KC_NAND3_X1 T10457 ( .Y(T10457_Y), .B(T9563_Y), .C(T6438_Y),     .A(T4181_Y));
KC_NAND3_X1 T9860 ( .Y(T9860_Y), .B(T2530_Y), .C(T16194_Y),     .A(T12785_Y));
KC_NAND3_X1 T9859 ( .Y(T9859_Y), .B(T2530_Y), .C(T16194_Y),     .A(T12785_Y));
KC_NAND3_X1 T10096 ( .Y(T10096_Y), .B(T12761_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T10095 ( .Y(T10095_Y), .B(T12761_Y), .C(T16194_Y),     .A(T3728_Y));
KC_NAND3_X1 T10888 ( .Y(T10888_Y), .B(T4392_Y), .C(T14943_Q),     .A(T4485_Y));
KC_NAND3_X1 T10914 ( .Y(T10914_Y), .B(T11402_Y), .C(T5788_Y),     .A(T14551_Q));
KC_NAND3_X1 T10910 ( .Y(T10910_Y), .B(T11393_Y), .C(T4486_Y),     .A(T5822_Y));
KC_NAND3_X1 T10902 ( .Y(T10902_Y), .B(T15845_Y), .C(T14942_Q),     .A(T4500_Y));
KC_NAND3_X1 T10901 ( .Y(T10901_Y), .B(T15872_Y), .C(T4383_Y),     .A(T3850_Y));
KC_NAND3_X1 T10925 ( .Y(T10925_Y), .B(T15570_Y), .C(T5862_Y),     .A(T4483_Y));
KC_NAND3_X1 T10924 ( .Y(T10924_Y), .B(T4483_Y), .C(T4492_Q),     .A(T5932_Y));
KC_NAND3_X1 T10922 ( .Y(T10922_Y), .B(T5853_Y), .C(T5854_Y),     .A(T15697_Y));
KC_NAND3_X1 T10631 ( .Y(T10631_Y), .B(T11520_Y), .C(T5932_Y),     .A(T4484_Q));
KC_NAND3_X1 T10939 ( .Y(T10939_Y), .B(T4489_Y), .C(T5929_Y),     .A(T4530_Y));
KC_NAND3_X1 T10938 ( .Y(T10938_Y), .B(T12197_Y), .C(T12209_Y),     .A(T12209_Y));
KC_NAND3_X1 T10937 ( .Y(T10937_Y), .B(T4489_Y), .C(T11453_Y),     .A(T4535_Y));
KC_NAND3_X1 T10931 ( .Y(T10931_Y), .B(T12355_Y), .C(T5889_Y),     .A(T4508_Y));
KC_NAND3_X1 T10951 ( .Y(T10951_Y), .B(T3943_Y), .C(T10943_Y),     .A(T11534_Y));
KC_NAND3_X1 T10950 ( .Y(T10950_Y), .B(T10943_Y), .C(T15592_Y),     .A(T5149_Y));
KC_NAND3_X1 T10948 ( .Y(T10948_Y), .B(T15988_Y), .C(T12229_Y),     .A(T4570_Y));
KC_NAND3_X1 T10943 ( .Y(T10943_Y), .B(T11540_Y), .C(T11537_Y),     .A(T12016_Y));
KC_NAND3_X1 T10957 ( .Y(T10957_Y), .B(T4602_Q), .C(T6016_Y),     .A(T4606_Q));
KC_NAND3_X1 T10576 ( .Y(T10576_Y), .B(T5512_Q), .C(T6104_Y),     .A(T13165_Q));
KC_NAND3_X1 T10989 ( .Y(T10989_Y), .B(T4758_Q), .C(T6203_Y),     .A(T4759_Q));
KC_NAND3_X1 T10981 ( .Y(T10981_Y), .B(T4757_Q), .C(T15629_Y),     .A(T4756_Q));
KC_NAND3_X1 T9477 ( .Y(T9477_Y), .B(T16187_Y), .C(T16189_Y),     .A(T15540_Y));
KC_NAND3_X1 T9372 ( .Y(T9372_Y), .B(T8767_Y), .C(T7644_Y), .A(T902_Y));
KC_NAND3_X1 T9435 ( .Y(T9435_Y), .B(T4872_Y), .C(T10880_Y),     .A(T9031_Y));
KC_NAND3_X1 T9330 ( .Y(T9330_Y), .B(T9329_Y), .C(T11879_Y),     .A(T8732_Y));
KC_NAND3_X1 T9329 ( .Y(T9329_Y), .B(T705_Q), .C(T9332_Y), .A(T6825_Y));
KC_NAND3_X1 T10372 ( .Y(T10372_Y), .B(T403_Y), .C(T6802_Y),     .A(T3653_Y));
KC_NAND3_X1 T10484 ( .Y(T10484_Y), .B(T10335_Y), .C(T15693_Y),     .A(T416_Y));
KC_NAND3_X1 T10483 ( .Y(T10483_Y), .B(T10333_Y), .C(T6753_Y),     .A(T416_Y));
KC_NAND3_X1 T10355 ( .Y(T10355_Y), .B(T10353_Y), .C(T15675_Y),     .A(T416_Y));
KC_NAND3_X1 T10354 ( .Y(T10354_Y), .B(T416_Y), .C(T6752_Y),     .A(T10364_Y));
KC_NAND3_X1 T16266 ( .Y(T16266_Y), .B(T10880_Y), .C(T10942_Y),     .A(T10941_Y));
KC_NAND3_X1 T11026 ( .Y(T11026_Y), .B(T11499_Y), .C(T2153_Q),     .A(T11551_Y));
KC_NAND3_X1 T11012 ( .Y(T11012_Y), .B(T2085_Y), .C(T4944_Y),     .A(T2108_Y));
KC_NAND3_X1 T10560 ( .Y(T10560_Y), .B(T12107_Y), .C(T16131_Y),     .A(T12102_Y));
KC_NAND3_X1 T10559 ( .Y(T10559_Y), .B(T16270_Y), .C(T12103_Y),     .A(T16131_Y));
KC_NAND3_X1 T10528 ( .Y(T10528_Y), .B(T16462_Q), .C(T16369_Y),     .A(T10100_Y));
KC_NAND3_X1 T10476 ( .Y(T10476_Y), .B(T1950_Y), .C(T15686_Y),     .A(T416_Y));
KC_NAND3_X1 T10441 ( .Y(T10441_Y), .B(T1621_Y), .C(T6458_Y),     .A(T414_Y));
KC_NAND3_X1 T11032 ( .Y(T11032_Y), .B(T11831_Y), .C(T6183_Y),     .A(T6182_Y));
KC_NAND3_X1 T11031 ( .Y(T11031_Y), .B(T5006_Y), .C(T16105_Y),     .A(T2857_Y));
KC_NAND3_X1 T11025 ( .Y(T11025_Y), .B(T5070_Y), .C(T6549_Q),     .A(T16035_Y));
KC_NAND3_X1 T11008 ( .Y(T11008_Y), .B(T2678_Y), .C(T5750_Y),     .A(T10281_Y));
KC_NAND3_X1 T10556 ( .Y(T10556_Y), .B(T5514_Y), .C(T11811_Y),     .A(T16133_Y));
KC_NAND3_X1 T10538 ( .Y(T10538_Y), .B(T10244_Y), .C(T10239_Y),     .A(T15815_Q));
KC_NAND3_X1 T10519 ( .Y(T10519_Y), .B(T2570_Q), .C(T5024_Y),     .A(T2584_Q));
KC_NAND3_X1 T10473 ( .Y(T10473_Y), .B(T3038_Y), .C(T15691_Y),     .A(T414_Y));
KC_NAND3_X1 T11018 ( .Y(T11018_Y), .B(T15598_Y), .C(T10961_Y),     .A(T5380_Q));
KC_NAND3_X1 T11015 ( .Y(T11015_Y), .B(T11989_Y), .C(T11990_Y),     .A(T11990_Y));
KC_NAND3_X1 T11014 ( .Y(T11014_Y), .B(T5788_Y), .C(T3844_Y),     .A(T16160_Y));
KC_NAND3_X1 T11027 ( .Y(T11027_Y), .B(T4147_Q), .C(T6045_Y),     .A(T5530_Q));
KC_NAND3_X1 T11024 ( .Y(T11024_Y), .B(T3965_Q), .C(T15587_Y),     .A(T3968_Q));
KC_NAND3_X1 T11023 ( .Y(T11023_Y), .B(T5986_Y), .C(T5973_Y),     .A(T11556_Y));
KC_NAND3_X1 T10505 ( .Y(T10505_Y), .B(T622_Y), .C(T6839_Y),     .A(T3677_Y));
KC_NAND3_X1 T10500 ( .Y(T10500_Y), .B(T622_Y), .C(T6802_Y),     .A(T3676_Y));
KC_NAND3_X1 T10470 ( .Y(T10470_Y), .B(T3677_Y), .C(T622_Y),     .A(T3676_Y));
KC_NAND3_X1 T11020 ( .Y(T11020_Y), .B(T4579_Q), .C(T15584_Y),     .A(T4573_Q));
KC_NAND3_X1 T11013 ( .Y(T11013_Y), .B(T15871_Y), .C(T14942_Q),     .A(T4457_Y));
KC_NAND3_X1 T10433 ( .Y(T10433_Y), .B(T12082_Y), .C(T16194_Y),     .A(T12785_Y));
KC_NAND3_X1 T10432 ( .Y(T10432_Y), .B(T12082_Y), .C(T16194_Y),     .A(T12785_Y));
KC_NAND3_X1 T10425 ( .Y(T10425_Y), .B(T3650_Y), .C(T403_Y),     .A(T3653_Y));
KC_NAND3_X1 T10413 ( .Y(T10413_Y), .B(T3072_Y), .C(T2451_Y),     .A(T3071_Y));
KC_NAND3_X1 T9647 ( .Y(T9647_Y), .B(T10399_Y), .C(T451_Y), .A(T416_Y));
KC_NAND3_X1 T10485 ( .Y(T10485_Y), .B(T10352_Y), .C(T6782_Y),     .A(T416_Y));
KC_NAND3_X1 T9756 ( .Y(T9756_Y), .B(T1645_Y), .C(T6770_Y), .A(T416_Y));
KC_NAND3_X1 T9738 ( .Y(T9738_Y), .B(T2451_Y), .C(T1633_Y),     .A(T3080_Y));
KC_NAND3_X1 T8678 ( .Y(T8678_Y), .B(T695_Q), .C(T7551_Y), .A(T6825_Y));
KC_NAND3_X1 T8658 ( .Y(T8658_Y), .B(T687_Q), .C(T10344_Y),     .A(T6825_Y));
KC_NAND3_X1 T9831 ( .Y(T9831_Y), .B(T3683_Y), .C(T1633_Y),     .A(T3080_Y));
KC_NAND3_X1 T8754 ( .Y(T8754_Y), .B(T7690_Y), .C(T6428_Y),     .A(T16336_Y));
KC_NAND3_X1 T8743 ( .Y(T8743_Y), .B(T8651_Y), .C(T9111_Y), .A(T382_Y));
KC_NAND3_X1 T9923 ( .Y(T9923_Y), .B(T1555_Y), .C(T7986_Y),     .A(T10318_Y));
KC_NAND3_X1 T9419 ( .Y(T9419_Y), .B(T8946_Y), .C(T16478_Y),     .A(T8120_Y));
KC_NAND3_X1 T8774 ( .Y(T8774_Y), .B(T8794_Y), .C(T931_Y), .A(T1095_Q));
KC_NAND3_X1 T10042 ( .Y(T10042_Y), .B(T8032_Y), .C(T1249_Q),     .A(T5376_Q));
KC_NAND3_X1 T8945 ( .Y(T8945_Y), .B(T8118_Y), .C(T16311_Y),     .A(T572_Q));
KC_NAND3_X1 T10904 ( .Y(T10904_Y), .B(T14540_Q), .C(T13307_Y),     .A(T3846_Y));
KC_NAND3_X1 T10949 ( .Y(T10949_Y), .B(T6549_Q), .C(T5070_Y),     .A(T3364_Y));
KC_NAND3_X1 T10946 ( .Y(T10946_Y), .B(T15942_Y), .C(T5983_Y),     .A(T1774_Q));
KC_NAND3_X1 T10956 ( .Y(T10956_Y), .B(T4590_Y), .C(T6022_Y),     .A(T4606_Q));
KC_NAND3_X1 T10952 ( .Y(T10952_Y), .B(T11675_Y), .C(T3516_Y),     .A(T6011_Y));
KC_NAND3_X1 T10972 ( .Y(T10972_Y), .B(T11645_Y), .C(T4021_Y),     .A(T11657_Y));
KC_NAND3_X1 T10963 ( .Y(T10963_Y), .B(T6043_Y), .C(T6044_Y),     .A(T4147_Q));
KC_NAND3_X1 T10591 ( .Y(T10591_Y), .B(T15623_Y), .C(T3436_Y),     .A(T6120_Y));
KC_NAND3_X1 T10996 ( .Y(T10996_Y), .B(T15637_Y), .C(T6207_Y),     .A(T11644_Y));
KC_NAND3_X1 T10980 ( .Y(T10980_Y), .B(T6197_Y), .C(T15633_Y),     .A(T12101_Y));
KC_ADDH_X1 T5644 ( .S(T5644_S), .B(T5641_Co), .Co(T5644_Co),     .A(T45_Q));
KC_ADDH_X1 T5641 ( .S(T5641_S), .B(T5639_Co), .Co(T5641_Co),     .A(T48_Q));
KC_ADDH_X1 T5640 ( .S(T5640_S), .B(T5644_Co), .Co(T5640_Co),     .A(T44_Q));
KC_ADDH_X1 T6850 ( .S(T6850_S), .B(T5643_Co), .Co(T6850_Co),     .A(T54_Q));
KC_ADDH_X1 T5643 ( .S(T5643_S), .B(T5609_Co), .Co(T5643_Co),     .A(T5189_Q));
KC_ADDH_X1 T5642 ( .S(T5642_S), .B(T5625_Co), .Co(T5642_Co),     .A(T5589_Q));
KC_ADDH_X1 T5625 ( .S(T5625_S), .B(T59_Co), .Co(T5625_Co),     .A(T5187_Q));
KC_ADDH_X1 T59 ( .S(T59_S), .B(T6850_Co), .Co(T59_Co), .A(T85_Q));
KC_ADDH_X1 T8993 ( .S(T8993_S), .B(T15099_Y), .Co(T8993_Co),     .A(T8972_Y));
KC_ADDH_X1 T9080 ( .S(T9080_S), .B(T1449_Y), .Co(T9080_Co),     .A(T9135_Y));
KC_ADDH_X1 T6855 ( .S(T6855_S), .B(T11052_Y), .Co(T6855_Co),     .A(T433_Y));
KC_ADDH_X1 T9141 ( .S(T9141_S), .B(T9047_Co), .Co(T9141_Co),     .A(T9469_Q));
KC_ADDH_X1 T9054 ( .S(T9054_S), .B(T9053_Co), .Co(T9054_Co),     .A(T4842_Y));
KC_ADDH_X1 T9053 ( .S(T9053_S), .B(T567_Q), .Co(T9053_Co), .A(T561_Q));
KC_ADDH_X1 T9047 ( .S(T9047_S), .B(T9046_Co), .Co(T9047_Co),     .A(T606_Q));
KC_ADDH_X1 T9046 ( .S(T9046_S), .B(T9054_Co), .Co(T9046_Co),     .A(T605_Q));
KC_ADDH_X1 T9159 ( .S(T9159_S), .B(T9142_Co), .Co(T9159_Co),     .A(T604_Q));
KC_ADDH_X1 T9142 ( .S(T9142_S), .B(T9141_Co), .Co(T9142_Co),     .A(T5406_Q));
KC_ADDH_X1 T9239 ( .S(T9239_S), .B(T781_Q), .Co(T9239_Co), .A(T784_Q));
KC_ADDH_X1 T9225 ( .S(T9225_S), .B(T9224_Co), .Co(T9225_Co),     .A(T5420_Q));
KC_ADDH_X1 T9224 ( .S(T9224_S), .B(T9239_Co), .Co(T9224_Co),     .A(T789_Q));
KC_ADDH_X1 T9188 ( .S(T9188_S), .B(T9225_Co), .Co(T9188_Co),     .A(T1022_Q));
KC_ADDH_X1 T6097 ( .S(T6097_S), .B(T2098_Y), .Co(T6097_Co),     .A(T2099_Y));
KC_ADDH_X1 T5825 ( .S(T5825_S), .B(T881_Y), .Co(T5825_Co),     .A(T2540_Y));
KC_ADDH_X1 T5869 ( .S(T5869_S), .B(T2573_Y), .Co(T5869_Co),     .A(T16412_Y));
KC_ADDH_X1 T6133 ( .S(T6133_S), .B(T2164_Y), .Co(T6133_Co),     .A(T2744_Y));
KC_ADDH_X1 T6231 ( .S(T6231_S), .B(T3295_Y), .Co(T6231_Co),     .A(T3303_Y));
KC_ADDH_X1 T6230 ( .S(T6230_S), .B(T3296_Y), .Co(T6230_Co),     .A(T5942_Y));
KC_ADDH_X1 T6776 ( .S(T6776_S), .B(T16002_Y), .Co(T6776_Co),     .A(T3327_Y));
KC_ADDH_X1 T6320 ( .S(T6320_S), .B(T6335_Y), .Co(T6320_Co),     .A(T7915_Y));
KC_ADDH_X1 T6031 ( .S(T6031_S), .B(T15554_Y), .Co(T6031_Co),     .A(T11315_Y));
KC_ADDH_X1 T6797 ( .S(T6797_S), .B(T15939_Y), .Co(T6797_Co),     .A(T3924_Y));
KC_ADDH_X1 T6146 ( .S(T6146_S), .B(T6142_Co), .Co(T6146_Co),     .A(T3877_Q));
KC_ADDH_X1 T6143 ( .S(T6143_S), .B(T6130_Co), .Co(T6143_Co),     .A(T3895_Q));
KC_ADDH_X1 T6142 ( .S(T6142_S), .B(T6132_Co), .Co(T6142_Co),     .A(T3878_Q));
KC_ADDH_X1 T6132 ( .S(T6132_S), .B(T6131_Co), .Co(T6132_Co),     .A(T5130_Q));
KC_ADDH_X1 T6131 ( .S(T6131_S), .B(T6143_Co), .Co(T6131_Co),     .A(T3883_Q));
KC_ADDH_X1 T6842 ( .S(T6842_S), .B(T6503_Co), .Co(T6842_Co),     .A(T15760_Q));
KC_ADDH_X1 T6841 ( .S(T6841_S), .B(T6504_Co), .Co(T6841_Co),     .A(T5528_Q));
KC_ADDH_X1 T6840 ( .S(T6840_S), .B(T3528_Q), .Co(T6840_Co),     .A(T4178_Q));
KC_ADDH_X1 T6534 ( .S(T6534_S), .B(T6549_Q), .Co(T6534_Co),     .A(T6526_Q));
KC_ADDH_X1 T6533 ( .S(T6533_S), .B(T6534_Co), .Co(T6533_Co),     .A(T6555_Q));
KC_ADDH_X1 T6504 ( .S(T6504_S), .B(T6840_Co), .Co(T6504_Co),     .A(T5532_Q));
KC_ADDH_X1 T6503 ( .S(T6503_S), .B(T6568_Co), .Co(T6503_Co),     .A(T5530_Q));
KC_ADDH_X1 T6614 ( .S(T6614_S), .B(T6591_Co), .Co(T6614_Co),     .A(T4164_Q));
KC_ADDH_X1 T6611 ( .S(T6611_S), .B(T6610_Co), .Co(T6611_Co),     .A(T4168_Q));
KC_ADDH_X1 T6610 ( .S(T6610_S), .B(T6614_Co), .Co(T6610_Co),     .A(T4171_Q));
KC_ADDH_X1 T6591 ( .S(T6591_S), .B(T6841_Co), .Co(T6591_Co),     .A(T4163_Q));
KC_ADDH_X1 T6590 ( .S(T6590_S), .B(T6842_Co), .Co(T6590_Co),     .A(T4179_Q));
KC_ADDH_X1 T6194 ( .S(T6194_S), .B(T4529_Y), .Co(T6194_Co),     .A(T4531_Y));
KC_ADDH_X1 T6420 ( .S(T6420_S), .B(T4754_Y), .Co(T6420_Co),     .A(T4717_Q));
KC_ADDH_X1 T6686 ( .S(T6686_S), .B(T4973_Y), .Co(T6686_Co),     .A(T635_Y));
KC_ADDH_X1 T5639 ( .S(T5639_S), .B(T5642_Co), .Co(T5639_Co),     .A(T5190_Q));
KC_ADDH_X1 T5609 ( .S(T5609_S), .B(T5220_Q), .Co(T5609_Co),     .A(T5184_Q));
KC_ADDH_X1 T6168 ( .S(T6168_S), .B(T3885_Q), .Co(T6168_Co),     .A(T4493_Q));
KC_ADDH_X1 T6167 ( .S(T6167_S), .B(T6168_Co), .Co(T6167_Co),     .A(T4491_Q));
KC_ADDH_X1 T6130 ( .S(T6130_S), .B(T6167_Co), .Co(T6130_Co),     .A(T3900_Q));
KC_ADDH_X1 T6568 ( .S(T6568_S), .B(T6567_Co), .Co(T6568_Co),     .A(T4147_Q));
KC_ADDH_X1 T6567 ( .S(T6567_S), .B(T6533_Co), .Co(T6567_Co),     .A(T5525_Q));
KC_NOR3_X1 T5628 ( .Y(T5628_Y), .B(T52_Y), .C(T5637_Y), .A(T79_Y));
KC_NOR3_X1 T5627 ( .Y(T5627_Y), .B(T5189_Q), .C(T8550_Y), .A(T48_Q));
KC_NOR3_X1 T55 ( .Y(T55_Y), .B(T5589_Q), .C(T5190_Q), .A(T44_Q));
KC_NOR3_X1 T5600 ( .Y(T5600_Y), .B(T12471_Y), .C(T5601_Y),     .A(T8538_Y));
KC_NOR3_X1 T5599 ( .Y(T5599_Y), .B(T12472_Y), .C(T12367_Y),     .A(T8544_Y));
KC_NOR3_X1 T9287 ( .Y(T9287_Y), .B(T260_Y), .C(T9288_Y), .A(T133_Q));
KC_NOR3_X1 T6968 ( .Y(T6968_Y), .B(T6969_Y), .C(T6971_Y), .A(T8608_Y));
KC_NOR3_X1 T9271 ( .Y(T9271_Y), .B(T5192_Q), .C(T9272_Y), .A(T131_Q));
KC_NOR3_X1 T9270 ( .Y(T9270_Y), .B(T257_Y), .C(T12382_Y), .A(T6319_Y));
KC_NOR3_X1 T7696 ( .Y(T7696_Y), .B(T224_Q), .C(T12418_Y), .A(T4803_Q));
KC_NOR3_X1 T7695 ( .Y(T7695_Y), .B(T16006_Y), .C(T908_Y), .A(T106_Q));
KC_NOR3_X1 T7681 ( .Y(T7681_Y), .B(T212_Q), .C(T7680_Y), .A(T207_Q));
KC_NOR3_X1 T7677 ( .Y(T7677_Y), .B(T15430_Y), .C(T7680_Y), .A(T647_Y));
KC_NOR3_X1 T7676 ( .Y(T7676_Y), .B(T207_Q), .C(T7678_Y), .A(T4803_Q));
KC_NOR3_X1 T7582 ( .Y(T7582_Y), .B(T645_Y), .C(T12418_Y), .A(T802_Y));
KC_NOR3_X1 T7581 ( .Y(T7581_Y), .B(T223_Q), .C(T645_Y), .A(T4803_Q));
KC_NOR3_X1 T7580 ( .Y(T7580_Y), .B(T223_Q), .C(T212_Q), .A(T224_Q));
KC_NOR3_X1 T6970 ( .Y(T6970_Y), .B(T9287_Y), .C(T6969_Y),     .A(T15354_Y));
KC_NOR3_X1 T6969 ( .Y(T6969_Y), .B(T5192_Q), .C(T6932_Y), .A(T5222_Q));
KC_NOR3_X1 T7660 ( .Y(T7660_Y), .B(T11183_Y), .C(T7566_Y),     .A(T11203_Y));
KC_NOR3_X1 T8072 ( .Y(T8072_Y), .B(T1323_Y), .C(T560_Y), .A(T566_Q));
KC_NOR3_X1 T8071 ( .Y(T8071_Y), .B(T8073_Y), .C(T8947_Y), .A(T5378_Q));
KC_NOR3_X1 T8070 ( .Y(T8070_Y), .B(T8065_Y), .C(T8947_Y), .A(T566_Q));
KC_NOR3_X1 T8059 ( .Y(T8059_Y), .B(T1323_Y), .C(T8062_Y), .A(T5378_Q));
KC_NOR3_X1 T8045 ( .Y(T8045_Y), .B(T8059_Y), .C(T8070_Y), .A(T5608_Y));
KC_NOR3_X1 T9164 ( .Y(T9164_Y), .B(T604_Q), .C(T9140_Y), .A(T9472_Q));
KC_NOR3_X1 T9145 ( .Y(T9145_Y), .B(T604_Q), .C(T9140_Y), .A(T9472_Q));
KC_NOR3_X1 T9144 ( .Y(T9144_Y), .B(T604_Q), .C(T9140_Y), .A(T9472_Q));
KC_NOR3_X1 T9102 ( .Y(T9102_Y), .B(T9472_Q), .C(T9065_Y), .A(T605_Q));
KC_NOR3_X1 T7263 ( .Y(T7263_Y), .B(T7417_Y), .C(T7093_Y), .A(T9276_Y));
KC_NOR3_X1 T7244 ( .Y(T7244_Y), .B(T7115_Y), .C(T7119_Y), .A(T7393_Y));
KC_NOR3_X1 T9242 ( .Y(T9242_Y), .B(T16511_Y), .C(T9226_Y),     .A(T9241_Y));
KC_NOR3_X1 T7555 ( .Y(T7555_Y), .B(T10942_Y), .C(T744_Y), .A(T7839_Y));
KC_NOR3_X1 T7838 ( .Y(T7838_Y), .B(T9393_Y), .C(T926_Y), .A(T4353_Y));
KC_NOR3_X1 T8996 ( .Y(T8996_Y), .B(T4847_Y), .C(T9436_Y),     .A(T16006_Y));
KC_NOR3_X1 T8058 ( .Y(T8058_Y), .B(T15800_Y), .C(T8975_Y), .A(T982_Q));
KC_NOR3_X1 T8031 ( .Y(T8031_Y), .B(T7879_Y), .C(T989_Y), .A(T9403_Y));
KC_NOR3_X1 T10048 ( .Y(T10048_Y), .B(T1133_Q), .C(T980_Q),     .A(T15500_Y));
KC_NOR3_X1 T10027 ( .Y(T10027_Y), .B(T10660_Y), .C(T8057_Y),     .A(T10004_Y));
KC_NOR3_X1 T8032 ( .Y(T8032_Y), .B(T1130_Q), .C(T927_Y), .A(T1133_Q));
KC_NOR3_X1 T10022 ( .Y(T10022_Y), .B(T10170_Y), .C(T7951_Y),     .A(T16119_Y));
KC_NOR3_X1 T10001 ( .Y(T10001_Y), .B(T10021_Y), .C(T10315_Y),     .A(T16118_Y));
KC_NOR3_X1 T10000 ( .Y(T10000_Y), .B(T11914_Y), .C(T12446_Y),     .A(T10152_Y));
KC_NOR3_X1 T1275 ( .Y(T1275_Y), .B(T1505_Y), .C(T13059_Q),     .A(T13054_Q));
KC_NOR3_X1 T7338 ( .Y(T7338_Y), .B(T3650_Y), .C(T7339_Y), .A(T3653_Y));
KC_NOR3_X1 T1359 ( .Y(T1359_Y), .B(T1357_Y), .C(T4825_Y), .A(T1738_Y));
KC_NOR3_X1 T7779 ( .Y(T7779_Y), .B(T4920_Y), .C(T10757_Y), .A(T803_Y));
KC_NOR3_X1 T8001 ( .Y(T8001_Y), .B(T3650_Y), .C(T8004_Y), .A(T3653_Y));
KC_NOR3_X1 T1743 ( .Y(T1743_Y), .B(T5380_Q), .C(T1744_Y),     .A(T16301_Q));
KC_NOR3_X1 T1764 ( .Y(T1764_Y), .B(T5903_Y), .C(T1772_Y), .A(T5945_Y));
KC_NOR3_X1 T1765 ( .Y(T1765_Y), .B(T5452_Q), .C(T2175_Y), .A(T2150_Q));
KC_NOR3_X1 T1767 ( .Y(T1767_Y), .B(T1769_Y), .C(T1770_Y),     .A(T15515_Y));
KC_NOR3_X1 T1769 ( .Y(T1769_Y), .B(T5452_Q), .C(T1772_Y), .A(T2150_Q));
KC_NOR3_X1 T1770 ( .Y(T1770_Y), .B(T5903_Y), .C(T5460_Y), .A(T5945_Y));
KC_NOR3_X1 T1997 ( .Y(T1997_Y), .B(T2005_Q), .C(T16378_Y),     .A(T2028_Q));
KC_NOR3_X1 T2033 ( .Y(T2033_Y), .B(T12100_Y), .C(T15812_Y),     .A(T12099_Y));
KC_NOR3_X1 T2100 ( .Y(T2100_Y), .B(T12165_Y), .C(T12165_Y),     .A(T5820_Y));
KC_NOR3_X1 T6324 ( .Y(T6324_Y), .B(T8317_Y), .C(T8326_Y), .A(T8318_Y));
KC_NOR3_X1 T2230 ( .Y(T2230_Y), .B(T2229_Y), .C(T2227_Y), .A(T2228_Y));
KC_NOR3_X1 T2263 ( .Y(T2263_Y), .B(T8470_Y), .C(T8347_Y), .A(T8353_Y));
KC_NOR3_X1 T2264 ( .Y(T2264_Y), .B(T8352_Q), .C(T16082_Q),     .A(T15138_Q));
KC_NOR3_X1 T2320 ( .Y(T2320_Y), .B(T6571_Y), .C(T12101_Y),     .A(T6225_Y));
KC_NOR3_X1 T2329 ( .Y(T2329_Y), .B(T10997_Y), .C(T5517_Y),     .A(T15633_Y));
KC_NOR3_X1 T2340 ( .Y(T2340_Y), .B(T2365_Y), .C(T2375_Y), .A(T3464_Y));
KC_NOR3_X1 T2550 ( .Y(T2550_Y), .B(T2545_Y), .C(T16363_Y),     .A(T2571_Q));
KC_NOR3_X1 T2562 ( .Y(T2562_Y), .B(T2561_Y), .C(T15477_Y),     .A(T5869_Co));
KC_NOR3_X1 T2656 ( .Y(T2656_Y), .B(T10271_Y), .C(T10242_Y),     .A(T10244_Y));
KC_NOR3_X1 T2702 ( .Y(T2702_Y), .B(T15804_Q), .C(T15807_Q),     .A(T15803_Q));
KC_NOR3_X1 T2727 ( .Y(T2727_Y), .B(T2726_Y), .C(T2725_Y), .A(T2728_Y));
KC_NOR3_X1 T2806 ( .Y(T2806_Y), .B(T12357_Y), .C(T964_Q),     .A(T16474_Y));
KC_NOR3_X1 T2819 ( .Y(T2819_Y), .B(T12322_Y), .C(T15615_Y),     .A(T2854_Y));
KC_NOR3_X1 T2823 ( .Y(T2823_Y), .B(T6214_Y), .C(T5512_Q), .A(T2839_Y));
KC_NOR3_X1 T2851 ( .Y(T2851_Y), .B(T6182_Y), .C(T6180_Y), .A(T2874_Q));
KC_NOR3_X1 T2855 ( .Y(T2855_Y), .B(T3425_Y), .C(T16084_Y),     .A(T2870_Y));
KC_NOR3_X1 T2856 ( .Y(T2856_Y), .B(T12065_Y), .C(T2859_Y),     .A(T6506_Y));
KC_NOR3_X1 T2857 ( .Y(T2857_Y), .B(T2860_Y), .C(T12853_Y),     .A(T6124_Y));
KC_NOR3_X1 T2906 ( .Y(T2906_Y), .B(T6192_Y), .C(T2915_Y), .A(T2910_Y));
KC_NOR3_X1 T3032 ( .Y(T3032_Y), .B(T2589_Y), .C(T3031_Y), .A(T3640_Y));
KC_NOR3_X1 T3054 ( .Y(T3054_Y), .B(T3081_Y), .C(T3051_Y), .A(T3080_Y));
KC_NOR3_X1 T3205 ( .Y(T3205_Y), .B(T12776_Y), .C(T5765_Y),     .A(T5765_Y));
KC_NOR3_X1 T3206 ( .Y(T3206_Y), .B(T11355_Y), .C(T12148_Y),     .A(T10243_Y));
KC_NOR3_X1 T3249 ( .Y(T3249_Y), .B(T15911_Y), .C(T15911_Y),     .A(T3278_Y));
KC_NOR3_X1 T3293 ( .Y(T3293_Y), .B(T3296_Y), .C(T3345_Y), .A(T3315_Y));
KC_NOR3_X1 T3318 ( .Y(T3318_Y), .B(T11022_Y), .C(T8273_Y),     .A(T6256_Y));
KC_NOR3_X1 T3320 ( .Y(T3320_Y), .B(T15579_Y), .C(T15982_Y),     .A(T5483_Y));
KC_NOR3_X1 T3321 ( .Y(T3321_Y), .B(T12963_Y), .C(T8486_Y),     .A(T8486_Y));
KC_NOR3_X1 T3346 ( .Y(T3346_Y), .B(T5478_Y), .C(T3340_Y), .A(T3349_Y));
KC_NOR3_X1 T3350 ( .Y(T3350_Y), .B(T3347_Y), .C(T16014_Y),     .A(T5478_Y));
KC_NOR3_X1 T3353 ( .Y(T3353_Y), .B(T3349_Y), .C(T3340_Y),     .A(T16014_Y));
KC_NOR3_X1 T3399 ( .Y(T3399_Y), .B(T3382_Y), .C(T5492_Y),     .A(T10962_Y));
KC_NOR3_X1 T3418 ( .Y(T3418_Y), .B(T3415_Y), .C(T5503_Y), .A(T6138_Y));
KC_NOR3_X1 T3419 ( .Y(T3419_Y), .B(T12045_Y), .C(T12877_Y),     .A(T16148_Y));
KC_NOR3_X1 T3420 ( .Y(T3420_Y), .B(T15616_Y), .C(T3416_Y),     .A(T16148_Y));
KC_NOR3_X1 T3442 ( .Y(T3442_Y), .B(T16141_Y), .C(T3385_Y),     .A(T3389_Y));
KC_NOR3_X1 T3517 ( .Y(T3517_Y), .B(T6510_Y), .C(T3510_Y), .A(T6512_Y));
KC_NOR3_X1 T3623 ( .Y(T3623_Y), .B(T5331_Y), .C(T3626_Y), .A(T5134_Y));
KC_NOR3_X1 T3636 ( .Y(T3636_Y), .B(T3650_Y), .C(T3621_Y), .A(T3653_Y));
KC_NOR3_X1 T3657 ( .Y(T3657_Y), .B(T9869_Y), .C(T3707_Y), .A(T3680_Y));
KC_NOR3_X1 T3792 ( .Y(T3792_Y), .B(T3202_Y), .C(T11330_Y),     .A(T15834_Y));
KC_NOR3_X1 T3813 ( .Y(T3813_Y), .B(T6041_Y), .C(T3812_Y),     .A(T11323_Y));
KC_NOR3_X1 T3814 ( .Y(T3814_Y), .B(T5430_Y), .C(T3810_Y),     .A(T12134_Y));
KC_NOR3_X1 T3828 ( .Y(T3828_Y), .B(T15888_Y), .C(T3856_Y),     .A(T11353_Y));
KC_NOR3_X1 T3838 ( .Y(T3838_Y), .B(T3241_Y), .C(T5842_Y), .A(T3242_Q));
KC_NOR3_X1 T3846 ( .Y(T3846_Y), .B(T5795_Y), .C(T5774_Y),     .A(T15871_Y));
KC_NOR3_X1 T3911 ( .Y(T3911_Y), .B(T12814_Y), .C(T11512_Y),     .A(T11484_Y));
KC_NOR3_X1 T3948 ( .Y(T3948_Y), .B(T5984_Y), .C(T15587_Y),     .A(T11576_Y));
KC_NOR3_X1 T3980 ( .Y(T3980_Y), .B(T3977_Y), .C(T12019_Y),     .A(T11618_Y));
KC_NOR3_X1 T4022 ( .Y(T4022_Y), .B(T6044_Y), .C(T10969_Y),     .A(T4179_Q));
KC_NOR3_X1 T4023 ( .Y(T4023_Y), .B(T10969_Y), .C(T4049_Y),     .A(T6043_Y));
KC_NOR3_X1 T4028 ( .Y(T4028_Y), .B(T4026_Y), .C(T4109_Y), .A(T3384_Y));
KC_NOR3_X1 T4029 ( .Y(T4029_Y), .B(T6048_Y), .C(T4032_Y), .A(T4176_Q));
KC_NOR3_X1 T4081 ( .Y(T4081_Y), .B(T4024_Y), .C(T5525_Q), .A(T4049_Y));
KC_NOR3_X1 T4087 ( .Y(T4087_Y), .B(T6134_Y), .C(T4083_Y), .A(T2752_Q));
KC_NOR3_X1 T4159 ( .Y(T4159_Y), .B(T4160_Y), .C(T4167_Y), .A(T4162_Y));
KC_NOR3_X1 T4181 ( .Y(T4181_Y), .B(T4191_Y), .C(T9563_Y),     .A(T12473_Y));
KC_NOR3_X1 T4271 ( .Y(T4271_Y), .B(T12656_Y), .C(T13900_Q),     .A(T5173_Y));
KC_NOR3_X1 T4397 ( .Y(T4397_Y), .B(T11365_Y), .C(T15832_Y),     .A(T5800_Y));
KC_NOR3_X1 T4466 ( .Y(T4466_Y), .B(T5854_Y), .C(T5778_Y),     .A(T14548_Q));
KC_NOR3_X1 T4469 ( .Y(T4469_Y), .B(T15572_Y), .C(T5873_Y),     .A(T5142_Y));
KC_NOR3_X1 T4474 ( .Y(T4474_Y), .B(T15935_Y), .C(T4497_Y),     .A(T10924_Y));
KC_NOR3_X1 T4475 ( .Y(T4475_Y), .B(T15934_Y), .C(T10628_Y),     .A(T4477_Y));
KC_NOR3_X1 T4476 ( .Y(T4476_Y), .B(T4708_Y), .C(T4495_Y), .A(T6165_Y));
KC_NOR3_X1 T4477 ( .Y(T4477_Y), .B(T4497_Y), .C(T10631_Y),     .A(T4492_Q));
KC_NOR3_X1 T4480 ( .Y(T4480_Y), .B(T4501_Y), .C(T6127_Y), .A(T5857_Y));
KC_NOR3_X1 T4512 ( .Y(T4512_Y), .B(T11507_Y), .C(T5139_Y),     .A(T15706_Y));
KC_NOR3_X1 T4513 ( .Y(T4513_Y), .B(T12959_Y), .C(T4511_Y),     .A(T4534_Y));
KC_NOR3_X1 T4514 ( .Y(T4514_Y), .B(T5892_Y), .C(T5907_Y),     .A(T11574_Y));
KC_NOR3_X1 T4517 ( .Y(T4517_Y), .B(T4516_Y), .C(T10925_Y),     .A(T4530_Y));
KC_NOR3_X1 T4518 ( .Y(T4518_Y), .B(T4535_Y), .C(T4489_Y), .A(T4530_Y));
KC_NOR3_X1 T4521 ( .Y(T4521_Y), .B(T4526_Q), .C(T4528_Q), .A(T4527_Q));
KC_NOR3_X1 T4552 ( .Y(T4552_Y), .B(T11573_Y), .C(T4571_Y),     .A(T10948_Y));
KC_NOR3_X1 T4561 ( .Y(T4561_Y), .B(T5157_Y), .C(T5947_Y), .A(T4556_Y));
KC_NOR3_X1 T4585 ( .Y(T4585_Y), .B(T4582_Y), .C(T6010_Y), .A(T4611_Y));
KC_NOR3_X1 T4586 ( .Y(T4586_Y), .B(T6016_Y), .C(T15604_Y),     .A(T4606_Q));
KC_NOR3_X1 T4587 ( .Y(T4587_Y), .B(T4602_Q), .C(T6021_Y), .A(T5159_Q));
KC_NOR3_X1 T4588 ( .Y(T4588_Y), .B(T4581_Y), .C(T10957_Y),     .A(T15604_Y));
KC_NOR3_X1 T4589 ( .Y(T4589_Y), .B(T15604_Y), .C(T4580_Y),     .A(T4602_Q));
KC_NOR3_X1 T4590 ( .Y(T4590_Y), .B(T15609_Y), .C(T15604_Y),     .A(T5158_Q));
KC_NOR3_X1 T4740 ( .Y(T4740_Y), .B(T4756_Q), .C(T4757_Q), .A(T4755_Q));
KC_NOR3_X1 T4743 ( .Y(T4743_Y), .B(T4758_Q), .C(T4759_Q), .A(T4760_Q));
KC_NOR3_X1 T9390 ( .Y(T9390_Y), .B(T15195_Y), .C(T7698_Y),     .A(T16318_Y));
KC_NOR3_X1 T9431 ( .Y(T9431_Y), .B(T1394_Y), .C(T9987_Y), .A(T4847_Y));
KC_NOR3_X1 T10297 ( .Y(T10297_Y), .B(T13121_Y), .C(T10171_Y),     .A(T16275_Y));
KC_NOR3_X1 T5109 ( .Y(T5109_Y), .B(T16143_Y), .C(T12071_Y),     .A(T4164_Q));
KC_NOR3_X1 T5115 ( .Y(T5115_Y), .B(T8163_Y), .C(T4761_Y), .A(T4180_Y));
KC_NOR3_X1 T5140 ( .Y(T5140_Y), .B(T4568_Q), .C(T5914_Y),     .A(T11570_Y));
KC_NOR3_X1 T5598 ( .Y(T5598_Y), .B(T5596_Y), .C(T5604_Y),     .A(T15316_Y));
KC_NOR3_X1 T8118 ( .Y(T8118_Y), .B(T5377_Q), .C(T8065_Y), .A(T556_Q));
KC_NOR3_X1 T8088 ( .Y(T8088_Y), .B(T15488_Y), .C(T8106_Y),     .A(T12723_Y));
KC_NOR3_X1 T5367 ( .Y(T5367_Y), .B(T5388_Q), .C(T16268_Y),     .A(T2957_Y));
KC_NOR3_X1 T9096 ( .Y(T9096_Y), .B(T5406_Q), .C(T9097_Y), .A(T606_Q));
KC_NOR3_X1 T5437 ( .Y(T5437_Y), .B(T5827_Y), .C(T5816_Y),     .A(T16154_Y));
KC_NOR3_X1 T5476 ( .Y(T5476_Y), .B(T4602_Q), .C(T15609_Y),     .A(T5159_Q));
KC_NOR3_X1 T5491 ( .Y(T5491_Y), .B(T4024_Y), .C(T4033_Y), .A(T3354_Y));
KC_NOR3_X1 T5515 ( .Y(T5515_Y), .B(T6225_Y), .C(T10992_Y),     .A(T12103_Y));
KC_OAI211B_X1 T5612 ( .C0N(T11262_Y), .B(T5599_Y), .A(T8557_Y),     .C1(T69_Y), .Y(T5612_Y));
KC_OAI211B_X1 T6856 ( .C0N(T5613_Y), .B(T14991_Y), .A(T5602_Y),     .C1(T6359_Q), .Y(T6856_Y));
KC_OAI211B_X1 T8989 ( .C0N(T1602_Y), .B(T247_Y), .A(T15091_Y),     .C1(T15489_Y), .Y(T8989_Y));
KC_OAI211B_X1 T7912 ( .C0N(T7863_Y), .B(T8874_Y), .A(T16418_Y),     .C1(T8872_Y), .Y(T7912_Y));
KC_OAI211B_X1 T7814 ( .C0N(T7578_Y), .B(T8785_Y), .A(T16327_Y),     .C1(T8780_Y), .Y(T7814_Y));
KC_OAI211B_X1 T9283 ( .C0N(T450_Q), .B(T297_Y), .A(T6272_Y),     .C1(T439_Q), .Y(T9283_Y));
KC_OAI211B_X1 T7893 ( .C0N(T5346_Q), .B(T16358_Y), .A(T15789_Y),     .C1(T16463_Y), .Y(T7893_Y));
KC_OAI211B_X1 T9055 ( .C0N(T605_Q), .B(T1587_Y), .A(T15801_Y),     .C1(T9062_Y), .Y(T9055_Y));
KC_OAI211B_X1 T5647 ( .C0N(T7533_Y), .B(T14739_Q), .A(T5028_Y),     .C1(T6765_Y), .Y(T5647_Y));
KC_OAI211B_X1 T2043 ( .C0N(T2042_Y), .B(T2058_Y), .A(T2058_Y),     .C1(T1495_Y), .Y(T2043_Y));
KC_OAI211B_X1 T2375 ( .C0N(T15645_Y), .B(T16472_Y), .A(T15645_Y),     .C1(T2365_Y), .Y(T2375_Y));
KC_OAI211B_X1 T2523 ( .C0N(T2540_Y), .B(T2540_Y), .A(T5825_Co),     .C1(T16169_Y), .Y(T2523_Y));
KC_OAI211B_X1 T2596 ( .C0N(T3741_Y), .B(T14342_Q), .A(T10239_Y),     .C1(T1114_Y), .Y(T2596_Y));
KC_OAI211B_X1 T2613 ( .C0N(T10064_Y), .B(T2624_Y), .A(T12098_Y),     .C1(T2625_Q), .Y(T2613_Y));
KC_OAI211B_X1 T2731 ( .C0N(T3283_Y), .B(T2753_Y), .A(T6150_Y),     .C1(T6133_Co), .Y(T2731_Y));
KC_OAI211B_X1 T3251 ( .C0N(T8352_Q), .B(T5447_Y), .A(T11522_Y),     .C1(T4471_Y), .Y(T3251_Y));
KC_OAI211B_X1 T3253 ( .C0N(T3252_Y), .B(T3269_Y), .A(T8223_Y),     .C1(T3254_Y), .Y(T3253_Y));
KC_OAI211B_X1 T3289 ( .C0N(T5922_Y), .B(T3298_Y), .A(T5921_Y),     .C1(T5921_Y), .Y(T3289_Y));
KC_OAI211B_X1 T3300 ( .C0N(T3286_Y), .B(T5921_Y), .A(T3289_Y),     .C1(T5067_Y), .Y(T3300_Y));
KC_OAI211B_X1 T3507 ( .C0N(T11817_Y), .B(T10993_Y), .A(T4155_Y),     .C1(T8430_Y), .Y(T3507_Y));
KC_OAI211B_X1 T3865 ( .C0N(T15138_Q), .B(T3862_Y), .A(T3920_Y),     .C1(T4471_Y), .Y(T3865_Y));
KC_OAI211B_X1 T3869 ( .C0N(T3884_Q), .B(T6228_Y), .A(T3867_Y),     .C1(T4471_Y), .Y(T3869_Y));
KC_OAI211B_X1 T3981 ( .C0N(T11577_Y), .B(T4583_Y), .A(T10956_Y),     .C1(T10958_Y), .Y(T3981_Y));
KC_OAI211B_X1 T4138 ( .C0N(T6503_S), .B(T4124_Y), .A(T12294_Y),     .C1(T6558_Y), .Y(T4138_Y));
KC_OAI211B_X1 T4153 ( .C0N(T4180_Y), .B(T8166_Y), .A(T3996_Y),     .C1(T3996_Y), .Y(T4153_Y));
KC_OAI211B_X1 T4162 ( .C0N(T11842_Y), .B(T4156_Y), .A(T4166_Y),     .C1(T9163_Y), .Y(T4162_Y));
KC_OAI211B_X1 T4451 ( .C0N(T11377_Y), .B(T12795_Y), .A(T11390_Y),     .C1(T6741_Y), .Y(T4451_Y));
KC_OAI211B_X1 T4543 ( .C0N(T3940_Y), .B(T4563_Y), .A(T15966_Y),     .C1(T4563_Y), .Y(T4543_Y));
KC_OAI211B_X1 T4591 ( .C0N(T4599_Y), .B(T8320_Y), .A(T4592_Y),     .C1(T4585_Y), .Y(T4591_Y));
KC_OAI211B_X1 T4592 ( .C0N(T4585_Y), .B(T6018_Y), .A(T4621_Y),     .C1(T6018_Y), .Y(T4592_Y));
KC_OAI211B_X1 T4597 ( .C0N(T16019_Y), .B(T4613_Y), .A(T4600_Y),     .C1(T4600_Y), .Y(T4597_Y));
KC_OAI211B_X1 T9268 ( .C0N(T9286_Y), .B(T7845_Y), .A(T9290_Y),     .C1(T161_Q), .Y(T9268_Y));
KC_OAI211B_X1 T4960 ( .C0N(T2671_Y), .B(T4939_Y), .A(T2190_Y),     .C1(T10959_Y), .Y(T4960_Y));
KC_OAI211B_X1 T5010 ( .C0N(T2815_Q), .B(T16156_Y), .A(T2276_Q),     .C1(T6070_Y), .Y(T5010_Y));
KC_OAI211B_X1 T5041 ( .C0N(T15559_Y), .B(T15562_Y), .A(T11989_Y),     .C1(T3210_Y), .Y(T5041_Y));
KC_OAI211B_X1 T5107 ( .C0N(T3825_Y), .B(T11377_Y), .A(T16153_Y),     .C1(T16154_Y), .Y(T5107_Y));
KC_OAI211B_X1 T5324 ( .C0N(T16462_Q), .B(T11252_Y), .A(T9972_Y),     .C1(T4934_Y), .Y(T5324_Y));
KC_OAI211B_X1 T5456 ( .C0N(T2762_Y), .B(T5941_Y), .A(T15928_Y),     .C1(T2734_Y), .Y(T5456_Y));
KC_OAI211B_X1 T5467 ( .C0N(T5457_Y), .B(T5470_Y), .A(T6284_Y),     .C1(T4557_Y), .Y(T5467_Y));
KC_OAI211B_X1 T5490 ( .C0N(T10973_Y), .B(T11666_Y), .A(T3369_Y),     .C1(T16057_Y), .Y(T5490_Y));
KC_OAI211B_X1 T5516 ( .C0N(T6568_S), .B(T11684_Y), .A(T4123_Y),     .C1(T11796_Y), .Y(T5516_Y));
KC_DFFRNHQ_X1 T964 ( .Q(T964_Q), .D(T962_Y), .RN(T15001_Y),     .CK(T971_Y));
KC_DFFRNHQ_X1 T1758 ( .Q(T1758_Q), .D(T1757_Y), .RN(T15011_Y),     .CK(T14554_Q));
KC_DFFRNHQ_X1 T2089 ( .Q(T2089_Q), .D(T15124_Y), .RN(T15008_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X1 T2091 ( .Q(T2091_Q), .D(T2090_Y), .RN(T15034_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X1 T2360 ( .Q(T2360_Q), .D(T12863_Y), .RN(T15037_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X1 T2361 ( .Q(T2361_Q), .D(T12469_Y), .RN(T15037_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X1 T2382 ( .Q(T2382_Q), .D(T2377_Y), .RN(T2709_Y),     .CK(T14560_Q));
KC_DFFRNHQ_X1 T2618 ( .Q(T2618_Q), .D(T15702_Y), .RN(T2063_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X1 T2640 ( .Q(T2640_Q), .D(T2641_Y), .RN(T2062_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X1 T2809 ( .Q(T2809_Q), .D(T11622_Y), .RN(T15020_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X1 T2844 ( .Q(T2844_Q), .D(T16053_Y), .RN(T15020_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X1 T4176 ( .Q(T4176_Q), .D(T8164_Y), .RN(T4047_Y),     .CK(T3496_Y));
KC_DFFRNHQ_X1 T4179 ( .Q(T4179_Q), .D(T11035_Y), .RN(T4047_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X1 T4538 ( .Q(T4538_Q), .D(T8263_Y), .RN(T3888_Y),     .CK(T14561_Q));
KC_DFFRNHQ_X1 T5380 ( .Q(T5380_Q), .D(T748_Y), .RN(T15001_Y),     .CK(T971_Y));
KC_DFFRNHQ_X1 T5480 ( .Q(T5480_Q), .D(T13156_Y), .RN(T15018_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X1 T5525 ( .Q(T5525_Q), .D(T11791_Y), .RN(T4047_Y),     .CK(T14575_Q));
KC_XOR2_X4 T2397 ( .A(T5640_Co), .B(T5586_Q), .Y(T2397_Y));
KC_XOR2_X4 T2312 ( .A(T8882_Y), .B(T8884_Y), .Y(T2312_Y));
KC_XOR2_X4 T2277 ( .A(T8842_Y), .B(T8788_Y), .Y(T2277_Y));
KC_XOR2_X4 T2242 ( .A(T8991_Y), .B(T11304_Y), .Y(T2242_Y));
KC_XOR2_X4 T2241 ( .A(T4807_Y), .B(T1445_Y), .Y(T2241_Y));
KC_XOR2_X4 T2130 ( .A(T239_Y), .B(T252_Y), .Y(T2130_Y));
KC_XOR2_X4 T2071 ( .A(T8969_Y), .B(T8957_Y), .Y(T2071_Y));
KC_XOR2_X4 T2049 ( .A(T5336_Y), .B(T15110_Y), .Y(T2049_Y));
KC_XOR2_X4 T1538 ( .A(T5284_Y), .B(T15098_Y), .Y(T1538_Y));
KC_XOR2_X4 T1523 ( .A(T9499_Y), .B(T9211_Y), .Y(T1523_Y));
KC_XOR2_X4 T1252 ( .A(T9249_Y), .B(T4816_Y), .Y(T1252_Y));
KC_XOR2_X4 T1167 ( .A(T9183_Y), .B(T9491_Y), .Y(T1167_Y));
KC_XOR2_X4 T1016 ( .A(T9492_Y), .B(T15095_Y), .Y(T1016_Y));
KC_XOR2_X4 T957 ( .A(T425_Y), .B(T9174_Y), .Y(T957_Y));
KC_XOR2_X4 T841 ( .A(T11303_Y), .B(T1345_Y), .Y(T841_Y));
KC_XOR2_X4 T776 ( .A(T11898_Y), .B(T12459_Y), .Y(T776_Y));
KC_XOR2_X4 T654 ( .A(T9201_Y), .B(T1354_Y), .Y(T654_Y));
KC_XOR2_X4 T620 ( .A(T9215_Y), .B(T9205_Y), .Y(T620_Y));
KC_XOR2_X4 T608 ( .A(T9217_Y), .B(T9218_Y), .Y(T608_Y));
KC_XOR2_X4 T591 ( .A(T9250_Y), .B(T9210_Y), .Y(T591_Y));
KC_XOR2_X4 T426 ( .A(T9202_Y), .B(T9208_Y), .Y(T426_Y));
KC_XOR2_X4 T425 ( .A(T9216_Y), .B(T9209_Y), .Y(T425_Y));
KC_XOR2_X4 T16516 ( .A(T9198_Y), .B(T9197_Y), .Y(T16516_Y));
KC_XOR2_X4 T16515 ( .A(T9159_Co), .B(T9472_Q), .Y(T16515_Y));
KC_XOR2_X4 T16514 ( .A(T15894_Q), .B(T15101_Y), .Y(T16514_Y));
KC_XOR2_X4 T16513 ( .A(T15894_Q), .B(T15102_Y), .Y(T16513_Y));
KC_XOR2_X4 T16512 ( .A(T7239_Y), .B(T15046_Y), .Y(T16512_Y));
KC_XOR2_X4 T16511 ( .A(T9466_Y), .B(T9225_S), .Y(T16511_Y));
KC_XOR2_X4 T16510 ( .A(T7088_Y), .B(T836_Y), .Y(T16510_Y));
KC_XOR2_X4 T16509 ( .A(T7870_Y), .B(T958_Y), .Y(T16509_Y));
KC_XOR2_X4 T16508 ( .A(T5417_Q), .B(T9188_Co), .Y(T16508_Y));
KC_XOR2_X4 T16507 ( .A(T15880_Q), .B(T15120_Y), .Y(T16507_Y));
KC_XOR2_X4 T16506 ( .A(T10127_Y), .B(T1268_Y), .Y(T16506_Y));
KC_XOR2_X4 T16505 ( .A(T13361_Q), .B(T16504_Y), .Y(T16505_Y));
KC_XOR2_X4 T16504 ( .A(T292_Y), .B(T6890_Y), .Y(T16504_Y));
KC_XOR2_X4 T4425 ( .A(T16461_Q), .B(T2055_Y), .Y(T4425_Y));
KC_XOR2_X4 T3342 ( .A(T15534_Y), .B(T10185_Y), .Y(T3342_Y));
KC_XOR2_X4 T3339 ( .A(T5070_Y), .B(T11489_Y), .Y(T3339_Y));
KC_XOR2_X4 T3338 ( .A(T11564_Y), .B(T12835_Y), .Y(T3338_Y));
KC_XOR2_X4 T3306 ( .A(T16008_Y), .B(T16009_Y), .Y(T3306_Y));
KC_XOR2_X4 T3304 ( .A(T5497_Q), .B(T12052_Y), .Y(T3304_Y));
KC_XOR2_X4 T3214 ( .A(T12315_Y), .B(T13170_Q), .Y(T3214_Y));
KC_XOR2_X4 T2960 ( .A(T5545_Y), .B(T6499_Y), .Y(T2960_Y));
KC_XOR2_X4 T2958 ( .A(T8159_Y), .B(T11839_Y), .Y(T2958_Y));
KC_XOR2_X4 T2957 ( .A(T9965_Y), .B(T2626_Q), .Y(T2957_Y));
KC_XOR2_X4 T2807 ( .A(T16068_Y), .B(T2639_Q), .Y(T2807_Y));
KC_XOR2_X4 T2788 ( .A(T15861_Y), .B(T12343_Y), .Y(T2788_Y));
KC_XOR2_X4 T2768 ( .A(T15930_Y), .B(T5016_Q), .Y(T2768_Y));
KC_XOR2_X4 T2765 ( .A(T14566_Q), .B(T12029_Y), .Y(T2765_Y));
KC_XOR2_X4 T4177 ( .A(T14563_Q), .B(T10641_Y), .Y(T4177_Y));
KC_XOR2_X4 T4174 ( .A(T13137_Y), .B(T11563_Y), .Y(T4174_Y));
KC_XOR2_X4 T4172 ( .A(T2798_Y), .B(T6776_S), .Y(T4172_Y));
KC_XOR2_X4 T4096 ( .A(T2836_Y), .B(T2955_Q), .Y(T4096_Y));
KC_XOR2_X4 T4055 ( .A(T6367_Y), .B(T2953_Q), .Y(T4055_Y));
KC_XOR2_X4 T4054 ( .A(T16473_Y), .B(T5541_Q), .Y(T4054_Y));
KC_XOR2_X4 T422 ( .A(T6413_Y), .B(T12944_Y), .Y(T422_Y));
KC_XOR2_X4 T3998 ( .A(T3219_Y), .B(T3206_Y), .Y(T3998_Y));
KC_XOR2_X4 T4384 ( .A(T11456_Y), .B(T3282_Y), .Y(T4384_Y));
KC_XOR2_X4 T3991 ( .A(T3291_Y), .B(T11515_Y), .Y(T3991_Y));
KC_XOR2_X4 T3921 ( .A(T11477_Y), .B(T11610_Y), .Y(T3921_Y));
KC_XOR2_X4 T3876 ( .A(T10637_Y), .B(T3337_Y), .Y(T3876_Y));
KC_XOR2_X4 T3451 ( .A(T15131_Y), .B(T11560_Y), .Y(T3451_Y));
KC_XOR2_X4 T3363 ( .A(T16001_Y), .B(T3316_Y), .Y(T3363_Y));
KC_XOR2_X4 T3344 ( .A(T3324_Y), .B(T3333_Y), .Y(T3344_Y));
KC_XOR2_X4 T16503 ( .A(T15984_Y), .B(T12244_Y), .Y(T16503_Y));
KC_XOR2_X4 T16502 ( .A(T12285_Y), .B(T15624_Y), .Y(T16502_Y));
KC_XOR2_X4 T421 ( .A(T11527_Y), .B(T4410_Y), .Y(T421_Y));
KC_XOR2_X4 T16501 ( .A(T6146_Co), .B(T5129_Q), .Y(T16501_Y));
KC_XOR2_X4 T16500 ( .A(T11483_Y), .B(T15581_Y), .Y(T16500_Y));
KC_XOR2_X4 T16417 ( .A(T8332_Y), .B(T13151_Q), .Y(T16417_Y));
KC_XOR2_X4 T16416 ( .A(T3990_Q), .B(T4591_Y), .Y(T16416_Y));
KC_XOR2_X4 T3281 ( .A(T13150_Q), .B(T11606_Y), .Y(T3281_Y));
KC_XOR2_X4 T4928 ( .A(T4037_Y), .B(T4069_Y), .Y(T4928_Y));
KC_XOR2_X4 T4748 ( .A(T5113_Y), .B(T4050_Q), .Y(T4748_Y));
KC_XOR2_X4 T4716 ( .A(T5504_Y), .B(T4691_Y), .Y(T4716_Y));
KC_XOR2_X4 T4662 ( .A(T4175_Y), .B(T3527_Y), .Y(T4662_Y));
KC_XOR2_X4 T4609 ( .A(T6611_Co), .B(T4169_Q), .Y(T4609_Y));
KC_XOR2_X4 T4540 ( .A(T6590_Co), .B(T4176_Q), .Y(T4540_Y));
KC_XOR2_X4 T420 ( .A(T4386_Y), .B(T5800_Y), .Y(T420_Y));
KC_XOR2_X4 T413 ( .A(T15156_Y), .B(T4455_Q), .Y(T413_Y));
KC_XOR2_X4 T4485 ( .A(T5761_Y), .B(T6027_Y), .Y(T4485_Y));
KC_XOR2_X4 T4483 ( .A(T8262_Y), .B(T15569_Y), .Y(T4483_Y));
KC_XOR2_X4 T16241 ( .A(T12151_Y), .B(T5165_Q), .Y(T16241_Y));
KC_XOR2_X4 T9487 ( .A(T3335_Y), .B(T4542_Y), .Y(T9487_Y));
KC_XOR2_X4 T9486 ( .A(T3982_Y), .B(T3942_Y), .Y(T9486_Y));
KC_XOR2_X4 T5466 ( .A(T5495_Q), .B(T15136_Y), .Y(T5466_Y));
KC_XOR2_X4 T5464 ( .A(T4721_Q), .B(T4712_Y), .Y(T5464_Y));
KC_XOR2_X4 T5339 ( .A(T4746_Q), .B(T12859_Y), .Y(T5339_Y));
KC_XOR2_X4 T5336 ( .A(T9493_Y), .B(T9248_Y), .Y(T5336_Y));
KC_XOR2_X4 T5284 ( .A(T9206_Y), .B(T9213_Y), .Y(T5284_Y));
KC_XOR2_X4 T5063 ( .A(T11552_Y), .B(T2370_Y), .Y(T5063_Y));
KC_XOR2_X4 T5021 ( .A(T12124_Y), .B(T3783_Y), .Y(T5021_Y));
KC_XOR2_X4 T5029 ( .A(T12460_Y), .B(T1_Y), .Y(T5029_Y));
KC_XOR2_X4 T16202 ( .A(T5061_Y), .B(T10642_Y), .Y(T16202_Y));
KC_XOR2_X4 T16201 ( .A(T3061_Y), .B(T2494_Y), .Y(T16201_Y));
KC_XOR2_X4 T15537 ( .A(T15927_Y), .B(T9923_Y), .Y(T15537_Y));
KC_XOR2_X4 T15328 ( .A(T7780_Y), .B(T7986_Y), .Y(T15328_Y));
KC_XOR2_X4 T5415 ( .A(T9237_Y), .B(T9204_Y), .Y(T5415_Y));
KC_XOR2_X4 T5414 ( .A(T1384_Y), .B(T10284_Y), .Y(T5414_Y));
KC_XOR2_X4 T5537 ( .A(T9482_Y), .B(T4916_Y), .Y(T5537_Y));
KC_XOR2_X4 T5484 ( .A(T3915_Y), .B(T5897_Y), .Y(T5484_Y));
KC_XOR2_X4 T5483 ( .A(T11490_Y), .B(T5895_Y), .Y(T5483_Y));
KC_XOR2_X4 T12843 ( .A(T4598_Y), .B(T4006_Q), .Y(T12843_Y));
KC_XOR2_X4 T7836 ( .A(T2951_Y), .B(T6539_Y), .Y(T7836_Y));
KC_OAI112B_X2 T16123 ( .C0(T955_Y), .B(T565_Y), .AN(T11273_Y),     .C1(T7872_Y), .Y(T16123_Y));
KC_OAI112B_X2 T16115 ( .C0(T910_Q), .B(T8725_Y), .AN(T7616_Y),     .C1(T15792_Y), .Y(T16115_Y));
KC_OAI112B_X2 T16117 ( .C0(T9915_Y), .B(T15466_Y), .AN(T9404_Y),     .C1(T1100_Q), .Y(T16117_Y));
KC_OAI112B_X2 T15830 ( .C0(T4992_Y), .B(T2693_Y), .AN(T11964_Y),     .C1(T14954_Q), .Y(T15830_Y));
KC_OAI112B_X2 T15834 ( .C0(T5772_Y), .B(T12139_Y), .AN(T3799_Y),     .C1(T5780_Y), .Y(T15834_Y));
KC_OAI112B_X2 T15955 ( .C0(T3917_Y), .B(T3907_Y), .AN(T13313_Y),     .C1(T3945_Y), .Y(T15955_Y));
KC_OAI112B_X2 T15899 ( .C0(T12798_Y), .B(T15898_Y), .AN(T11423_Y),     .C1(T4465_Q), .Y(T15899_Y));
KC_OAI112B_X2 T15838 ( .C0(T5770_Y), .B(T16154_Y), .AN(T15888_Y),     .C1(T11349_Y), .Y(T15838_Y));
KC_OAI112B_X2 T6528 ( .C0(T12467_Y), .B(T3518_Y), .AN(T12968_Y),     .C1(T2865_Y), .Y(T6528_Y));
KC_NAND2B_X1 T52 ( .B(T44_Q), .Y(T52_Y), .AN(T5220_Q));
KC_NAND2B_X1 T79 ( .B(T85_Q), .Y(T79_Y), .AN(T5187_Q));
KC_NAND2B_X1 T247 ( .B(T15490_Y), .Y(T247_Y), .AN(T15489_Y));
KC_NAND2B_X1 T349 ( .B(T9353_Q), .Y(T349_Y), .AN(T337_Q));
KC_NAND2B_X1 T378 ( .B(T8782_Y), .Y(T378_Y), .AN(T8747_Y));
KC_NAND2B_X1 T387 ( .B(T9449_Y), .Y(T387_Y), .AN(T9078_Y));
KC_NAND2B_X1 T419 ( .B(T9119_Y), .Y(T419_Y), .AN(T9125_Y));
KC_NAND2B_X1 T513 ( .B(T9378_Y), .Y(T513_Y), .AN(T722_Q));
KC_NAND2B_X1 T540 ( .B(T8838_Y), .Y(T540_Y), .AN(T8747_Y));
KC_NAND2B_X1 T558 ( .B(T8983_Y), .Y(T558_Y), .AN(T7829_Y));
KC_NAND2B_X1 T559 ( .B(T8119_Y), .Y(T559_Y), .AN(T8980_Y));
KC_NAND2B_X1 T597 ( .B(T11233_Y), .Y(T597_Y), .AN(T12447_Y));
KC_NAND2B_X1 T598 ( .B(T9065_Y), .Y(T598_Y), .AN(T4842_Y));
KC_NAND2B_X1 T667 ( .B(T7599_Y), .Y(T667_Y), .AN(T9373_Y));
KC_NAND2B_X1 T673 ( .B(T12395_Y), .Y(T673_Y), .AN(T6485_Y));
KC_NAND2B_X1 T720 ( .B(T757_Y), .Y(T720_Y), .AN(T756_Y));
KC_NAND2B_X1 T832 ( .B(T8630_Y), .Y(T832_Y), .AN(T12393_Y));
KC_NAND2B_X1 T833 ( .B(T4853_Y), .Y(T833_Y), .AN(T7088_Y));
KC_NAND2B_X1 T919 ( .B(T1724_Y), .Y(T919_Y), .AN(T9361_Y));
KC_NAND2B_X1 T952 ( .B(T8845_Y), .Y(T952_Y), .AN(T8799_Y));
KC_NAND2B_X1 T979 ( .B(T16420_Y), .Y(T979_Y), .AN(T952_Y));
KC_NAND2B_X1 T1039 ( .B(T1048_Q), .Y(T1039_Y), .AN(T15775_Y));
KC_NAND2B_X1 T1125 ( .B(T8032_Y), .Y(T1125_Y), .AN(T5376_Q));
KC_NAND2B_X1 T1772 ( .B(T2186_Q), .Y(T1772_Y), .AN(T1760_Q));
KC_NAND2B_X1 T2009 ( .B(T9968_Y), .Y(T2009_Y), .AN(T9882_Y));
KC_NAND2B_X1 T2020 ( .B(T2014_Y), .Y(T2020_Y), .AN(T1998_Y));
KC_NAND2B_X1 T2025 ( .B(T1119_Y), .Y(T2025_Y), .AN(T1107_Y));
KC_NAND2B_X1 T2048 ( .B(T16411_Y), .Y(T2048_Y), .AN(T9967_Y));
KC_NAND2B_X1 T2070 ( .B(T6593_Y), .Y(T2070_Y), .AN(T16234_Y));
KC_NAND2B_X1 T2110 ( .B(T2165_Y), .Y(T2110_Y), .AN(T11970_Y));
KC_NAND2B_X1 T2158 ( .B(T2145_Y), .Y(T2158_Y), .AN(T11436_Y));
KC_NAND2B_X1 T2175 ( .B(T1760_Q), .Y(T2175_Y), .AN(T2186_Q));
KC_NAND2B_X1 T2176 ( .B(T15974_Y), .Y(T2176_Y), .AN(T11500_Y));
KC_NAND2B_X1 T2185 ( .B(T15974_Y), .Y(T2185_Y), .AN(T11517_Y));
KC_NAND2B_X1 T2310 ( .B(T10612_Y), .Y(T2310_Y), .AN(T2311_Q));
KC_NAND2B_X1 T2362 ( .B(T2336_Y), .Y(T2362_Y), .AN(T11773_Y));
KC_NAND2B_X1 T2363 ( .B(T2336_Y), .Y(T2363_Y), .AN(T2373_Y));
KC_NAND2B_X1 T2383 ( .B(T2371_Y), .Y(T2383_Y), .AN(T2393_Y));
KC_NAND2B_X1 T2393 ( .B(T4963_Y), .Y(T2393_Y), .AN(T4979_Y));
KC_NAND2B_X1 T2496 ( .B(T1535_Y), .Y(T2496_Y), .AN(T3061_Y));
KC_NAND2B_X1 T2539 ( .B(T8453_Y), .Y(T2539_Y), .AN(T2541_Y));
KC_NAND2B_X1 T2540 ( .B(T1101_Y), .Y(T2540_Y), .AN(T881_Y));
KC_NAND2B_X1 T2641 ( .B(T2633_Y), .Y(T2641_Y), .AN(T2566_Y));
KC_NAND2B_X1 T2674 ( .B(T2677_Y), .Y(T2674_Y), .AN(T2676_Y));
KC_NAND2B_X1 T2698 ( .B(T15849_Y), .Y(T2698_Y), .AN(T14957_Q));
KC_NAND2B_X1 T2720 ( .B(T5860_Y), .Y(T2720_Y), .AN(T3257_Q));
KC_NAND2B_X1 T2784 ( .B(T6279_Y), .Y(T2784_Y), .AN(T2789_Y));
KC_NAND2B_X1 T2812 ( .B(T16024_Y), .Y(T2812_Y), .AN(T3423_Y));
KC_NAND2B_X1 T2836 ( .B(T2840_Y), .Y(T2836_Y), .AN(T12252_Y));
KC_NAND2B_X1 T2879 ( .B(T5567_Q), .Y(T2879_Y), .AN(T3214_Y));
KC_NAND2B_X1 T2926 ( .B(T2903_Y), .Y(T2926_Y), .AN(T2329_Y));
KC_NAND2B_X1 T2947 ( .B(T2933_Y), .Y(T2947_Y), .AN(T6516_Y));
KC_NAND2B_X1 T3076 ( .B(T3078_Y), .Y(T3076_Y), .AN(T3728_Y));
KC_NAND2B_X1 T3211 ( .B(T14949_Q), .Y(T3211_Y), .AN(T10266_Y));
KC_NAND2B_X1 T3212 ( .B(T12147_Y), .Y(T3212_Y), .AN(T12132_Y));
KC_NAND2B_X1 T3260 ( .B(T3250_Y), .Y(T3260_Y), .AN(T3266_Y));
KC_NAND2B_X1 T3261 ( .B(T5860_Y), .Y(T3261_Y), .AN(T13096_Q));
KC_NAND2B_X1 T3262 ( .B(T15129_Y), .Y(T3262_Y), .AN(T15929_Y));
KC_NAND2B_X1 T3270 ( .B(T3274_Y), .Y(T3270_Y), .AN(T3263_Y));
KC_NAND2B_X1 T3271 ( .B(T5860_Y), .Y(T3271_Y), .AN(T13110_Q));
KC_NAND2B_X1 T3275 ( .B(T5860_Y), .Y(T3275_Y), .AN(T13298_Q));
KC_NAND2B_X1 T3301 ( .B(T5860_Y), .Y(T3301_Y), .AN(T3256_Q));
KC_NAND2B_X1 T3302 ( .B(T5860_Y), .Y(T3302_Y), .AN(T12980_Q));
KC_NAND2B_X1 T3312 ( .B(T8267_Y), .Y(T3312_Y), .AN(T11486_Y));
KC_NAND2B_X1 T3313 ( .B(T5860_Y), .Y(T3313_Y), .AN(T5462_Q));
KC_NAND2B_X1 T3408 ( .B(T10585_Y), .Y(T3408_Y), .AN(T10970_Y));
KC_NAND2B_X1 T3455 ( .B(T3456_Y), .Y(T3455_Y), .AN(T3428_Y));
KC_NAND2B_X1 T3458 ( .B(T3435_Y), .Y(T3458_Y), .AN(T3389_Y));
KC_NAND2B_X1 T3497 ( .B(T3474_Y), .Y(T3497_Y), .AN(T10554_Y));
KC_NAND2B_X1 T3526 ( .B(T11832_Y), .Y(T3526_Y), .AN(T3508_Y));
KC_NAND2B_X1 T3818 ( .B(T11984_Y), .Y(T3818_Y), .AN(T3831_Y));
KC_NAND2B_X1 T3880 ( .B(T11414_Y), .Y(T3880_Y), .AN(T2700_Y));
KC_NAND2B_X1 T3930 ( .B(T15961_Y), .Y(T3930_Y), .AN(T11023_Y));
KC_NAND2B_X1 T3931 ( .B(T11590_Y), .Y(T3931_Y), .AN(T3906_Y));
KC_NAND2B_X1 T3932 ( .B(T3933_Y), .Y(T3932_Y), .AN(T5120_Y));
KC_NAND2B_X1 T3933 ( .B(T10937_Y), .Y(T3933_Y), .AN(T3966_Y));
KC_NAND2B_X1 T3960 ( .B(T5985_Y), .Y(T3960_Y), .AN(T12164_Y));
KC_NAND2B_X1 T3983 ( .B(T5860_Y), .Y(T3983_Y), .AN(T3281_Y));
KC_NAND2B_X1 T3985 ( .B(T5860_Y), .Y(T3985_Y), .AN(T5479_Q));
KC_NAND2B_X1 T3986 ( .B(T5860_Y), .Y(T3986_Y), .AN(T12843_Y));
KC_NAND2B_X1 T3987 ( .B(T5860_Y), .Y(T3987_Y), .AN(T13154_Q));
KC_NAND2B_X1 T4009 ( .B(T12957_Y), .Y(T4009_Y), .AN(T5992_Y));
KC_NAND2B_X1 T4049 ( .B(T11626_Y), .Y(T4049_Y), .AN(T3354_Y));
KC_NAND2B_X1 T4099 ( .B(T11745_Y), .Y(T4099_Y), .AN(T4070_Y));
KC_NAND2B_X1 T4101 ( .B(T10580_Y), .Y(T4101_Y), .AN(T10577_Y));
KC_NAND2B_X1 T4104 ( .B(T11636_Y), .Y(T4104_Y), .AN(T2849_Y));
KC_NAND2B_X1 T4146 ( .B(T5522_Y), .Y(T4146_Y), .AN(T12041_Y));
KC_NAND2B_X1 T4149 ( .B(T4140_Y), .Y(T4149_Y), .AN(T13179_Y));
KC_NAND2B_X1 T4180 ( .B(T3996_Y), .Y(T4180_Y), .AN(T4761_Y));
KC_NAND2B_X1 T4284 ( .B(T4272_Y), .Y(T4284_Y), .AN(T15782_Y));
KC_NAND2B_X1 T4494 ( .B(T4481_Y), .Y(T4494_Y), .AN(T15934_Y));
KC_NAND2B_X1 T4503 ( .B(T4480_Y), .Y(T4503_Y), .AN(T4502_Y));
KC_NAND2B_X1 T4532 ( .B(T4518_Y), .Y(T4532_Y), .AN(T10925_Y));
KC_NAND2B_X1 T4599 ( .B(T4582_Y), .Y(T4599_Y), .AN(T6010_Y));
KC_NAND2B_X1 T4614 ( .B(T4615_Y), .Y(T4614_Y), .AN(T5485_Y));
KC_NAND2B_X1 T4664 ( .B(T6467_Y), .Y(T4664_Y), .AN(T11706_Y));
KC_NAND2B_X1 T4687 ( .B(T4665_Y), .Y(T4687_Y), .AN(T4690_Y));
KC_NAND2B_X1 T4751 ( .B(T4752_Y), .Y(T4751_Y), .AN(T13184_Y));
KC_NAND2B_X1 T4850 ( .B(T15485_Y), .Y(T4850_Y), .AN(T15660_Y));
KC_NAND2B_X1 T4919 ( .B(T10757_Y), .Y(T4919_Y), .AN(T16468_Q));
KC_NAND2B_X1 T4931 ( .B(T6737_Y), .Y(T4931_Y), .AN(T2133_Y));
KC_NAND2B_X1 T4978 ( .B(T8427_Y), .Y(T4978_Y), .AN(T4963_Y));
KC_NAND2B_X1 T5017 ( .B(T5860_Y), .Y(T5017_Y), .AN(T13299_Q));
KC_NAND2B_X1 T5019 ( .B(T10280_Y), .Y(T5019_Y), .AN(T2664_Y));
KC_NAND2B_X1 T5065 ( .B(T8486_Y), .Y(T5065_Y), .AN(T8488_Y));
KC_NAND2B_X1 T5077 ( .B(T10266_Y), .Y(T5077_Y), .AN(T14949_Q));
KC_NAND2B_X1 T5122 ( .B(T15878_Y), .Y(T5122_Y), .AN(T5472_Y));
KC_NAND2B_X1 T5124 ( .B(T12349_Y), .Y(T5124_Y), .AN(T12349_Y));
KC_NAND2B_X1 T5433 ( .B(T15833_Y), .Y(T5433_Y), .AN(T3791_Y));
KC_NAND2B_X1 T5450 ( .B(T5860_Y), .Y(T5450_Y), .AN(T5451_Q));
KC_NAND2B_X1 T5472 ( .B(T5860_Y), .Y(T5472_Y), .AN(T13119_Q));
KC_NAND2B_X1 T5535 ( .B(T11844_Y), .Y(T5535_Y), .AN(T8160_Y));
KC_NAND2B_X1 T5539 ( .B(T11843_Y), .Y(T5539_Y), .AN(T3513_Y));
KC_NAND2B_X1 T5545 ( .B(T1844_Y), .Y(T5545_Y), .AN(T1843_Y));
KC_BUF_X3 T18 ( .Y(T18_Y), .A(T1243_Y));
KC_BUF_X3 T19 ( .Y(T19_Y), .A(T2380_Y));
KC_BUF_X3 T20 ( .Y(T20_Y), .A(T4187_Y));
KC_BUF_X3 T1006 ( .Y(T1006_Y), .A(T974_Q));
KC_BUF_X3 T1024 ( .Y(T1024_Y), .A(T16168_Y));
KC_BUF_X3 T1169 ( .Y(T1169_Y), .A(T1753_Q));
KC_BUF_X3 T1170 ( .Y(T1170_Y), .A(T14965_Y));
KC_BUF_X3 T1244 ( .Y(T1244_Y), .A(T15230_Y));
KC_BUF_X3 T1616 ( .Y(T1616_Y), .A(T15924_Y));
KC_BUF_X3 T1745 ( .Y(T1745_Y), .A(T13108_Q));
KC_BUF_X3 T1746 ( .Y(T1746_Y), .A(T4930_Q));
KC_BUF_X3 T1755 ( .Y(T1755_Y), .A(T2153_Q));
KC_BUF_X3 T1756 ( .Y(T1756_Y), .A(T2129_Q));
KC_BUF_X3 T1850 ( .Y(T1850_Y), .A(T1846_Y));
KC_BUF_X3 T1835 ( .Y(T1835_Y), .A(T1835_A));
KC_BUF_X3 T1848 ( .Y(T1848_Y), .A(T1831_Y));
KC_BUF_X3 T1849 ( .Y(T1849_Y), .A(T1831_Y));
KC_BUF_X3 T2081 ( .Y(T2081_Y), .A(T15230_Y));
KC_BUF_X3 T2379 ( .Y(T2379_Y), .A(T2384_Y));
KC_BUF_X3 T2380 ( .Y(T2380_Y), .A(T2342_Y));
KC_BUF_X3 T2401 ( .Y(T2401_Y), .A(T15019_Y));
KC_BUF_X3 T2709 ( .Y(T2709_Y), .A(T2081_Y));
KC_BUF_X3 T4186 ( .Y(T4186_Y), .A(T4784_Y));
KC_BUF_X3 T4187 ( .Y(T4187_Y), .A(T18_Y));
KC_BUF_X3 T4783 ( .Y(T4783_Y), .A(T2379_Y));
KC_BUF_X3 T4784 ( .Y(T4784_Y), .A(T3999_Y));
KC_BUF_X3 T5443 ( .Y(T5443_Y), .A(T1759_Q));
KC_BUF_X3 T5547 ( .Y(T5547_Y), .A(T2248_Y));
KC_OAI112BB_X1 T15818 ( .B(T11961_Y), .AN(T2660_Y), .C0N(T11337_Y),     .C1(T3204_Y), .Y(T15818_Y));
KC_OAI21_X2 T15737 ( .B(T7553_Y), .A0(T11872_Y), .A1(T886_Y),     .Y(T15737_Y));
KC_OAI21_X2 T15310 ( .B(T7437_Y), .A0(T13239_Y), .A1(T886_Y),     .Y(T15310_Y));
KC_OAI21_X2 T6828 ( .B(T7363_Y), .A0(T11139_Y), .A1(T886_Y),     .Y(T6828_Y));
KC_OAI21_X2 T16116 ( .B(T7561_Y), .A0(T11199_Y), .A1(T886_Y),     .Y(T16116_Y));
KC_OAI21_X2 T8389 ( .B(T7560_Y), .A0(T11192_Y), .A1(T886_Y),     .Y(T8389_Y));
KC_OAI21_X2 T8384 ( .B(T7683_Y), .A0(T11197_Y), .A1(T886_Y),     .Y(T8384_Y));
KC_OAI21_X2 T16127 ( .B(T10596_Y), .A0(T12067_Y), .A1(T2867_Y),     .Y(T16127_Y));
KC_OAI21_X2 T15878 ( .B(T5860_Y), .A0(T3200_Y), .A1(T12148_Y),     .Y(T15878_Y));
KC_OAI21_X2 T16448 ( .B(T16451_Y), .A0(T2632_Y), .A1(T10934_Y),     .Y(T16448_Y));
KC_OAI21_X2 T6829 ( .B(T7415_Y), .A0(T11143_Y), .A1(T886_Y),     .Y(T6829_Y));
KC_OAI21_X2 T16449 ( .B(T16450_Y), .A0(T2632_Y), .A1(T13121_Y),     .Y(T16449_Y));
KC_OAI21_X1 T87 ( .B(T5633_Y), .A0(T98_Q), .A1(T8564_Y), .Y(T87_Y));
KC_OAI21_X1 T243 ( .B(T11296_Y), .A0(T9078_Y), .A1(T16285_Y),     .Y(T243_Y));
KC_OAI21_X1 T248 ( .B(T8960_Y), .A0(T1386_Y), .A1(T8993_Co),     .Y(T248_Y));
KC_OAI21_X1 T253 ( .B(T9203_Y), .A0(T1353_Y), .A1(T8142_Y),     .Y(T253_Y));
KC_OAI21_X1 T297 ( .B(T9266_Y), .A0(T288_Q), .A1(T265_Y), .Y(T297_Y));
KC_OAI21_X1 T300 ( .B(T9260_Y), .A0(T306_Q), .A1(T332_Y), .Y(T300_Y));
KC_OAI21_X1 T303 ( .B(T7084_Y), .A0(T313_Q), .A1(T318_Y), .Y(T303_Y));
KC_OAI21_X1 T307 ( .B(T7104_Y), .A0(T275_Q), .A1(T321_Y), .Y(T307_Y));
KC_OAI21_X1 T308 ( .B(T7121_Y), .A0(T158_Q), .A1(T348_Y), .Y(T308_Y));
KC_OAI21_X1 T340 ( .B(T8667_Y), .A0(T9353_Q), .A1(T569_Y), .Y(T340_Y));
KC_OAI21_X1 T388 ( .B(T4820_Y), .A0(T1440_Y), .A1(T1438_Y),     .Y(T388_Y));
KC_OAI21_X1 T415 ( .B(T9136_Y), .A0(T4817_Y), .A1(T9124_Y),     .Y(T415_Y));
KC_OAI21_X1 T476 ( .B(T7097_Y), .A0(T460_Q), .A1(T347_Y), .Y(T476_Y));
KC_OAI21_X1 T486 ( .B(T7306_Y), .A0(T5265_Q), .A1(T6348_Y),     .Y(T486_Y));
KC_OAI21_X1 T516 ( .B(T13260_Y), .A0(T543_Q), .A1(T517_Q), .Y(T516_Y));
KC_OAI21_X1 T518 ( .B(T8803_Y), .A0(T551_Q), .A1(T5356_Q), .Y(T518_Y));
KC_OAI21_X1 T555 ( .B(T8125_Y), .A0(T567_Q), .A1(T1593_Y), .Y(T555_Y));
KC_OAI21_X1 T571 ( .B(T12458_Y), .A0(T8079_Y), .A1(T1214_Y),     .Y(T571_Y));
KC_OAI21_X1 T592 ( .B(T1839_Y), .A0(T604_Q), .A1(T1593_Y), .Y(T592_Y));
KC_OAI21_X1 T599 ( .B(T955_Y), .A0(T10140_Y), .A1(T1593_Y),     .Y(T599_Y));
KC_OAI21_X1 T603 ( .B(T955_Y), .A0(T1593_Y), .A1(T9065_Y), .Y(T603_Y));
KC_OAI21_X1 T614 ( .B(T15538_Y), .A0(T168_Y), .A1(T9194_Y),     .Y(T614_Y));
KC_OAI21_X1 T691 ( .B(T8851_Y), .A0(T669_Q), .A1(T9314_Y), .Y(T691_Y));
KC_OAI21_X1 T16427 ( .B(T16354_Y), .A0(T9409_Y), .A1(T7892_Y),     .Y(T16427_Y));
KC_OAI21_X1 T16426 ( .B(T16356_Y), .A0(T9410_Y), .A1(T7892_Y),     .Y(T16426_Y));
KC_OAI21_X1 T16425 ( .B(T7887_Y), .A0(T9412_Y), .A1(T7892_Y),     .Y(T16425_Y));
KC_OAI21_X1 T721 ( .B(T7885_Y), .A0(T9408_Y), .A1(T7892_Y),     .Y(T721_Y));
KC_OAI21_X1 T732 ( .B(T7888_Y), .A0(T8893_Y), .A1(T7892_Y),     .Y(T732_Y));
KC_OAI21_X1 T733 ( .B(T7884_Y), .A0(T8802_Y), .A1(T7892_Y),     .Y(T733_Y));
KC_OAI21_X1 T734 ( .B(T7882_Y), .A0(T8851_Y), .A1(T7892_Y),     .Y(T734_Y));
KC_OAI21_X1 T735 ( .B(T7886_Y), .A0(T8853_Y), .A1(T7892_Y),     .Y(T735_Y));
KC_OAI21_X1 T909 ( .B(T755_Y), .A0(T8748_Y), .A1(T744_Y), .Y(T909_Y));
KC_OAI21_X1 T922 ( .B(T7618_Y), .A0(T7629_Y), .A1(T7617_Y),     .Y(T922_Y));
KC_OAI21_X1 T937 ( .B(T15454_Y), .A0(T16149_Y), .A1(T953_Y),     .Y(T937_Y));
KC_OAI21_X1 T953 ( .B(T15223_Y), .A0(T7839_Y), .A1(T12612_Y),     .Y(T953_Y));
KC_OAI21_X1 T989 ( .B(T10027_Y), .A0(T941_Y), .A1(T8849_Y),     .Y(T989_Y));
KC_OAI21_X1 T1010 ( .B(T972_Y), .A0(T9436_Y), .A1(T10142_Y),     .Y(T1010_Y));
KC_OAI21_X1 T1034 ( .B(T585_Y), .A0(T11880_Y), .A1(T6822_Y),     .Y(T1034_Y));
KC_OAI21_X1 T6796 ( .B(T585_Y), .A0(T11918_Y), .A1(T6822_Y),     .Y(T6796_Y));
KC_OAI21_X1 T1043 ( .B(T9723_Y), .A0(T5359_Q), .A1(T11087_Y),     .Y(T1043_Y));
KC_OAI21_X1 T1049 ( .B(T585_Y), .A0(T515_Y), .A1(T6822_Y),     .Y(T1049_Y));
KC_OAI21_X1 T1052 ( .B(T498_Y), .A0(T12400_Y), .A1(T7499_Y),     .Y(T1052_Y));
KC_OAI21_X1 T1053 ( .B(T585_Y), .A0(T8724_Y), .A1(T6822_Y),     .Y(T1053_Y));
KC_OAI21_X1 T1056 ( .B(T585_Y), .A0(T514_Y), .A1(T6822_Y),     .Y(T1056_Y));
KC_OAI21_X1 T1063 ( .B(T8029_Y), .A0(T1113_Q), .A1(T7976_Y),     .Y(T1063_Y));
KC_OAI21_X1 T1075 ( .B(T8029_Y), .A0(T1128_Q), .A1(T7976_Y),     .Y(T1075_Y));
KC_OAI21_X1 T16431 ( .B(T7845_Y), .A0(T7844_Y), .A1(T378_Y),     .Y(T16431_Y));
KC_OAI21_X1 T1087 ( .B(T8029_Y), .A0(T5334_Q), .A1(T7976_Y),     .Y(T1087_Y));
KC_OAI21_X1 T1090 ( .B(T7845_Y), .A0(T7844_Y), .A1(T540_Y),     .Y(T1090_Y));
KC_OAI21_X1 T1099 ( .B(T7845_Y), .A0(T7844_Y), .A1(T1062_Y),     .Y(T1099_Y));
KC_OAI21_X1 T1104 ( .B(T7845_Y), .A0(T7844_Y), .A1(T1042_Y),     .Y(T1104_Y));
KC_OAI21_X1 T16309 ( .B(T9986_Y), .A0(T1134_Y), .A1(T8110_Y),     .Y(T16309_Y));
KC_OAI21_X1 T1126 ( .B(T10660_Y), .A0(T927_Y), .A1(T1481_Y),     .Y(T1126_Y));
KC_OAI21_X1 T1144 ( .B(T1342_Y), .A0(T5353_Q), .A1(T9400_Y),     .Y(T1144_Y));
KC_OAI21_X1 T1150 ( .B(T972_Y), .A0(T10301_Y), .A1(T10142_Y),     .Y(T1150_Y));
KC_OAI21_X1 T1168 ( .B(T12114_Y), .A0(T1174_Y), .A1(T15798_Q),     .Y(T1168_Y));
KC_OAI21_X1 T1193 ( .B(T10040_Y), .A0(T1094_Q), .A1(T5337_Q),     .Y(T1193_Y));
KC_OAI21_X1 T1218 ( .B(T10024_Y), .A0(T1113_Q), .A1(T5341_Q),     .Y(T1218_Y));
KC_OAI21_X1 T1237 ( .B(T10024_Y), .A0(T1129_Q), .A1(T1223_Q),     .Y(T1237_Y));
KC_OAI21_X1 T1238 ( .B(T10040_Y), .A0(T5373_Q), .A1(T1232_Q),     .Y(T1238_Y));
KC_OAI21_X1 T1239 ( .B(T10048_Y), .A0(T10170_Y), .A1(T10021_Y),     .Y(T1239_Y));
KC_OAI21_X1 T1257 ( .B(T10157_Y), .A0(T15529_Y), .A1(T4838_Y),     .Y(T1257_Y));
KC_OAI21_X1 T6836 ( .B(T1453_Y), .A0(T7490_Y), .A1(T9720_Y),     .Y(T6836_Y));
KC_OAI21_X1 T1347 ( .B(T1453_Y), .A0(T7541_Y), .A1(T7490_Y),     .Y(T1347_Y));
KC_OAI21_X1 T1348 ( .B(T4885_Y), .A0(T7542_Y), .A1(T9720_Y),     .Y(T1348_Y));
KC_OAI21_X1 T1401 ( .B(T1419_Y), .A0(T10389_Y), .A1(T10380_Y),     .Y(T1401_Y));
KC_OAI21_X1 T6442 ( .B(T1418_Y), .A0(T6993_Y), .A1(T6982_Y),     .Y(T6442_Y));
KC_OAI21_X1 T6441 ( .B(T1418_Y), .A0(T6991_Y), .A1(T9542_Y),     .Y(T6441_Y));
KC_OAI21_X1 T1404 ( .B(T1418_Y), .A0(T6983_Y), .A1(T6982_Y),     .Y(T1404_Y));
KC_OAI21_X1 T1406 ( .B(T1418_Y), .A0(T6982_Y), .A1(T9543_Y),     .Y(T1406_Y));
KC_OAI21_X1 T1407 ( .B(T1418_Y), .A0(T6993_Y), .A1(T6991_Y),     .Y(T1407_Y));
KC_OAI21_X1 T1408 ( .B(T1418_Y), .A0(T6991_Y), .A1(T9543_Y),     .Y(T1408_Y));
KC_OAI21_X1 T1409 ( .B(T1418_Y), .A0(T6983_Y), .A1(T6991_Y),     .Y(T1409_Y));
KC_OAI21_X1 T1410 ( .B(T1418_Y), .A0(T6982_Y), .A1(T9542_Y),     .Y(T1410_Y));
KC_OAI21_X1 T6823 ( .B(T1453_Y), .A0(T7490_Y), .A1(T9721_Y),     .Y(T6823_Y));
KC_OAI21_X1 T1451 ( .B(T1453_Y), .A0(T7542_Y), .A1(T9721_Y),     .Y(T1451_Y));
KC_OAI21_X1 T1452 ( .B(T1453_Y), .A0(T7489_Y), .A1(T7542_Y),     .Y(T1452_Y));
KC_OAI21_X1 T1459 ( .B(T1492_Y), .A0(T7782_Y), .A1(T9810_Y),     .Y(T1459_Y));
KC_OAI21_X1 T16307 ( .B(T1493_Y), .A0(T10016_Y), .A1(T10014_Y),     .Y(T16307_Y));
KC_OAI21_X1 T16298 ( .B(T1493_Y), .A0(T9995_Y), .A1(T10014_Y),     .Y(T16298_Y));
KC_OAI21_X1 T1500 ( .B(T1493_Y), .A0(T10016_Y), .A1(T10015_Y),     .Y(T1500_Y));
KC_OAI21_X1 T1501 ( .B(T1493_Y), .A0(T10018_Y), .A1(T10016_Y),     .Y(T1501_Y));
KC_OAI21_X1 T1502 ( .B(T1493_Y), .A0(T10017_Y), .A1(T10016_Y),     .Y(T1502_Y));
KC_OAI21_X1 T1503 ( .B(T1493_Y), .A0(T10018_Y), .A1(T9995_Y),     .Y(T1503_Y));
KC_OAI21_X1 T1504 ( .B(T1493_Y), .A0(T10017_Y), .A1(T9995_Y),     .Y(T1504_Y));
KC_OAI21_X1 T1507 ( .B(T1493_Y), .A0(T9995_Y), .A1(T10015_Y),     .Y(T1507_Y));
KC_OAI21_X1 T1520 ( .B(T1419_Y), .A0(T6990_Y), .A1(T9540_Y),     .Y(T1520_Y));
KC_OAI21_X1 T6439 ( .B(T1419_Y), .A0(T6990_Y), .A1(T9541_Y),     .Y(T6439_Y));
KC_OAI21_X1 T1526 ( .B(T1419_Y), .A0(T10389_Y), .A1(T6990_Y),     .Y(T1526_Y));
KC_OAI21_X1 T16179 ( .B(T1492_Y), .A0(T7705_Y), .A1(T9787_Y),     .Y(T16179_Y));
KC_OAI21_X1 T1552 ( .B(T1492_Y), .A0(T7782_Y), .A1(T9787_Y),     .Y(T1552_Y));
KC_OAI21_X1 T1553 ( .B(T1492_Y), .A0(T7781_Y), .A1(T7705_Y),     .Y(T1553_Y));
KC_OAI21_X1 T1556 ( .B(T1492_Y), .A0(T7704_Y), .A1(T7782_Y),     .Y(T1556_Y));
KC_OAI21_X1 T1557 ( .B(T1492_Y), .A0(T7704_Y), .A1(T7705_Y),     .Y(T1557_Y));
KC_OAI21_X1 T1559 ( .B(T1492_Y), .A0(T7781_Y), .A1(T7782_Y),     .Y(T1559_Y));
KC_OAI21_X1 T15883 ( .B(T2722_Y), .A0(T15916_Y), .A1(T15858_Y),     .Y(T15883_Y));
KC_OAI21_X1 T1757 ( .B(T2722_Y), .A0(T15916_Y), .A1(T15857_Y),     .Y(T1757_Y));
KC_OAI21_X1 T1776 ( .B(T10947_Y), .A0(T94_Y), .A1(T15974_Y),     .Y(T1776_Y));
KC_OAI21_X1 T1843 ( .B(T6494_Y), .A0(T1834_Y), .A1(T1834_Y),     .Y(T1843_Y));
KC_OAI21_X1 T1844 ( .B(T2400_Y), .A0(T6494_Y), .A1(T6496_Y),     .Y(T1844_Y));
KC_OAI21_X1 T2010 ( .B(T12097_Y), .A0(T2009_Y), .A1(T5369_Y),     .Y(T2010_Y));
KC_OAI21_X1 T2017 ( .B(T1992_Y), .A0(T1118_Y), .A1(T1142_Y),     .Y(T2017_Y));
KC_OAI21_X1 T2056 ( .B(T4936_Y), .A0(T16269_Y), .A1(T1509_Y),     .Y(T2056_Y));
KC_OAI21_X1 T2057 ( .B(T16305_Y), .A0(T1485_Y), .A1(T16411_Y),     .Y(T2057_Y));
KC_OAI21_X1 T15850 ( .B(T5436_Y), .A0(T15916_Y), .A1(T10245_Y),     .Y(T15850_Y));
KC_OAI21_X1 T2088 ( .B(T4943_Y), .A0(T15916_Y), .A1(T15912_Y),     .Y(T2088_Y));
KC_OAI21_X1 T2090 ( .B(T2132_Y), .A0(T15916_Y), .A1(T15855_Y),     .Y(T2090_Y));
KC_OAI21_X1 T2092 ( .B(T2104_Y), .A0(T15916_Y), .A1(T2719_Y),     .Y(T2092_Y));
KC_OAI21_X1 T2093 ( .B(T2104_Y), .A0(T15916_Y), .A1(T2127_Y),     .Y(T2093_Y));
KC_OAI21_X1 T2094 ( .B(T5436_Y), .A0(T15916_Y), .A1(T15853_Y),     .Y(T2094_Y));
KC_OAI21_X1 T2096 ( .B(T2132_Y), .A0(T15916_Y), .A1(T1748_Y),     .Y(T2096_Y));
KC_OAI21_X1 T2116 ( .B(T2165_Y), .A0(T15916_Y), .A1(T15895_Y),     .Y(T2116_Y));
KC_OAI21_X1 T2120 ( .B(T2140_Y), .A0(T15916_Y), .A1(T16474_Y),     .Y(T2120_Y));
KC_OAI21_X1 T2123 ( .B(T4943_Y), .A0(T15916_Y), .A1(T2751_Y),     .Y(T2123_Y));
KC_OAI21_X1 T2126 ( .B(T2145_Y), .A0(T15916_Y), .A1(T15854_Y),     .Y(T2126_Y));
KC_OAI21_X1 T2154 ( .B(T15943_Y), .A0(T10933_Y), .A1(T2168_Y),     .Y(T2154_Y));
KC_OAI21_X1 T2155 ( .B(T15942_Y), .A0(T5058_Y), .A1(T15574_Y),     .Y(T2155_Y));
KC_OAI21_X1 T2159 ( .B(T2140_Y), .A0(T15916_Y), .A1(T15856_Y),     .Y(T2159_Y));
KC_OAI21_X1 T2212 ( .B(T2802_Y), .A0(T16098_Y), .A1(T2217_Y),     .Y(T2212_Y));
KC_OAI21_X1 T2238 ( .B(T10959_Y), .A0(T2236_Q), .A1(T2217_Y),     .Y(T2238_Y));
KC_OAI21_X1 T2251 ( .B(T6070_Y), .A0(T12958_Y), .A1(T11599_Y),     .Y(T2251_Y));
KC_OAI21_X1 T2348 ( .B(T2349_Y), .A0(T16129_Y), .A1(T15713_Y),     .Y(T2348_Y));
KC_OAI21_X1 T2357 ( .B(T5520_Y), .A0(T5517_Y), .A1(T2325_Y),     .Y(T2357_Y));
KC_OAI21_X1 T2530 ( .B(T5979_Y), .A0(T16267_Y), .A1(T9849_Y),     .Y(T2530_Y));
KC_OAI21_X1 T2534 ( .B(T5979_Y), .A0(T2068_Y), .A1(T9849_Y),     .Y(T2534_Y));
KC_OAI21_X1 T2577 ( .B(T5869_S), .A0(T2573_Y), .A1(T9971_Y),     .Y(T2577_Y));
KC_OAI21_X1 T16293 ( .B(T5389_Q), .A0(T2575_Q), .A1(T15518_Y),     .Y(T16293_Y));
KC_OAI21_X1 T2621 ( .B(T10091_Y), .A0(T2360_Q), .A1(T12091_Y),     .Y(T2621_Y));
KC_OAI21_X1 T2622 ( .B(T10091_Y), .A0(T2361_Q), .A1(T12091_Y),     .Y(T2622_Y));
KC_OAI21_X1 T2624 ( .B(T15518_Y), .A0(T2844_Q), .A1(T10104_Y),     .Y(T2624_Y));
KC_OAI21_X1 T2629 ( .B(T16411_Y), .A0(T16367_Y), .A1(T1987_Y),     .Y(T2629_Y));
KC_OAI21_X1 T2643 ( .B(T15535_Y), .A0(T5408_Q), .A1(T5409_Y),     .Y(T2643_Y));
KC_OAI21_X1 T2648 ( .B(T5979_Y), .A0(T4896_Y), .A1(T2065_Y),     .Y(T2648_Y));
KC_OAI21_X1 T2666 ( .B(T14954_Q), .A0(T10271_Y), .A1(T10242_Y),     .Y(T2666_Y));
KC_OAI21_X1 T2690 ( .B(T10272_Y), .A0(T6061_Y), .A1(T2683_Y),     .Y(T2690_Y));
KC_OAI21_X1 T2691 ( .B(T2681_Y), .A0(T11357_Y), .A1(T5758_Y),     .Y(T2691_Y));
KC_OAI21_X1 T2694 ( .B(T4995_Y), .A0(T2683_Y), .A1(T8441_Y),     .Y(T2694_Y));
KC_OAI21_X1 T2696 ( .B(T15696_Y), .A0(T15752_Y), .A1(T14954_Q),     .Y(T2696_Y));
KC_OAI21_X1 T2697 ( .B(T12136_Y), .A0(T5766_Y), .A1(T2677_Y),     .Y(T2697_Y));
KC_OAI21_X1 T2742 ( .B(T8209_Y), .A0(T2751_Y), .A1(T13110_Q),     .Y(T2742_Y));
KC_OAI21_X1 T2743 ( .B(T11462_Y), .A0(T2281_Q), .A1(T8238_Y),     .Y(T2743_Y));
KC_OAI21_X1 T2745 ( .B(T11461_Y), .A0(T2249_Q), .A1(T8238_Y),     .Y(T2745_Y));
KC_OAI21_X1 T2750 ( .B(T5861_Y), .A0(T3283_Y), .A1(T6133_S),     .Y(T2750_Y));
KC_OAI21_X1 T2792 ( .B(T10959_Y), .A0(T5987_Q), .A1(T2217_Y),     .Y(T2792_Y));
KC_OAI21_X1 T2847 ( .B(T8503_Y), .A0(T3399_Y), .A1(T12831_Y),     .Y(T2847_Y));
KC_OAI21_X1 T2873 ( .B(T6183_Y), .A0(T2876_Y), .A1(T10592_Y),     .Y(T2873_Y));
KC_OAI21_X1 T2875 ( .B(T6583_Y), .A0(T3429_Y), .A1(T6180_Y),     .Y(T2875_Y));
KC_OAI21_X1 T2920 ( .B(T12306_Y), .A0(T8261_Y), .A1(T11808_Y),     .Y(T2920_Y));
KC_OAI21_X1 T2921 ( .B(T12312_Y), .A0(T16099_Y), .A1(T2908_Y),     .Y(T2921_Y));
KC_OAI21_X1 T2922 ( .B(T6196_Y), .A0(T2891_Y), .A1(T2889_Y),     .Y(T2922_Y));
KC_OAI21_X1 T2923 ( .B(T2898_Y), .A0(T15953_Y), .A1(T6240_Y),     .Y(T2923_Y));
KC_OAI21_X1 T2924 ( .B(T2896_Y), .A0(T11810_Y), .A1(T15633_Y),     .Y(T2924_Y));
KC_OAI21_X1 T2925 ( .B(T5521_Y), .A0(T6240_Y), .A1(T6583_Y),     .Y(T2925_Y));
KC_OAI21_X1 T2928 ( .B(T6196_Y), .A0(T10987_Y), .A1(T11767_Y),     .Y(T2928_Y));
KC_OAI21_X1 T8153 ( .B(T2950_Y), .A0(T11005_Y), .A1(T3509_Y),     .Y(T8153_Y));
KC_OAI21_X1 T2950 ( .B(T2949_Q), .A0(T3509_Y), .A1(T10570_Y),     .Y(T2950_Y));
KC_OAI21_X1 T3186 ( .B(T5747_Y), .A0(T14516_Q), .A1(T5748_Y),     .Y(T3186_Y));
KC_OAI21_X1 T3220 ( .B(T15694_Y), .A0(T3816_Y), .A1(T5101_Y),     .Y(T3220_Y));
KC_OAI21_X1 T3278 ( .B(T8206_Y), .A0(T3282_Y), .A1(T4384_Y),     .Y(T3278_Y));
KC_OAI21_X1 T16044 ( .B(T3374_Y), .A0(T15760_Q), .A1(T16031_Y),     .Y(T16044_Y));
KC_OAI21_X1 T16034 ( .B(T11996_Y), .A0(T6044_Y), .A1(T6034_Y),     .Y(T16034_Y));
KC_OAI21_X1 T3405 ( .B(T6045_Y), .A0(T11663_Y), .A1(T5116_Y),     .Y(T3405_Y));
KC_OAI21_X1 T3406 ( .B(T15622_Y), .A0(T16105_Y), .A1(T10965_Y),     .Y(T3406_Y));
KC_OAI21_X1 T3410 ( .B(T6045_Y), .A0(T11661_Y), .A1(T11647_Y),     .Y(T3410_Y));
KC_OAI21_X1 T3452 ( .B(T6139_Y), .A0(T11725_Y), .A1(T10975_Y),     .Y(T3452_Y));
KC_OAI21_X1 T3453 ( .B(T6067_Y), .A0(T15623_Y), .A1(T8342_Y),     .Y(T3453_Y));
KC_OAI21_X1 T3456 ( .B(T11831_Y), .A0(T11739_Y), .A1(T10620_Y),     .Y(T3456_Y));
KC_OAI21_X1 T3457 ( .B(T10587_Y), .A0(T4081_Y), .A1(T4079_Y),     .Y(T3457_Y));
KC_OAI21_X1 T3459 ( .B(T11746_Y), .A0(T6112_Y), .A1(T10588_Y),     .Y(T3459_Y));
KC_OAI21_X1 T3460 ( .B(T8510_Y), .A0(T3404_Y), .A1(T11719_Y),     .Y(T3460_Y));
KC_OAI21_X1 T3461 ( .B(T10975_Y), .A0(T3412_Q), .A1(T6120_Y),     .Y(T3461_Y));
KC_OAI21_X1 T3494 ( .B(T6561_Y), .A0(T12056_Y), .A1(T13191_Y),     .Y(T3494_Y));
KC_OAI21_X1 T3495 ( .B(T3447_Y), .A0(T8361_Y), .A1(T6824_Y),     .Y(T3495_Y));
KC_OAI21_X1 T3499 ( .B(T4122_Y), .A0(T2356_Y), .A1(T3489_Y),     .Y(T3499_Y));
KC_OAI21_X1 T3500 ( .B(T10984_Y), .A0(T6209_Y), .A1(T12870_Y),     .Y(T3500_Y));
KC_OAI21_X1 T16246 ( .B(T3735_Y), .A0(T16251_Y), .A1(T10096_Y),     .Y(T16246_Y));
KC_OAI21_X1 T3773 ( .B(T3735_Y), .A0(T16250_Y), .A1(T10096_Y),     .Y(T3773_Y));
KC_OAI21_X1 T3819 ( .B(T5763_Y), .A0(T15868_Y), .A1(T11389_Y),     .Y(T3819_Y));
KC_OAI21_X1 T3820 ( .B(T4465_Q), .A0(T5801_Y), .A1(T3797_Y),     .Y(T3820_Y));
KC_OAI21_X1 T3821 ( .B(T3802_Y), .A0(T16241_Y), .A1(T4486_Y),     .Y(T3821_Y));
KC_OAI21_X1 T3852 ( .B(T15896_Y), .A0(T3830_Y), .A1(T5790_Y),     .Y(T3852_Y));
KC_OAI21_X1 T3853 ( .B(T3826_Y), .A0(T15908_Y), .A1(T5789_Y),     .Y(T3853_Y));
KC_OAI21_X1 T3855 ( .B(T5826_Y), .A0(T11353_Y), .A1(T5789_Y),     .Y(T3855_Y));
KC_OAI21_X1 T3882 ( .B(T11519_Y), .A0(T2700_Y), .A1(T2699_Y),     .Y(T3882_Y));
KC_OAI21_X1 T3899 ( .B(T3896_Y), .A0(T4505_Y), .A1(T12804_Y),     .Y(T3899_Y));
KC_OAI21_X1 T3927 ( .B(T5905_Y), .A0(T5907_Y), .A1(T3932_Y),     .Y(T3927_Y));
KC_OAI21_X1 T3928 ( .B(T3911_Y), .A0(T3906_Y), .A1(T3914_Y),     .Y(T3928_Y));
KC_OAI21_X1 T3953 ( .B(T3980_Y), .A0(T3941_Y), .A1(T11577_Y),     .Y(T3953_Y));
KC_OAI21_X1 T3966 ( .B(T6265_Y), .A0(T5914_Y), .A1(T4549_Y),     .Y(T3966_Y));
KC_OAI21_X1 T3967 ( .B(T10937_Y), .A0(T15586_Y), .A1(T15968_Y),     .Y(T3967_Y));
KC_OAI21_X1 T4007 ( .B(T15622_Y), .A0(T2723_Y), .A1(T2849_Y),     .Y(T4007_Y));
KC_OAI21_X1 T4038 ( .B(T8505_Y), .A0(T6155_Y), .A1(T4015_Y),     .Y(T4038_Y));
KC_OAI21_X1 T4098 ( .B(T6806_Y), .A0(T5056_Y), .A1(T10972_Y),     .Y(T4098_Y));
KC_OAI21_X1 T4100 ( .B(T6098_Y), .A0(T8373_Y), .A1(T4049_Y),     .Y(T4100_Y));
KC_OAI21_X1 T6562 ( .B(T4119_Y), .A0(T6207_Y), .A1(T6587_Y),     .Y(T6562_Y));
KC_OAI21_X1 T4150 ( .B(T4140_Y), .A0(T2865_Y), .A1(T6558_Y),     .Y(T4150_Y));
KC_OAI21_X1 T4170 ( .B(T4152_Y), .A0(T2865_Y), .A1(T12860_Y),     .Y(T4170_Y));
KC_OAI21_X1 T4189 ( .B(T5721_Y), .A0(T5712_Y), .A1(T6645_Y),     .Y(T4189_Y));
KC_OAI21_X1 T6447 ( .B(T3025_Y), .A0(T4202_Y), .A1(T10432_Y),     .Y(T6447_Y));
KC_OAI21_X1 T4210 ( .B(T3025_Y), .A0(T4205_Y), .A1(T10433_Y),     .Y(T4210_Y));
KC_OAI21_X1 T4211 ( .B(T3585_Y), .A0(T4204_Y), .A1(T4202_Y),     .Y(T4211_Y));
KC_OAI21_X1 T4212 ( .B(T3585_Y), .A0(T4203_Y), .A1(T4202_Y),     .Y(T4212_Y));
KC_OAI21_X1 T4213 ( .B(T3025_Y), .A0(T4204_Y), .A1(T4205_Y),     .Y(T4213_Y));
KC_OAI21_X1 T4214 ( .B(T3025_Y), .A0(T4203_Y), .A1(T4205_Y),     .Y(T4214_Y));
KC_OAI21_X1 T4215 ( .B(T3025_Y), .A0(T4202_Y), .A1(T10433_Y),     .Y(T4215_Y));
KC_OAI21_X1 T4216 ( .B(T3025_Y), .A0(T4205_Y), .A1(T10432_Y),     .Y(T4216_Y));
KC_OAI21_X1 T4286 ( .B(T4283_Y), .A0(T4267_Y), .A1(T4265_Y),     .Y(T4286_Y));
KC_OAI21_X1 T4274 ( .B(T4283_Y), .A0(T4266_Y), .A1(T4268_Y),     .Y(T4274_Y));
KC_OAI21_X1 T4276 ( .B(T4283_Y), .A0(T4266_Y), .A1(T4265_Y),     .Y(T4276_Y));
KC_OAI21_X1 T4277 ( .B(T15782_Y), .A0(T5173_Y), .A1(T16444_Y),     .Y(T4277_Y));
KC_OAI21_X1 T4278 ( .B(T4283_Y), .A0(T4268_Y), .A1(T9859_Y),     .Y(T4278_Y));
KC_OAI21_X1 T4279 ( .B(T4283_Y), .A0(T4265_Y), .A1(T9859_Y),     .Y(T4279_Y));
KC_OAI21_X1 T4280 ( .B(T4283_Y), .A0(T4268_Y), .A1(T9860_Y),     .Y(T4280_Y));
KC_OAI21_X1 T4281 ( .B(T4283_Y), .A0(T4267_Y), .A1(T4268_Y),     .Y(T4281_Y));
KC_OAI21_X1 T4285 ( .B(T4283_Y), .A0(T4265_Y), .A1(T9860_Y),     .Y(T4285_Y));
KC_OAI21_X1 T16292 ( .B(T3735_Y), .A0(T4318_Y), .A1(T16251_Y),     .Y(T16292_Y));
KC_OAI21_X1 T4326 ( .B(T3735_Y), .A0(T4318_Y), .A1(T16250_Y),     .Y(T4326_Y));
KC_OAI21_X1 T16247 ( .B(T3735_Y), .A0(T16248_Y), .A1(T16250_Y),     .Y(T16247_Y));
KC_OAI21_X1 T4405 ( .B(T5781_Y), .A0(T11976_Y), .A1(T5815_Y),     .Y(T4405_Y));
KC_OAI21_X1 T4420 ( .B(T11428_Y), .A0(T11322_Y), .A1(T13071_Y),     .Y(T4420_Y));
KC_OAI21_X1 T4421 ( .B(T10888_Y), .A0(T15557_Y), .A1(T4485_Y),     .Y(T4421_Y));
KC_OAI21_X1 T15876 ( .B(T4445_Y), .A0(T16153_Y), .A1(T8184_Y),     .Y(T15876_Y));
KC_OAI21_X1 T4458 ( .B(T11977_Y), .A0(T14551_Q), .A1(T11393_Y),     .Y(T4458_Y));
KC_OAI21_X1 T4460 ( .B(T3856_Y), .A0(T11421_Y), .A1(T11973_Y),     .Y(T4460_Y));
KC_OAI21_X1 T4461 ( .B(T15872_Y), .A0(T5815_Y), .A1(T4500_Y),     .Y(T4461_Y));
KC_OAI21_X1 T4464 ( .B(T4463_Y), .A0(T16153_Y), .A1(T4478_Y),     .Y(T4464_Y));
KC_OAI21_X1 T4504 ( .B(T5107_Y), .A0(T8444_Y), .A1(T6128_Y),     .Y(T4504_Y));
KC_OAI21_X1 T4536 ( .B(T10931_Y), .A0(T16302_Y), .A1(T4557_Y),     .Y(T4536_Y));
KC_OAI21_X1 T4566 ( .B(T15970_Y), .A0(T12352_Y), .A1(T3940_Y),     .Y(T4566_Y));
KC_OAI21_X1 T4567 ( .B(T4560_Y), .A0(T3945_Y), .A1(T4551_Y),     .Y(T4567_Y));
KC_OAI21_X1 T4569 ( .B(T4474_Y), .A0(T5969_Y), .A1(T4550_Y),     .Y(T4569_Y));
KC_OAI21_X1 T16062 ( .B(T16061_Y), .A0(T4644_Y), .A1(T4667_Y),     .Y(T16062_Y));
KC_OAI21_X1 T16061 ( .B(T4675_Q), .A0(T4667_Y), .A1(T12032_Y),     .Y(T16061_Y));
KC_OAI21_X1 T16060 ( .B(T5501_Q), .A0(T4645_Y), .A1(T12032_Y),     .Y(T16060_Y));
KC_OAI21_X1 T16059 ( .B(T4674_Y), .A0(T4642_Y), .A1(T4639_Y),     .Y(T16059_Y));
KC_OAI21_X1 T16048 ( .B(T4056_Q), .A0(T4666_Y), .A1(T12032_Y),     .Y(T16048_Y));
KC_OAI21_X1 T16046 ( .B(T4685_Q), .A0(T4654_Y), .A1(T12032_Y),     .Y(T16046_Y));
KC_OAI21_X1 T4666 ( .B(T4726_Y), .A0(T11706_Y), .A1(T16110_Y),     .Y(T4666_Y));
KC_OAI21_X1 T4667 ( .B(T12855_Y), .A0(T11706_Y), .A1(T16110_Y),     .Y(T4667_Y));
KC_OAI21_X1 T4670 ( .B(T4672_Y), .A0(T4655_Y), .A1(T4640_Y),     .Y(T4670_Y));
KC_OAI21_X1 T4671 ( .B(T16049_Q), .A0(T4658_Y), .A1(T12032_Y),     .Y(T4671_Y));
KC_OAI21_X1 T4672 ( .B(T4686_Q), .A0(T4640_Y), .A1(T12032_Y),     .Y(T4672_Y));
KC_OAI21_X1 T4673 ( .B(T16060_Y), .A0(T4647_Y), .A1(T4645_Y),     .Y(T4673_Y));
KC_OAI21_X1 T4674 ( .B(T4714_Q), .A0(T4639_Y), .A1(T11705_Y),     .Y(T4674_Y));
KC_OAI21_X1 T4676 ( .B(T5502_Q), .A0(T12032_Y), .A1(T16047_Y),     .Y(T4676_Y));
KC_OAI21_X1 T4677 ( .B(T16046_Y), .A0(T4656_Y), .A1(T4654_Y),     .Y(T4677_Y));
KC_OAI21_X1 T4678 ( .B(T4693_Q), .A0(T12032_Y), .A1(T4657_Y),     .Y(T4678_Y));
KC_OAI21_X1 T4679 ( .B(T4682_Y), .A0(T4660_Y), .A1(T4643_Y),     .Y(T4679_Y));
KC_OAI21_X1 T4680 ( .B(T16048_Y), .A0(T4659_Y), .A1(T4666_Y),     .Y(T4680_Y));
KC_OAI21_X1 T4681 ( .B(T5496_Q), .A0(T11705_Y), .A1(T4646_Y),     .Y(T4681_Y));
KC_OAI21_X1 T4682 ( .B(T4043_Q), .A0(T4643_Y), .A1(T11705_Y),     .Y(T4682_Y));
KC_OAI21_X1 T4683 ( .B(T4671_Y), .A0(T4653_Y), .A1(T4658_Y),     .Y(T4683_Y));
KC_OAI21_X1 T4684 ( .B(T4663_Q), .A0(T11705_Y), .A1(T4652_Y),     .Y(T4684_Y));
KC_OAI21_X1 T4725 ( .B(T6467_Y), .A0(T4719_Q), .A1(T10989_Y),     .Y(T4725_Y));
KC_OAI21_X1 T4726 ( .B(T6448_Y), .A0(T4719_Q), .A1(T10981_Y),     .Y(T4726_Y));
KC_OAI21_X1 T4727 ( .B(T5153_Y), .A0(T4648_Y), .A1(T4637_Y),     .Y(T4727_Y));
KC_OAI21_X1 T6548 ( .B(T4742_Y), .A0(T12302_Y), .A1(T286_Y),     .Y(T6548_Y));
KC_OAI21_X1 T4753 ( .B(T4738_Y), .A0(T11777_Y), .A1(T15625_Y),     .Y(T4753_Y));
KC_OAI21_X1 T9474 ( .B(T216_Y), .A0(T605_Q), .A1(T15538_Y),     .Y(T9474_Y));
KC_OAI21_X1 T4824 ( .B(T16335_Y), .A0(T7826_Y), .A1(T16333_Y),     .Y(T4824_Y));
KC_OAI21_X1 T4834 ( .B(T7249_Y), .A0(T4835_Q), .A1(T6346_Y),     .Y(T4834_Y));
KC_OAI21_X1 T4857 ( .B(T585_Y), .A0(T11171_Y), .A1(T6822_Y),     .Y(T4857_Y));
KC_OAI21_X1 T4859 ( .B(T8029_Y), .A0(T1094_Q), .A1(T7976_Y),     .Y(T4859_Y));
KC_OAI21_X1 T4863 ( .B(T585_Y), .A0(T11193_Y), .A1(T6822_Y),     .Y(T4863_Y));
KC_OAI21_X1 T4892 ( .B(T1492_Y), .A0(T7705_Y), .A1(T9810_Y),     .Y(T4892_Y));
KC_OAI21_X1 T4972 ( .B(T2604_Y), .A0(T16371_Y), .A1(T5369_Y),     .Y(T4972_Y));
KC_OAI21_X1 T5060 ( .B(T3467_Y), .A0(T11598_Y), .A1(T6515_Y),     .Y(T5060_Y));
KC_OAI21_X1 T16257 ( .B(T3735_Y), .A0(T16250_Y), .A1(T10095_Y),     .Y(T16257_Y));
KC_OAI21_X1 T5120 ( .B(T12205_Y), .A0(T11555_Y), .A1(T11024_Y),     .Y(T5120_Y));
KC_OAI21_X1 T5125 ( .B(T15997_Y), .A0(T16453_Q), .A1(T16454_Q),     .Y(T5125_Y));
KC_OAI21_X1 T5126 ( .B(T15622_Y), .A0(T6011_Y), .A1(T2849_Y),     .Y(T5126_Y));
KC_OAI21_X1 T5151 ( .B(T4706_Y), .A0(T15756_Y), .A1(T4735_Y),     .Y(T5151_Y));
KC_OAI21_X1 T5153 ( .B(T5513_Q), .A0(T4637_Y), .A1(T11705_Y),     .Y(T5153_Y));
KC_OAI21_X1 T5155 ( .B(T3258_Q), .A0(T4521_Y), .A1(T15964_Y),     .Y(T5155_Y));
KC_OAI21_X1 T5183 ( .B(T1419_Y), .A0(T10380_Y), .A1(T9541_Y),     .Y(T5183_Y));
KC_OAI21_X1 T5217 ( .B(T1419_Y), .A0(T6992_Y), .A1(T6990_Y),     .Y(T5217_Y));
KC_OAI21_X1 T5218 ( .B(T1419_Y), .A0(T6992_Y), .A1(T10380_Y),     .Y(T5218_Y));
KC_OAI21_X1 T5219 ( .B(T1419_Y), .A0(T10380_Y), .A1(T9540_Y),     .Y(T5219_Y));
KC_OAI21_X1 T6837 ( .B(T4885_Y), .A0(T7541_Y), .A1(T7542_Y),     .Y(T6837_Y));
KC_OAI21_X1 T5273 ( .B(T1453_Y), .A0(T7489_Y), .A1(T7490_Y),     .Y(T5273_Y));
KC_OAI21_X1 T5296 ( .B(T8939_Y), .A0(T5348_Q), .A1(T725_Q),     .Y(T5296_Y));
KC_OAI21_X1 T5312 ( .B(T12330_Y), .A0(T1107_Y), .A1(T16406_Y),     .Y(T5312_Y));
KC_OAI21_X1 T5352 ( .B(T7883_Y), .A0(T8854_Y), .A1(T7892_Y),     .Y(T5352_Y));
KC_OAI21_X1 T5370 ( .B(T10023_Y), .A0(T1128_Q), .A1(T5340_Q),     .Y(T5370_Y));
KC_OAI21_X1 T5372 ( .B(T10023_Y), .A0(T1135_Q), .A1(T1220_Q),     .Y(T5372_Y));
KC_OAI21_X1 T5395 ( .B(T2057_Y), .A0(T15503_Y), .A1(T15501_Y),     .Y(T5395_Y));
KC_OAI21_X1 T5410 ( .B(T3735_Y), .A0(T16248_Y), .A1(T16251_Y),     .Y(T5410_Y));
KC_OAI21_X1 T5430 ( .B(T6059_Y), .A0(T3795_Y), .A1(T5783_Y),     .Y(T5430_Y));
KC_OAI21_X1 T5431 ( .B(T3797_Y), .A0(T11969_Y), .A1(T3794_Y),     .Y(T5431_Y));
KC_OAI21_X1 T5435 ( .B(T15865_Y), .A0(T11370_Y), .A1(T11983_Y),     .Y(T5435_Y));
KC_OAI21_X1 T5440 ( .B(T5826_Y), .A0(T8202_Y), .A1(T13089_Y),     .Y(T5440_Y));
KC_OAI21_X1 T5471 ( .B(T10959_Y), .A0(T2809_Q), .A1(T2217_Y),     .Y(T5471_Y));
KC_OAI21_X1 T5487 ( .B(T2235_Y), .A0(T2854_Y), .A1(T12220_Y),     .Y(T5487_Y));
KC_OAI21_X1 T5500 ( .B(T10967_Y), .A0(T8468_Y), .A1(T10971_Y),     .Y(T5500_Y));
KC_OAI21_X1 T16125 ( .B(T6806_Y), .A0(T15623_Y), .A1(T10972_Y),     .Y(T16125_Y));
KC_OAI21_X1 T5509 ( .B(T12284_Y), .A0(T10625_Y), .A1(T2871_Y),     .Y(T5509_Y));
KC_OAI21_X1 T16252 ( .B(T3735_Y), .A0(T16251_Y), .A1(T10095_Y),     .Y(T16252_Y));
KC_MXI2B_X2 T16418 ( .Y(T16418_Y), .A(T8082_Y), .BN(T8916_Y),     .S0(T7908_Y));
KC_MXI2B_X2 T16327 ( .Y(T16327_Y), .A(T9387_Y), .BN(T9379_Y),     .S0(T7575_Y));
KC_MXI2B_X2 T3277 ( .Y(T3277_Y), .A(T526_Q), .BN(T183_Q), .S0(T166_Q));
KC_MXI2B_X2 T16430 ( .Y(T16430_Y), .A(T15059_Y), .BN(T8692_Y),     .S0(T745_Y));
KC_MXI2B_X2 T8835 ( .Y(T8835_Y), .A(T15062_Y), .BN(T8694_Y),     .S0(T745_Y));
KC_MXI2B_X2 T16428 ( .Y(T16428_Y), .A(T15065_Y), .BN(T8691_Y),     .S0(T745_Y));
KC_MXI2B_X2 T8809 ( .Y(T8809_Y), .A(T15143_Y), .BN(T8689_Y),     .S0(T745_Y));
KC_MXI2B_X2 T16419 ( .Y(T16419_Y), .A(T15074_Y), .BN(T8690_Y),     .S0(T745_Y));
KC_MXI2B_X2 T5143 ( .Y(T5143_Y), .A(T15066_Y), .BN(T8738_Y),     .S0(T745_Y));
KC_MXI2B_X2 T5108 ( .Y(T5108_Y), .A(T15063_Y), .BN(T8695_Y),     .S0(T745_Y));
KC_MXI2B_X2 T6834 ( .Y(T6834_Y), .A(T5280_Q), .BN(T689_Q),     .S0(T697_Q));
KC_MXI2B_X2 T16423 ( .Y(T16423_Y), .A(T1100_Q), .BN(T10022_Y),     .S0(T8936_Y));
KC_MXI2B_X2 T5030 ( .Y(T5030_Y), .A(T16422_Q), .BN(T10001_Y),     .S0(T950_Y));
KC_MXI2B_X2 T4354 ( .Y(T4354_Y), .A(T13301_Y), .BN(T5793_Y),     .S0(T11971_Y));
KC_MXI2B_X2 T6570 ( .Y(T6570_Y), .A(T2358_Y), .BN(T2317_Y),     .S0(T12869_Y));
KC_MXI2B_X2 T10077 ( .Y(T10077_Y), .A(T2609_Y), .BN(T2628_Q),     .S0(T12735_Y));
KC_MXI2B_X2 T10194 ( .Y(T10194_Y), .A(T10936_Y), .BN(T14534_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T2861 ( .Y(T2861_Y), .A(T10880_Y), .BN(T14498_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T3783 ( .Y(T3783_Y), .A(T13131_Y), .BN(T14500_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T16195 ( .Y(T16195_Y), .A(T10941_Y), .BN(T14499_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T3782 ( .Y(T3782_Y), .A(T6118_Y), .BN(T16081_Q),     .S0(T6436_Y));
KC_MXI2B_X2 T3781 ( .Y(T3781_Y), .A(T10934_Y), .BN(T14956_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T3780 ( .Y(T3780_Y), .A(T13121_Y), .BN(T14529_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T3779 ( .Y(T3779_Y), .A(T10936_Y), .BN(T14517_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T1708 ( .Y(T1708_Y), .A(T16012_Y), .BN(T3348_Y),     .S0(T4172_Y));
KC_MXI2B_X2 T10238 ( .Y(T10238_Y), .A(T5736_Y), .BN(T14460_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T3778 ( .Y(T3778_Y), .A(T15688_Y), .BN(T14488_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T3777 ( .Y(T3777_Y), .A(T15548_Y), .BN(T14486_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T3776 ( .Y(T3776_Y), .A(T15688_Y), .BN(T14901_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T3775 ( .Y(T3775_Y), .A(T10934_Y), .BN(T14952_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T3774 ( .Y(T3774_Y), .A(T13121_Y), .BN(T14518_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T16229 ( .Y(T16229_Y), .A(T15550_Y), .BN(T14489_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16228 ( .Y(T16228_Y), .A(T5734_Y), .BN(T14468_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16227 ( .Y(T16227_Y), .A(T5563_Y), .BN(T14461_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16226 ( .Y(T16226_Y), .A(T5704_Y), .BN(T14513_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16225 ( .Y(T16225_Y), .A(T5405_Y), .BN(T14511_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16224 ( .Y(T16224_Y), .A(T5704_Y), .BN(T14512_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16223 ( .Y(T16223_Y), .A(T5706_Y), .BN(T14509_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16222 ( .Y(T16222_Y), .A(T5544_Y), .BN(T14946_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16221 ( .Y(T16221_Y), .A(T5706_Y), .BN(T14945_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16220 ( .Y(T16220_Y), .A(T15548_Y), .BN(T14472_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16219 ( .Y(T16219_Y), .A(T15549_Y), .BN(T14471_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16218 ( .Y(T16218_Y), .A(T15549_Y), .BN(T14485_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16217 ( .Y(T16217_Y), .A(T15550_Y), .BN(T14473_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16216 ( .Y(T16216_Y), .A(T5734_Y), .BN(T14487_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16215 ( .Y(T16215_Y), .A(T5729_Y), .BN(T14470_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16214 ( .Y(T16214_Y), .A(T5736_Y), .BN(T14463_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16213 ( .Y(T16213_Y), .A(T5738_Y), .BN(T14466_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16212 ( .Y(T16212_Y), .A(T5729_Y), .BN(T14469_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16211 ( .Y(T16211_Y), .A(T5790_Y), .BN(T3830_Y),     .S0(T6068_Y));
KC_MXI2B_X2 T15962 ( .Y(T15962_Y), .A(T6173_Y), .BN(T12195_Y),     .S0(T12194_Y));
KC_MXI2B_X2 T16210 ( .Y(T16210_Y), .A(T12278_Y), .BN(T4048_Q),     .S0(T12286_Y));
KC_MXI2B_X2 T16209 ( .Y(T16209_Y), .A(T5741_Y), .BN(T14894_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16208 ( .Y(T16208_Y), .A(T5740_Y), .BN(T14483_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16207 ( .Y(T16207_Y), .A(T5740_Y), .BN(T14467_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16206 ( .Y(T16206_Y), .A(T5563_Y), .BN(T14459_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16205 ( .Y(T16205_Y), .A(T5405_Y), .BN(T14508_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T16204 ( .Y(T16204_Y), .A(T5741_Y), .BN(T14484_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T16203 ( .Y(T16203_Y), .A(T5738_Y), .BN(T14482_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T4410 ( .Y(T4410_Y), .A(T12803_Y), .BN(T3896_Y),     .S0(T3899_Y));
KC_MXI2B_X2 T8247 ( .Y(T8247_Y), .A(T15971_Y), .BN(T5885_Y),     .S0(T5888_Y));
KC_MXI2B_X2 T16473 ( .Y(T16473_Y), .A(T2389_Y), .BN(T14969_Y),     .S0(T6356_Y));
KC_MXI2B_X2 T16193 ( .Y(T16193_Y), .A(T13125_Y), .BN(T14530_Q),     .S0(T2640_Q));
KC_MXI2B_X2 T16114 ( .Y(T16114_Y), .A(T15546_Y), .BN(T14943_Q),     .S0(T15825_Y));
KC_MXI2B_X2 T5148 ( .Y(T5148_Y), .A(T5544_Y), .BN(T14507_Q),     .S0(T15835_Y));
KC_MXI2B_X2 T5548 ( .Y(T5548_Y), .A(T13125_Y), .BN(T14521_Q),     .S0(T2640_Q));
KC_AOI22B_X2 T16133 ( .B1(T10560_Y), .B0(T15712_Y), .A1(T12102_Y),     .Y(T16133_Y), .A0N(T10559_Y));
KC_AO22_X1 T15779 ( .B0(T10651_Y), .B1(T1070_Q), .A1(T1075_Y),     .A0(T1071_Q), .Y(T15779_Y));
KC_AO22_X1 T15777 ( .B0(T10651_Y), .B1(T1072_Q), .A1(T1063_Y),     .A0(T1073_Q), .Y(T15777_Y));
KC_AO22_X1 T15776 ( .B0(T10651_Y), .B1(T1069_Q), .A1(T1075_Y),     .A0(T1061_Q), .Y(T15776_Y));
KC_AO22_X1 T15775 ( .B0(T10651_Y), .B1(T1067_Q), .A1(T1063_Y),     .A0(T1064_Q), .Y(T15775_Y));
KC_AO22_X1 T15773 ( .B0(T10651_Y), .B1(T1076_Q), .A1(T4859_Y),     .A0(T1078_Q), .Y(T15773_Y));
KC_AO22_X1 T15792 ( .B0(T10651_Y), .B1(T1091_Q), .A1(T1087_Y),     .A0(T8834_Q), .Y(T15792_Y));
KC_AO22_X1 T15781 ( .B0(T1065_Q), .B1(T15466_Y), .A1(T15664_Y),     .A0(T1183_Q), .Y(T15781_Y));
KC_AO22_X1 T15778 ( .B0(T5293_Q), .B1(T15466_Y), .A1(T15664_Y),     .A0(T1186_Q), .Y(T15778_Y));
KC_AO22_X1 T15774 ( .B0(T5292_Q), .B1(T15466_Y), .A1(T15664_Y),     .A0(T1185_Q), .Y(T15774_Y));
KC_AO22_X1 T15810 ( .B0(T2073_Y), .B1(T15085_Y), .A1(T10160_Y),     .A0(T8975_Y), .Y(T15810_Y));
KC_AO22_X1 T15893 ( .B0(T16156_Y), .B1(T12100_Y), .A1(T2104_Y),     .A0(T2112_Q), .Y(T15893_Y));
KC_AO22_X1 T15885 ( .B0(T16156_Y), .B1(T12099_Y), .A1(T4943_Y),     .A0(T2118_Q), .Y(T15885_Y));
KC_AO22_X1 T15884 ( .B0(T16156_Y), .B1(T15812_Y), .A1(T2145_Y),     .A0(T2119_Q), .Y(T15884_Y));
KC_AO22_X1 T15913 ( .B0(T16156_Y), .B1(T16471_Q), .A1(T2132_Y),     .A0(T6071_Q), .Y(T15913_Y));
KC_AO22_X1 T15958 ( .B0(T16156_Y), .B1(T10739_Y), .A1(T13117_Y),     .A0(T5463_Q), .Y(T15958_Y));
KC_AO22_X1 T15975 ( .B0(T11586_Y), .B1(T2113_Q), .A1(T16072_Y),     .A0(T15232_Y), .Y(T15975_Y));
KC_AO22_X1 T6505 ( .B0(T2386_Y), .B1(T2956_Y), .A1(T8432_Y),     .A0(T2951_Y), .Y(T6505_Y));
KC_AO22_X1 T16098 ( .B0(T10203_Y), .B1(T2515_Y), .A1(T3166_Y),     .A0(T16236_Y), .Y(T16098_Y));
KC_AO22_X1 T16097 ( .B0(T10203_Y), .B1(T2469_Y), .A1(T3713_Y),     .A0(T16236_Y), .Y(T16097_Y));
KC_AO22_X1 T16096 ( .B0(T10203_Y), .B1(T2485_Y), .A1(T4291_Y),     .A0(T16236_Y), .Y(T16096_Y));
KC_AO22_X1 T16076 ( .B0(T10203_Y), .B1(T2516_Y), .A1(T3177_Y),     .A0(T16236_Y), .Y(T16076_Y));
KC_AO22_X1 T16075 ( .B0(T10203_Y), .B1(T2470_Y), .A1(T3692_Y),     .A0(T16236_Y), .Y(T16075_Y));
KC_AO22_X1 T16074 ( .B0(T10203_Y), .B1(T2483_Y), .A1(T3685_Y),     .A0(T16236_Y), .Y(T16074_Y));
KC_AO22_X1 T16073 ( .B0(T10203_Y), .B1(T2461_Y), .A1(T5322_Y),     .A0(T16236_Y), .Y(T16073_Y));
KC_AO22_X1 T16072 ( .B0(T10203_Y), .B1(T2468_Y), .A1(T4307_Y),     .A0(T16236_Y), .Y(T16072_Y));
KC_AO22_X1 T16071 ( .B0(T10203_Y), .B1(T2514_Y), .A1(T3742_Y),     .A0(T16236_Y), .Y(T16071_Y));
KC_AO22_X1 T16069 ( .B0(T10203_Y), .B1(T4987_Y), .A1(T3739_Y),     .A0(T16236_Y), .Y(T16069_Y));
KC_AO22_X1 T16053 ( .B0(T6066_Y), .B1(T2844_Q), .A1(T8362_Y),     .A0(T11666_Y), .Y(T16053_Y));
KC_AO22_X1 T15944 ( .B0(T5942_Y), .B1(T3309_Y), .A1(T3285_Y),     .A0(T8266_Y), .Y(T15944_Y));
KC_AO22_X1 T15998 ( .B0(T12960_Y), .B1(T6772_Y), .A1(T15992_Y),     .A0(T12216_Y), .Y(T15998_Y));
KC_AO22_X1 T15931 ( .B0(T3890_Q), .B1(T10634_Y), .A1(T10635_Y),     .A0(T3873_Q), .Y(T15931_Y));
KC_AO22_X1 T16027 ( .B0(T5992_Y), .B1(T4042_Y), .A1(T16029_Y),     .A0(T5992_Y), .Y(T16027_Y));
KC_AO22_X1 T6525 ( .B0(T4153_Y), .B1(T4175_Y), .A1(T4761_Y),     .A0(T3996_Y), .Y(T6525_Y));
KC_AO22_X1 T15909 ( .B0(T4479_Y), .B1(T3222_Y), .A1(T4503_Y),     .A0(T5857_Y), .Y(T15909_Y));
KC_AO22_X1 T15946 ( .B0(T4524_Y), .B1(T4524_Y), .A1(T5156_Y),     .A0(T4524_Y), .Y(T15946_Y));
KC_AO22_X1 T16087 ( .B0(T15492_Y), .B1(T9080_S), .A1(T9451_Y),     .A0(T15077_Y), .Y(T16087_Y));
KC_AO22_X1 T16086 ( .B0(T972_Y), .B1(T9443_Y), .A1(T10069_Y),     .A0(T601_Y), .Y(T16086_Y));
KC_AO22_X1 T16092 ( .B0(T10651_Y), .B1(T4860_Q), .A1(T1087_Y),     .A0(T1122_Q), .Y(T16092_Y));
KC_AO22_X1 T16091 ( .B0(T10651_Y), .B1(T1088_Q), .A1(T4859_Y),     .A0(T1121_Q), .Y(T16091_Y));
KC_AO22_X1 T15972 ( .B0(T16156_Y), .B1(T10659_Y), .A1(T13314_Y),     .A0(T5473_Q), .Y(T15972_Y));
KC_AO22_X1 T6546 ( .B0(T12069_Y), .B1(T6545_Y), .A1(T11038_Y),     .A0(T11038_Y), .Y(T6546_Y));
KC_AO22_X1 T15780 ( .B0(T5294_Q), .B1(T15466_Y), .A1(T15664_Y),     .A0(T1184_Q), .Y(T15780_Y));
KC_AO22_X1 T15772 ( .B0(T1077_Q), .B1(T15466_Y), .A1(T15664_Y),     .A0(T1187_Q), .Y(T15772_Y));
KC_AO22_X1 T15813 ( .B0(T15518_Y), .B1(T2360_Q), .A1(T2622_Y),     .A0(T5388_Q), .Y(T15813_Y));
KC_AO22_X1 T16070 ( .B0(T10203_Y), .B1(T2511_Y), .A1(T3161_Y),     .A0(T16236_Y), .Y(T16070_Y));
KC_AO22_X1 T16012 ( .B0(T3327_Y), .B1(T12961_Y), .A1(T6776_S),     .A0(T3327_Y), .Y(T16012_Y));
KC_AO22_X1 T16090 ( .B0(T5333_Q), .B1(T15466_Y), .A1(T15664_Y),     .A0(T1189_Q), .Y(T16090_Y));
KC_AO21_X2 T16429 ( .A0(T8868_Y), .B(T13246_Y), .Y(T16429_Y),     .A1(T7912_Y));
KC_AO21_X2 T10264 ( .A0(T8741_Y), .B(T13238_Y), .Y(T10264_Y),     .A1(T7814_Y));
KC_AO21_X2 T15999 ( .A0(T3294_Y), .B(T4052_Q), .Y(T15999_Y),     .A1(T6769_Y));
KC_DFFRNHQ_X3 T6359 ( .RN(T7073_Y), .Q(T6359_Q), .D(T15336_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T6358 ( .RN(T14975_Y), .Q(T6358_Q), .D(T736_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T6357 ( .RN(T14975_Y), .Q(T6357_Q), .D(T11209_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T6355 ( .RN(T7073_Y), .Q(T6355_Q), .D(T53_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T2319 ( .RN(T7609_Y), .Q(T2319_Q), .D(T8723_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6379 ( .RN(T7609_Y), .Q(T6379_Q), .D(T7812_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6371 ( .RN(T7609_Y), .Q(T6371_Q), .D(T11205_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6369 ( .RN(T7609_Y), .Q(T6369_Q), .D(T16376_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6364 ( .RN(T7609_Y), .Q(T6364_Q), .D(T15786_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6684 ( .RN(T7675_Y), .Q(T6684_Q), .D(T8808_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6412 ( .RN(T7609_Y), .Q(T6412_Q), .D(T15722_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6411 ( .RN(T7609_Y), .Q(T6411_Q), .D(T10264_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6401 ( .RN(T7609_Y), .Q(T6401_Q), .D(T11208_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6391 ( .RN(T7609_Y), .Q(T6391_Q), .D(T7385_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6425 ( .RN(T7675_Y), .Q(T6425_Q), .D(T11235_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6424 ( .RN(T7675_Y), .Q(T6424_Q), .D(T15839_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6423 ( .RN(T7675_Y), .Q(T6423_Q), .D(T7813_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6422 ( .RN(T7675_Y), .Q(T6422_Q), .D(T16162_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6416 ( .RN(T7675_Y), .Q(T6416_Q), .D(T7623_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T16085 ( .RN(T7675_Y), .Q(T16085_Q), .D(T15031_Y),     .CK(T4828_Y));
KC_DFFRNHQ_X3 T6430 ( .RN(T7675_Y), .Q(T6430_Q), .D(T15840_Y),     .CK(T4828_Y));
KC_DFFRNHQ_X3 T6432 ( .RN(T7074_Y), .Q(T6432_Q), .D(T7607_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T6361 ( .RN(T7073_Y), .Q(T6361_Q), .D(T7810_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T6417 ( .RN(T7675_Y), .Q(T6417_Q), .D(T11238_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T15795 ( .RN(T14997_Y), .Q(T15795_Q), .D(T11291_Y),     .CK(T594_Y));
KC_DFFRNHQ_X3 T16301 ( .RN(T15001_Y), .Q(T16301_Q), .D(T9004_Y),     .CK(T971_Y));
KC_DFFRNHQ_X3 T15798 ( .RN(T15001_Y), .Q(T15798_Q), .D(T1739_Y),     .CK(T971_Y));
KC_DFFRNHQ_X3 T15797 ( .RN(T15001_Y), .Q(T15797_Q), .D(T973_Y),     .CK(T971_Y));
KC_DFFRNHQ_X3 T15796 ( .RN(T15001_Y), .Q(T15796_Q), .D(T9037_Y),     .CK(T971_Y));
KC_DFFRNHQ_X3 T16088 ( .RN(T10727_Y), .Q(T16088_Q), .D(T9039_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T16299 ( .RN(T10727_Y), .Q(T16299_Q), .D(T4805_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T15844 ( .RN(T15002_Y), .Q(T15844_Q), .D(T9003_Y),     .CK(T971_Y));
KC_DFFRNHQ_X3 T15808 ( .RN(T10727_Y), .Q(T15808_Q), .D(T1732_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T15807 ( .RN(T10727_Y), .Q(T15807_Q), .D(T1634_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T15806 ( .RN(T1283_RN), .Q(T15806_Q), .D(T1283_Q),     .CK(T5725_Y));
KC_DFFRNHQ_X3 T15805 ( .RN(T10727_Y), .Q(T15805_Q), .D(T16086_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T15804 ( .RN(T10661_Y), .Q(T15804_Q), .D(T8998_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T15828 ( .RN(T15008_Y), .Q(T15828_Q), .D(T2120_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X3 T16007 ( .RN(T15018_Y), .Q(T16007_Q), .D(T8485_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X3 T15990 ( .RN(T15018_Y), .Q(T15990_Q), .D(T8283_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X3 T16018 ( .RN(T15018_Y), .Q(T16018_Q), .D(T12832_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X3 T16010 ( .RN(T15018_Y), .Q(T16010_Q), .D(T11623_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X3 T16081 ( .RN(T15021_Y), .Q(T16081_Q), .D(T3782_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X3 T6555 ( .RN(T15037_Y), .Q(T6555_Q), .D(T11783_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X3 T15894 ( .RN(T15013_Y), .Q(T15894_Q), .D(T10899_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X3 T15880 ( .RN(T15013_Y), .Q(T15880_Q), .D(T10913_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X3 T15879 ( .RN(T15008_Y), .Q(T15879_Q), .D(T10909_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X3 T5987 ( .RN(T2169_Y), .Q(T5987_Q), .D(T8287_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X3 T16023 ( .RN(T15020_Y), .Q(T16023_Q), .D(T11611_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X3 T6431 ( .RN(T2081_Y), .Q(T6431_Q), .D(T11679_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X3 T6526 ( .RN(T4047_Y), .Q(T6526_Q), .D(T4145_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X3 T15313 ( .RN(T7675_Y), .Q(T15313_Q), .D(T11234_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6730 ( .RN(T7609_Y), .Q(T6730_Q), .D(T16429_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6683 ( .RN(T7675_Y), .Q(T6683_Q), .D(T8861_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6479 ( .RN(T14975_Y), .Q(T6479_Q), .D(T8739_Y),     .CK(T175_Y));
KC_DFFRNHQ_X3 T6363 ( .RN(T7073_Y), .Q(T6363_Q), .D(T15731_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T6362 ( .RN(T7074_Y), .Q(T6362_Q), .D(T305_Y),     .CK(T138_Y));
KC_DFFRNHQ_X3 T6426 ( .RN(T7675_Y), .Q(T6426_Q), .D(T8837_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6418 ( .RN(T7675_Y), .Q(T6418_Q), .D(T11198_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T6415 ( .RN(T7675_Y), .Q(T6415_Q), .D(T16382_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X3 T15815 ( .RN(T14999_Y), .Q(T15815_Q), .D(T1714_Q),     .CK(T2050_Y));
KC_DFFRNHQ_X3 T15809 ( .RN(T10727_Y), .Q(T15809_Q), .D(T1697_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T15803 ( .RN(T10727_Y), .Q(T15803_Q), .D(T1567_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T15802 ( .RN(T10661_Y), .Q(T15802_Q), .D(T9057_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X3 T16079 ( .RN(T2063_Y), .Q(T16079_Q), .D(T5988_Y),     .CK(T14497_Q));
KC_DFFRNHQ_X3 T15860 ( .RN(T15008_Y), .Q(T15860_Q), .D(T10886_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X3 T15891 ( .RN(T15013_Y), .Q(T15891_Q), .D(T10919_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X3 T8352 ( .RN(T15021_Y), .Q(T8352_Q), .D(T2256_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X3 T15138 ( .RN(T15021_Y), .Q(T15138_Q), .D(T4947_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X3 T16082 ( .RN(T15021_Y), .Q(T16082_Q), .D(T4949_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X3 T6549 ( .RN(T4047_Y), .Q(T6549_Q), .D(T11760_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X3 T15760 ( .RN(T4047_Y), .Q(T15760_Q), .D(T12058_Y),     .CK(T14575_Q));
KC_AO12B_X2 T6446 ( .Y(T6446_Y), .B(T12083_Y), .A(T3070_Y),     .C(T1419_Y));
KC_INV_X1 T13294 ( .Y(T13294_Y), .A(T54_Q));
KC_INV_X1 T15169 ( .Y(T15169_Y), .A(T84_Q));
KC_INV_X1 T15324 ( .Y(T15324_Y), .A(T101_Q));
KC_INV_X1 T15320 ( .Y(T15320_Y), .A(T162_Q));
KC_INV_X1 T15319 ( .Y(T15319_Y), .A(T114_Q));
KC_INV_X1 T15317 ( .Y(T15317_Y), .A(T8554_Y));
KC_INV_X1 T15316 ( .Y(T15316_Y), .A(T107_Q));
KC_INV_X1 T15315 ( .Y(T15315_Y), .A(T5202_Q));
KC_INV_X1 T16479 ( .Y(T16479_Y), .A(T5203_Q));
KC_INV_X1 T15318 ( .Y(T15318_Y), .A(T8546_Y));
KC_INV_X1 T15314 ( .Y(T15314_Y), .A(T8544_Y));
KC_INV_X1 T15312 ( .Y(T15312_Y), .A(T8556_Y));
KC_INV_X1 T15336 ( .Y(T15336_Y), .A(T6856_Y));
KC_INV_X1 T6319 ( .Y(T6319_Y), .A(T136_Q));
KC_INV_X1 T6318 ( .Y(T6318_Y), .A(T5225_Q));
KC_INV_X1 T6317 ( .Y(T6317_Y), .A(T131_Q));
KC_INV_X1 T260 ( .Y(T260_Y), .A(T5192_Q));
KC_INV_X1 T257 ( .Y(T257_Y), .A(T133_Q));
KC_INV_X1 T255 ( .Y(T255_Y), .A(T9289_Y));
KC_INV_X1 T236 ( .Y(T236_Y), .A(T150_Q));
KC_INV_X1 T228 ( .Y(T228_Y), .A(T350_Y));
KC_INV_X1 T15358 ( .Y(T15358_Y), .A(T5222_Q));
KC_INV_X1 T15356 ( .Y(T15356_Y), .A(T9287_Y));
KC_INV_X1 T15353 ( .Y(T15353_Y), .A(T8602_Y));
KC_INV_X1 T878 ( .Y(T878_Y), .A(T16006_Y));
KC_INV_X1 T322 ( .Y(T322_Y), .A(T9268_Y));
KC_INV_X1 T6233 ( .Y(T6233_Y), .A(T163_Q));
KC_INV_X1 T802 ( .Y(T802_Y), .A(T4803_Q));
KC_INV_X1 T650 ( .Y(T650_Y), .A(T4802_Q));
KC_INV_X1 T648 ( .Y(T648_Y), .A(T12614_Y));
KC_INV_X1 T647 ( .Y(T647_Y), .A(T207_Q));
KC_INV_X1 T646 ( .Y(T646_Y), .A(T12608_Y));
KC_INV_X1 T645 ( .Y(T645_Y), .A(T224_Q));
KC_INV_X1 T15430 ( .Y(T15430_Y), .A(T212_Q));
KC_INV_X1 T15656 ( .Y(T15656_Y), .A(T7677_Y));
KC_INV_X1 T16289 ( .Y(T16289_Y), .A(T9453_Y));
KC_INV_X1 T1449 ( .Y(T1449_Y), .A(T1340_Y));
KC_INV_X1 T1430 ( .Y(T1430_Y), .A(T243_Y));
KC_INV_X1 T1386 ( .Y(T1386_Y), .A(T15080_Y));
KC_INV_X1 T1378 ( .Y(T1378_Y), .A(T247_Y));
KC_INV_X1 T1353 ( .Y(T1353_Y), .A(T8990_Y));
KC_INV_X1 T1340 ( .Y(T1340_Y), .A(T8972_Y));
KC_INV_X1 T1339 ( .Y(T1339_Y), .A(T8971_Y));
KC_INV_X1 T1245 ( .Y(T1245_Y), .A(T8924_Y));
KC_INV_X1 T15492 ( .Y(T15492_Y), .A(T9024_Y));
KC_INV_X1 T15490 ( .Y(T15490_Y), .A(T15082_Y));
KC_INV_X1 T15489 ( .Y(T15489_Y), .A(T2242_Y));
KC_INV_X1 T15488 ( .Y(T15488_Y), .A(T16287_Y));
KC_INV_X1 T4818 ( .Y(T4818_Y), .A(T15118_Y));
KC_INV_X1 T4817 ( .Y(T4817_Y), .A(T9174_Y));
KC_INV_X1 T4816 ( .Y(T4816_Y), .A(T9207_Y));
KC_INV_X1 T4801 ( .Y(T4801_Y), .A(T15091_Y));
KC_INV_X1 T4800 ( .Y(T4800_Y), .A(T15150_Y));
KC_INV_X1 T1603 ( .Y(T1603_Y), .A(T9083_Y));
KC_INV_X1 T16478 ( .Y(T16478_Y), .A(T12457_Y));
KC_INV_X1 T265 ( .Y(T265_Y), .A(T277_Q));
KC_INV_X1 T264 ( .Y(T264_Y), .A(T293_Q));
KC_INV_X1 T251 ( .Y(T251_Y), .A(T296_Q));
KC_INV_X1 T15357 ( .Y(T15357_Y), .A(T5226_Q));
KC_INV_X1 T15354 ( .Y(T15354_Y), .A(T6944_Y));
KC_INV_X1 T6465 ( .Y(T6465_Y), .A(T151_Q));
KC_INV_X1 T6471 ( .Y(T6471_Y), .A(T4823_Q));
KC_INV_X1 T954 ( .Y(T954_Y), .A(T5243_Q));
KC_INV_X1 T348 ( .Y(T348_Y), .A(T5562_Q));
KC_INV_X1 T332 ( .Y(T332_Y), .A(T282_Q));
KC_INV_X1 T331 ( .Y(T331_Y), .A(T5241_Q));
KC_INV_X1 T327 ( .Y(T327_Y), .A(T5239_Q));
KC_INV_X1 T321 ( .Y(T321_Y), .A(T289_Q));
KC_INV_X1 T318 ( .Y(T318_Y), .A(T5242_Q));
KC_INV_X1 T15373 ( .Y(T15373_Y), .A(T4822_Q));
KC_INV_X1 T15372 ( .Y(T15372_Y), .A(T5564_Q));
KC_INV_X1 T6608 ( .Y(T6608_Y), .A(T177_Q));
KC_INV_X1 T6603 ( .Y(T6603_Y), .A(T5559_Q));
KC_INV_X1 T6351 ( .Y(T6351_Y), .A(T323_Q));
KC_INV_X1 T399 ( .Y(T399_Y), .A(T5255_Q));
KC_INV_X1 T397 ( .Y(T397_Y), .A(T172_Q));
KC_INV_X1 T396 ( .Y(T396_Y), .A(T171_Q));
KC_INV_X1 T389 ( .Y(T389_Y), .A(T5251_Q));
KC_INV_X1 T386 ( .Y(T386_Y), .A(T316_Q));
KC_INV_X1 T15388 ( .Y(T15388_Y), .A(T169_Q));
KC_INV_X1 T6809 ( .Y(T6809_Y), .A(T684_Y));
KC_INV_X1 T6723 ( .Y(T6723_Y), .A(T319_Q));
KC_INV_X1 T569 ( .Y(T569_Y), .A(T204_Q));
KC_INV_X1 T568 ( .Y(T568_Y), .A(T189_Q));
KC_INV_X1 T535 ( .Y(T535_Y), .A(T191_Q));
KC_INV_X1 T507 ( .Y(T507_Y), .A(T9352_Q));
KC_INV_X1 T506 ( .Y(T506_Y), .A(T184_Q));
KC_INV_X1 T505 ( .Y(T505_Y), .A(T9349_Q));
KC_INV_X1 T6681 ( .Y(T6681_Y), .A(T362_Q));
KC_INV_X1 T797 ( .Y(T797_Y), .A(T7569_Y));
KC_INV_X1 T743 ( .Y(T743_Y), .A(T208_Q));
KC_INV_X1 T740 ( .Y(T740_Y), .A(T8697_Y));
KC_INV_X1 T739 ( .Y(T739_Y), .A(T9388_Y));
KC_INV_X1 T738 ( .Y(T738_Y), .A(T11207_Y));
KC_INV_X1 T682 ( .Y(T682_Y), .A(T16320_Y));
KC_INV_X1 T15429 ( .Y(T15429_Y), .A(T350_Y));
KC_INV_X1 T16331 ( .Y(T16331_Y), .A(T9386_Y));
KC_INV_X1 T16329 ( .Y(T16329_Y), .A(T7827_Y));
KC_INV_X1 T16319 ( .Y(T16319_Y), .A(T7576_Y));
KC_INV_X1 T970 ( .Y(T970_Y), .A(T8137_Y));
KC_INV_X1 T968 ( .Y(T968_Y), .A(T9110_Y));
KC_INV_X1 T967 ( .Y(T967_Y), .A(T8865_Y));
KC_INV_X1 T941 ( .Y(T941_Y), .A(T7582_Y));
KC_INV_X1 T936 ( .Y(T936_Y), .A(T8812_Y));
KC_INV_X1 T924 ( .Y(T924_Y), .A(T9381_Y));
KC_INV_X1 T921 ( .Y(T921_Y), .A(T5354_Q));
KC_INV_X1 T918 ( .Y(T918_Y), .A(T7828_Y));
KC_INV_X1 T917 ( .Y(T917_Y), .A(T9384_Y));
KC_INV_X1 T15655 ( .Y(T15655_Y), .A(T7670_Y));
KC_INV_X1 T15453 ( .Y(T15453_Y), .A(T16480_Q));
KC_INV_X1 T15452 ( .Y(T15452_Y), .A(T7831_Y));
KC_INV_X1 T15451 ( .Y(T15451_Y), .A(T12455_Y));
KC_INV_X1 T1440 ( .Y(T1440_Y), .A(T9092_Y));
KC_INV_X1 T1439 ( .Y(T1439_Y), .A(T9079_Y));
KC_INV_X1 T1438 ( .Y(T1438_Y), .A(T9158_Y));
KC_INV_X1 T1429 ( .Y(T1429_Y), .A(T9093_Y));
KC_INV_X1 T1427 ( .Y(T1427_Y), .A(T16278_Y));
KC_INV_X1 T1354 ( .Y(T1354_Y), .A(T9203_Y));
KC_INV_X1 T1335 ( .Y(T1335_Y), .A(T12723_Y));
KC_INV_X1 T1334 ( .Y(T1334_Y), .A(T8104_Y));
KC_INV_X1 T1321 ( .Y(T1321_Y), .A(T7918_Y));
KC_INV_X1 T1287 ( .Y(T1287_Y), .A(T7902_Y));
KC_INV_X1 T1286 ( .Y(T1286_Y), .A(T8079_Y));
KC_INV_X1 T1284 ( .Y(T1284_Y), .A(T7917_Y));
KC_INV_X1 T1278 ( .Y(T1278_Y), .A(T8101_Y));
KC_INV_X1 T1273 ( .Y(T1273_Y), .A(T8949_Y));
KC_INV_X1 T1272 ( .Y(T1272_Y), .A(T8078_Y));
KC_INV_X1 T1266 ( .Y(T1266_Y), .A(T8103_Y));
KC_INV_X1 T1225 ( .Y(T1225_Y), .A(T7909_Y));
KC_INV_X1 T1217 ( .Y(T1217_Y), .A(T7905_Y));
KC_INV_X1 T1213 ( .Y(T1213_Y), .A(T8100_Y));
KC_INV_X1 T1206 ( .Y(T1206_Y), .A(T8950_Y));
KC_INV_X1 T16191 ( .Y(T16191_Y), .A(T9484_Y));
KC_INV_X1 T2392 ( .Y(T2392_Y), .A(T15092_Y));
KC_INV_X1 T2390 ( .Y(T2390_Y), .A(T15093_Y));
KC_INV_X1 T15524 ( .Y(T15524_Y), .A(T9169_Y));
KC_INV_X1 T15523 ( .Y(T15523_Y), .A(T9168_Y));
KC_INV_X1 T5274 ( .Y(T5274_Y), .A(T9115_Y));
KC_INV_X1 T5228 ( .Y(T5228_Y), .A(T427_Y));
KC_INV_X1 T217 ( .Y(T217_Y), .A(T5193_Q));
KC_INV_X1 T108 ( .Y(T108_Y), .A(T438_Q));
KC_INV_X1 T6313 ( .Y(T6313_Y), .A(T439_Q));
KC_INV_X1 T311 ( .Y(T311_Y), .A(T274_Q));
KC_INV_X1 T250 ( .Y(T250_Y), .A(T5204_Q));
KC_INV_X1 T15352 ( .Y(T15352_Y), .A(T432_Q));
KC_INV_X1 T6348 ( .Y(T6348_Y), .A(T7085_Q));
KC_INV_X1 T347 ( .Y(T347_Y), .A(T160_Q));
KC_INV_X1 T342 ( .Y(T342_Y), .A(T459_Q));
KC_INV_X1 T15371 ( .Y(T15371_Y), .A(T5260_Q));
KC_INV_X1 T6613 ( .Y(T6613_Y), .A(T5253_Q));
KC_INV_X1 T6609 ( .Y(T6609_Y), .A(T320_Q));
KC_INV_X1 T6346 ( .Y(T6346_Y), .A(T281_Q));
KC_INV_X1 T391 ( .Y(T391_Y), .A(T170_Q));
KC_INV_X1 T385 ( .Y(T385_Y), .A(T330_Q));
KC_INV_X1 T381 ( .Y(T381_Y), .A(T672_Q));
KC_INV_X1 T15389 ( .Y(T15389_Y), .A(T5257_Q));
KC_INV_X1 T6713 ( .Y(T6713_Y), .A(T5276_Q));
KC_INV_X1 T6712 ( .Y(T6712_Y), .A(T5560_Q));
KC_INV_X1 T6397 ( .Y(T6397_Y), .A(T190_Q));
KC_INV_X1 T564 ( .Y(T564_Y), .A(T501_Q));
KC_INV_X1 T563 ( .Y(T563_Y), .A(T181_Q));
KC_INV_X1 T562 ( .Y(T562_Y), .A(T341_Q));
KC_INV_X1 T527 ( .Y(T527_Y), .A(T681_Q));
KC_INV_X1 T504 ( .Y(T504_Y), .A(T5304_Q));
KC_INV_X1 T502 ( .Y(T502_Y), .A(T5282_Q));
KC_INV_X1 T499 ( .Y(T499_Y), .A(T9351_Q));
KC_INV_X1 T15412 ( .Y(T15412_Y), .A(T526_Q));
KC_INV_X1 T6671 ( .Y(T6671_Y), .A(T523_Q));
KC_INV_X1 T6670 ( .Y(T6670_Y), .A(T519_Q));
KC_INV_X1 T6662 ( .Y(T6662_Y), .A(T5306_Q));
KC_INV_X1 T794 ( .Y(T794_Y), .A(T8777_Y));
KC_INV_X1 T742 ( .Y(T742_Y), .A(T9111_Y));
KC_INV_X1 T684 ( .Y(T684_Y), .A(T8722_Y));
KC_INV_X1 T642 ( .Y(T642_Y), .A(T7564_Y));
KC_INV_X1 T15434 ( .Y(T15434_Y), .A(T8803_Y));
KC_INV_X1 T16420 ( .Y(T16420_Y), .A(T12368_Y));
KC_INV_X1 T9378 ( .Y(T9378_Y), .A(T5342_Q));
KC_INV_X1 T966 ( .Y(T966_Y), .A(T7901_Y));
KC_INV_X1 T960 ( .Y(T960_Y), .A(T8067_Y));
KC_INV_X1 T933 ( .Y(T933_Y), .A(T9269_Y));
KC_INV_X1 T920 ( .Y(T920_Y), .A(T612_Y));
KC_INV_X1 T916 ( .Y(T916_Y), .A(T9411_Y));
KC_INV_X1 T915 ( .Y(T915_Y), .A(T551_Q));
KC_INV_X1 T914 ( .Y(T914_Y), .A(T541_Q));
KC_INV_X1 T913 ( .Y(T913_Y), .A(T5350_Q));
KC_INV_X1 T16311 ( .Y(T16311_Y), .A(T566_Q));
KC_INV_X1 T1422 ( .Y(T1422_Y), .A(T390_Y));
KC_INV_X1 T1421 ( .Y(T1421_Y), .A(T9418_Y));
KC_INV_X1 T1352 ( .Y(T1352_Y), .A(T561_Q));
KC_INV_X1 T1350 ( .Y(T1350_Y), .A(T556_Q));
KC_INV_X1 T1349 ( .Y(T1349_Y), .A(T8947_Y));
KC_INV_X1 T1328 ( .Y(T1328_Y), .A(T572_Q));
KC_INV_X1 T1214 ( .Y(T1214_Y), .A(T16391_Y));
KC_INV_X1 T1205 ( .Y(T1205_Y), .A(T16310_Y));
KC_INV_X1 T1201 ( .Y(T1201_Y), .A(T9007_Y));
KC_INV_X1 T1200 ( .Y(T1200_Y), .A(T8072_Y));
KC_INV_X1 T1199 ( .Y(T1199_Y), .A(T8945_Y));
KC_INV_X1 T10140 ( .Y(T10140_Y), .A(T9113_Y));
KC_INV_X1 T16184 ( .Y(T16184_Y), .A(T9166_Y));
KC_INV_X1 T16183 ( .Y(T16183_Y), .A(T604_Q));
KC_INV_X1 T4815 ( .Y(T4815_Y), .A(T5406_Q));
KC_INV_X1 T4814 ( .Y(T4814_Y), .A(T605_Q));
KC_INV_X1 T4813 ( .Y(T4813_Y), .A(T606_Q));
KC_INV_X1 T1842 ( .Y(T1842_Y), .A(T606_Q));
KC_INV_X1 T1841 ( .Y(T1841_Y), .A(T9469_Q));
KC_INV_X1 T1599 ( .Y(T1599_Y), .A(T567_Q));
KC_INV_X1 T1594 ( .Y(T1594_Y), .A(T955_Y));
KC_INV_X1 T1593 ( .Y(T1593_Y), .A(T8123_Y));
KC_INV_X1 T168 ( .Y(T168_Y), .A(T9193_Y));
KC_INV_X1 T15540 ( .Y(T15540_Y), .A(T1279_Y));
KC_INV_X1 T15538 ( .Y(T15538_Y), .A(T16507_Y));
KC_INV_X1 T110 ( .Y(T110_Y), .A(T5199_Q));
KC_INV_X1 T109 ( .Y(T109_Y), .A(T12374_Y));
KC_INV_X1 T15331 ( .Y(T15331_Y), .A(T627_Q));
KC_INV_X1 T15171 ( .Y(T15171_Y), .A(T624_Q));
KC_INV_X1 T6304 ( .Y(T6304_Y), .A(T452_Q));
KC_INV_X1 T6300 ( .Y(T6300_Y), .A(T6270_Y));
KC_INV_X1 T6289 ( .Y(T6289_Y), .A(T814_Q));
KC_INV_X1 T6288 ( .Y(T6288_Y), .A(T5195_Q));
KC_INV_X1 T310 ( .Y(T310_Y), .A(T5205_Q));
KC_INV_X1 T302 ( .Y(T302_Y), .A(T12381_Y));
KC_INV_X1 T299 ( .Y(T299_Y), .A(T6919_Y));
KC_INV_X1 T249 ( .Y(T249_Y), .A(T5200_Q));
KC_INV_X1 T246 ( .Y(T246_Y), .A(T449_Q));
KC_INV_X1 T244 ( .Y(T244_Y), .A(T625_Q));
KC_INV_X1 T242 ( .Y(T242_Y), .A(T12385_Y));
KC_INV_X1 T237 ( .Y(T237_Y), .A(T456_Q));
KC_INV_X1 T15355 ( .Y(T15355_Y), .A(T790_Q));
KC_INV_X1 T15350 ( .Y(T15350_Y), .A(T12378_Y));
KC_INV_X1 T15349 ( .Y(T15349_Y), .A(T630_Q));
KC_INV_X1 T6332 ( .Y(T6332_Y), .A(T441_Q));
KC_INV_X1 T6331 ( .Y(T6331_Y), .A(T4846_Q));
KC_INV_X1 T339 ( .Y(T339_Y), .A(T435_Q));
KC_INV_X1 T333 ( .Y(T333_Y), .A(T5206_Q));
KC_INV_X1 T324 ( .Y(T324_Y), .A(T657_Q));
KC_INV_X1 T15648 ( .Y(T15648_Y), .A(T12392_Y));
KC_INV_X1 T15367 ( .Y(T15367_Y), .A(T12394_Y));
KC_INV_X1 T6485 ( .Y(T6485_Y), .A(T5206_Q));
KC_INV_X1 T6699 ( .Y(T6699_Y), .A(T680_Q));
KC_INV_X1 T557 ( .Y(T557_Y), .A(T11885_Y));
KC_INV_X1 T15406 ( .Y(T15406_Y), .A(T712_Q));
KC_INV_X1 T737 ( .Y(T737_Y), .A(T711_Q));
KC_INV_X1 T641 ( .Y(T641_Y), .A(T11886_Y));
KC_INV_X1 T16388 ( .Y(T16388_Y), .A(T8117_Y));
KC_INV_X1 T16387 ( .Y(T16387_Y), .A(T9416_Y));
KC_INV_X1 T944 ( .Y(T944_Y), .A(T11887_Y));
KC_INV_X1 T932 ( .Y(T932_Y), .A(T9001_Y));
KC_INV_X1 T931 ( .Y(T931_Y), .A(T8976_Y));
KC_INV_X1 T928 ( .Y(T928_Y), .A(T7844_Y));
KC_INV_X1 T912 ( .Y(T912_Y), .A(T5348_Q));
KC_INV_X1 T908 ( .Y(T908_Y), .A(T758_Y));
KC_INV_X1 T907 ( .Y(T907_Y), .A(T13241_Q));
KC_INV_X1 T906 ( .Y(T906_Y), .A(T729_Q));
KC_INV_X1 T905 ( .Y(T905_Y), .A(T8939_Y));
KC_INV_X1 T904 ( .Y(T904_Y), .A(T11888_Y));
KC_INV_X1 T902 ( .Y(T902_Y), .A(T7868_Y));
KC_INV_X1 T900 ( .Y(T900_Y), .A(T8805_Y));
KC_INV_X1 T1255 ( .Y(T1255_Y), .A(T9096_Y));
KC_INV_X1 T1198 ( .Y(T1198_Y), .A(T8905_Y));
KC_INV_X1 T209 ( .Y(T209_Y), .A(T209_A));
KC_INV_X1 T192 ( .Y(T192_Y), .A(T185_Y));
KC_INV_X1 T185 ( .Y(T185_Y), .A(T209_Y));
KC_INV_X1 T6290 ( .Y(T6290_Y), .A(T824_Q));
KC_INV_X1 T301 ( .Y(T301_Y), .A(T816_Q));
KC_INV_X1 T245 ( .Y(T245_Y), .A(T793_Q));
KC_INV_X1 T6172 ( .Y(T6172_Y), .A(T671_Q));
KC_INV_X1 T345 ( .Y(T345_Y), .A(T831_Q));
KC_INV_X1 T334 ( .Y(T334_Y), .A(T811_Q));
KC_INV_X1 T317 ( .Y(T317_Y), .A(T813_Q));
KC_INV_X1 T315 ( .Y(T315_Y), .A(T825_Q));
KC_INV_X1 T6638 ( .Y(T6638_Y), .A(T666_Q));
KC_INV_X1 T6630 ( .Y(T6630_Y), .A(T663_Q));
KC_INV_X1 T6629 ( .Y(T6629_Y), .A(T668_Q));
KC_INV_X1 T6625 ( .Y(T6625_Y), .A(T665_Q));
KC_INV_X1 T5938 ( .Y(T5938_Y), .A(T679_Q));
KC_INV_X1 T384 ( .Y(T384_Y), .A(T9301_Y));
KC_INV_X1 T380 ( .Y(T380_Y), .A(T5565_Q));
KC_INV_X1 T379 ( .Y(T379_Y), .A(T4855_Q));
KC_INV_X1 T377 ( .Y(T377_Y), .A(T829_Q));
KC_INV_X1 T15659 ( .Y(T15659_Y), .A(T694_Q));
KC_INV_X1 T15647 ( .Y(T15647_Y), .A(T674_Q));
KC_INV_X1 T15391 ( .Y(T15391_Y), .A(T676_Q));
KC_INV_X1 T15390 ( .Y(T15390_Y), .A(T670_Q));
KC_INV_X1 T15387 ( .Y(T15387_Y), .A(T677_Q));
KC_INV_X1 T6691 ( .Y(T6691_Y), .A(T8758_Y));
KC_INV_X1 T578 ( .Y(T578_Y), .A(T8707_Y));
KC_INV_X1 T577 ( .Y(T577_Y), .A(T7437_Y));
KC_INV_X1 T573 ( .Y(T573_Y), .A(T9334_Y));
KC_INV_X1 T553 ( .Y(T553_Y), .A(T9370_Y));
KC_INV_X1 T552 ( .Y(T552_Y), .A(T7412_Y));
KC_INV_X1 T549 ( .Y(T549_Y), .A(T8762_Y));
KC_INV_X1 T548 ( .Y(T548_Y), .A(T7413_Y));
KC_INV_X1 T547 ( .Y(T547_Y), .A(T896_Y));
KC_INV_X1 T546 ( .Y(T546_Y), .A(T7415_Y));
KC_INV_X1 T545 ( .Y(T545_Y), .A(T7414_Y));
KC_INV_X1 T542 ( .Y(T542_Y), .A(T7363_Y));
KC_INV_X1 T497 ( .Y(T497_Y), .A(T9360_Y));
KC_INV_X1 T15650 ( .Y(T15650_Y), .A(T9303_Y));
KC_INV_X1 T15413 ( .Y(T15413_Y), .A(T692_Y));
KC_INV_X1 T15408 ( .Y(T15408_Y), .A(T8670_Y));
KC_INV_X1 T16163 ( .Y(T16163_Y), .A(T7591_Y));
KC_INV_X1 T6659 ( .Y(T6659_Y), .A(T9331_Y));
KC_INV_X1 T6650 ( .Y(T6650_Y), .A(T7553_Y));
KC_INV_X1 T791 ( .Y(T791_Y), .A(T8771_Y));
KC_INV_X1 T786 ( .Y(T786_Y), .A(T7867_Y));
KC_INV_X1 T783 ( .Y(T783_Y), .A(T8828_Y));
KC_INV_X1 T764 ( .Y(T764_Y), .A(T8792_Y));
KC_INV_X1 T763 ( .Y(T763_Y), .A(T8831_Y));
KC_INV_X1 T755 ( .Y(T755_Y), .A(T8770_Y));
KC_INV_X1 T744 ( .Y(T744_Y), .A(T8763_Y));
KC_INV_X1 T731 ( .Y(T731_Y), .A(T15840_Y));
KC_INV_X1 T728 ( .Y(T728_Y), .A(T15839_Y));
KC_INV_X1 T727 ( .Y(T727_Y), .A(T9359_Y));
KC_INV_X1 T726 ( .Y(T726_Y), .A(T7561_Y));
KC_INV_X1 T719 ( .Y(T719_Y), .A(T7635_Y));
KC_INV_X1 T703 ( .Y(T703_Y), .A(T7618_Y));
KC_INV_X1 T702 ( .Y(T702_Y), .A(T9312_Y));
KC_INV_X1 T700 ( .Y(T700_Y), .A(T7560_Y));
KC_INV_X1 T660 ( .Y(T660_Y), .A(T7590_Y));
KC_INV_X1 T652 ( .Y(T652_Y), .A(T15223_Y));
KC_INV_X1 T651 ( .Y(T651_Y), .A(T9313_Y));
KC_INV_X1 T639 ( .Y(T639_Y), .A(T934_Y));
KC_INV_X1 T638 ( .Y(T638_Y), .A(T16092_Y));
KC_INV_X1 T637 ( .Y(T637_Y), .A(T9362_Y));
KC_INV_X1 T636 ( .Y(T636_Y), .A(T910_Q));
KC_INV_X1 T15432 ( .Y(T15432_Y), .A(T7683_Y));
KC_INV_X1 T15431 ( .Y(T15431_Y), .A(T7614_Y));
KC_INV_X1 T15428 ( .Y(T15428_Y), .A(T5302_Y));
KC_INV_X1 T15841 ( .Y(T15841_Y), .A(T7845_Y));
KC_INV_X1 T16421 ( .Y(T16421_Y), .A(T8936_Y));
KC_INV_X1 T951 ( .Y(T951_Y), .A(T7878_Y));
KC_INV_X1 T950 ( .Y(T950_Y), .A(T7846_Y));
KC_INV_X1 T948 ( .Y(T948_Y), .A(T938_Q));
KC_INV_X1 T947 ( .Y(T947_Y), .A(T940_Q));
KC_INV_X1 T926 ( .Y(T926_Y), .A(T13201_Y));
KC_INV_X1 T925 ( .Y(T925_Y), .A(T7841_Y));
KC_INV_X1 T903 ( .Y(T903_Y), .A(T1247_Q));
KC_INV_X1 T15654 ( .Y(T15654_Y), .A(T8829_Y));
KC_INV_X1 T15458 ( .Y(T15458_Y), .A(T939_Q));
KC_INV_X1 T15457 ( .Y(T15457_Y), .A(T981_Q));
KC_INV_X1 T15454 ( .Y(T15454_Y), .A(T7839_Y));
KC_INV_X1 T1395 ( .Y(T1395_Y), .A(T9000_Y));
KC_INV_X1 T1346 ( .Y(T1346_Y), .A(T140_Y));
KC_INV_X1 T1342 ( .Y(T1342_Y), .A(T10660_Y));
KC_INV_X1 T1197 ( .Y(T1197_Y), .A(T965_Y));
KC_INV_X1 T1196 ( .Y(T1196_Y), .A(T16006_Y));
KC_INV_X1 T15487 ( .Y(T15487_Y), .A(T9998_Y));
KC_INV_X1 T15486 ( .Y(T15486_Y), .A(T1134_Y));
KC_INV_X1 T15485 ( .Y(T15485_Y), .A(T16006_Y));
KC_INV_X1 T1551 ( .Y(T1551_Y), .A(T1012_Q));
KC_INV_X1 T15520 ( .Y(T15520_Y), .A(T8093_Y));
KC_INV_X1 T383 ( .Y(T383_Y), .A(T5297_Q));
KC_INV_X1 T6822 ( .Y(T6822_Y), .A(T8716_Y));
KC_INV_X1 T6651 ( .Y(T6651_Y), .A(T10344_Y));
KC_INV_X1 T596 ( .Y(T596_Y), .A(T15777_Y));
KC_INV_X1 T585 ( .Y(T585_Y), .A(T8727_Y));
KC_INV_X1 T515 ( .Y(T515_Y), .A(T8717_Y));
KC_INV_X1 T514 ( .Y(T514_Y), .A(T8683_Y));
KC_INV_X1 T498 ( .Y(T498_Y), .A(T7592_Y));
KC_INV_X1 T15751 ( .Y(T15751_Y), .A(T15779_Y));
KC_INV_X1 T15750 ( .Y(T15750_Y), .A(T10345_Y));
KC_INV_X1 T718 ( .Y(T718_Y), .A(T1084_Q));
KC_INV_X1 T715 ( .Y(T715_Y), .A(T7636_Y));
KC_INV_X1 T658 ( .Y(T658_Y), .A(T9332_Y));
KC_INV_X1 T656 ( .Y(T656_Y), .A(T15773_Y));
KC_INV_X1 T15665 ( .Y(T15665_Y), .A(T15776_Y));
KC_INV_X1 T15440 ( .Y(T15440_Y), .A(T7799_Y));
KC_INV_X1 T15433 ( .Y(T15433_Y), .A(T5310_Q));
KC_INV_X1 T16401 ( .Y(T16401_Y), .A(T10331_Y));
KC_INV_X1 T16394 ( .Y(T16394_Y), .A(T1128_Q));
KC_INV_X1 T16384 ( .Y(T16384_Y), .A(T8800_Y));
KC_INV_X1 T16381 ( .Y(T16381_Y), .A(T5561_Q));
KC_INV_X1 T1062 ( .Y(T1062_Y), .A(T8781_Y));
KC_INV_X1 T1050 ( .Y(T1050_Y), .A(T378_Y));
KC_INV_X1 T1042 ( .Y(T1042_Y), .A(T8783_Y));
KC_INV_X1 T1009 ( .Y(T1009_Y), .A(T1113_Q));
KC_INV_X1 T1008 ( .Y(T1008_Y), .A(T1094_Q));
KC_INV_X1 T1007 ( .Y(T1007_Y), .A(T9891_Y));
KC_INV_X1 T987 ( .Y(T987_Y), .A(T5334_Q));
KC_INV_X1 T986 ( .Y(T986_Y), .A(T10316_Y));
KC_INV_X1 T946 ( .Y(T946_Y), .A(T1130_Q));
KC_INV_X1 T927 ( .Y(T927_Y), .A(T1131_Q));
KC_INV_X1 T15664 ( .Y(T15664_Y), .A(T1100_Q));
KC_INV_X1 T15466 ( .Y(T15466_Y), .A(T16422_Q));
KC_INV_X1 T15461 ( .Y(T15461_Y), .A(T540_Y));
KC_INV_X1 T15455 ( .Y(T15455_Y), .A(T12444_Y));
KC_INV_X1 T1481 ( .Y(T1481_Y), .A(T10048_Y));
KC_INV_X1 T1469 ( .Y(T1469_Y), .A(T10169_Y));
KC_INV_X1 T1458 ( .Y(T1458_Y), .A(T10004_Y));
KC_INV_X1 T1457 ( .Y(T1457_Y), .A(T1135_Q));
KC_INV_X1 T1394 ( .Y(T1394_Y), .A(T10298_Y));
KC_INV_X1 T1246 ( .Y(T1246_Y), .A(T10008_Y));
KC_INV_X1 T15500 ( .Y(T15500_Y), .A(T1130_Q));
KC_INV_X1 T15497 ( .Y(T15497_Y), .A(T1129_Q));
KC_INV_X1 T9056 ( .Y(T9056_Y), .A(T10175_Y));
KC_INV_X1 T4848 ( .Y(T4848_Y), .A(T10299_Y));
KC_INV_X1 T16414 ( .Y(T16414_Y), .A(T5373_Q));
KC_INV_X1 T16393 ( .Y(T16393_Y), .A(T10044_Y));
KC_INV_X1 T16377 ( .Y(T16377_Y), .A(T9899_Y));
KC_INV_X1 T1089 ( .Y(T1089_Y), .A(T1204_Q));
KC_INV_X1 T1086 ( .Y(T1086_Y), .A(T10328_Y));
KC_INV_X1 T1085 ( .Y(T1085_Y), .A(T7845_Y));
KC_INV_X1 T1060 ( .Y(T1060_Y), .A(T1209_Q));
KC_INV_X1 T1059 ( .Y(T1059_Y), .A(T11011_Y));
KC_INV_X1 T15472 ( .Y(T15472_Y), .A(T9898_Y));
KC_INV_X1 T15471 ( .Y(T15471_Y), .A(T1191_Q));
KC_INV_X1 T15464 ( .Y(T15464_Y), .A(T10329_Y));
KC_INV_X1 T15463 ( .Y(T15463_Y), .A(T10916_Y));
KC_INV_X1 T16308 ( .Y(T16308_Y), .A(T5375_Q));
KC_INV_X1 T4847 ( .Y(T4847_Y), .A(T10130_Y));
KC_INV_X1 T4838 ( .Y(T4838_Y), .A(T10139_Y));
KC_INV_X1 T4831 ( .Y(T4831_Y), .A(T5814_Y));
KC_INV_X1 T4819 ( .Y(T4819_Y), .A(T1281_Y));
KC_INV_X1 T15527 ( .Y(T15527_Y), .A(T1358_Y));
KC_INV_X1 T5382 ( .Y(T5382_Y), .A(T13056_Q));
KC_INV_X1 T5381 ( .Y(T5381_Y), .A(T13059_Q));
KC_INV_X1 T372 ( .Y(T372_Y), .A(T7236_Y));
KC_INV_X1 T367 ( .Y(T367_Y), .A(T7235_Y));
KC_INV_X1 T361 ( .Y(T361_Y), .A(T14980_Y));
KC_INV_X1 T356 ( .Y(T356_Y), .A(T7182_Y));
KC_INV_X1 T355 ( .Y(T355_Y), .A(T7233_Y));
KC_INV_X1 T15378 ( .Y(T15378_Y), .A(T7351_Y));
KC_INV_X1 T6748 ( .Y(T6748_Y), .A(T7339_Y));
KC_INV_X1 T6747 ( .Y(T6747_Y), .A(T1338_Y));
KC_INV_X1 T15677 ( .Y(T15677_Y), .A(T5674_Y));
KC_INV_X1 T852 ( .Y(T852_Y), .A(T7776_Y));
KC_INV_X1 T1083 ( .Y(T1083_Y), .A(T10037_Y));
KC_INV_X1 T1082 ( .Y(T1082_Y), .A(T7975_Y));
KC_INV_X1 T15470 ( .Y(T15470_Y), .A(T7942_Y));
KC_INV_X1 T4825 ( .Y(T4825_Y), .A(T10725_Y));
KC_INV_X1 T15543 ( .Y(T15543_Y), .A(T6431_Q));
KC_INV_X1 T370 ( .Y(T370_Y), .A(T7017_Y));
KC_INV_X1 T369 ( .Y(T369_Y), .A(T6984_Y));
KC_INV_X1 T366 ( .Y(T366_Y), .A(T7026_Y));
KC_INV_X1 T365 ( .Y(T365_Y), .A(T7160_Y));
KC_INV_X1 T364 ( .Y(T364_Y), .A(T7151_Y));
KC_INV_X1 T358 ( .Y(T358_Y), .A(T7227_Y));
KC_INV_X1 T354 ( .Y(T354_Y), .A(T7159_Y));
KC_INV_X1 T353 ( .Y(T353_Y), .A(T6997_Y));
KC_INV_X1 T351 ( .Y(T351_Y), .A(T7232_Y));
KC_INV_X1 T15671 ( .Y(T15671_Y), .A(T7219_Y));
KC_INV_X1 T15670 ( .Y(T15670_Y), .A(T7703_Y));
KC_INV_X1 T15379 ( .Y(T15379_Y), .A(T7036_Y));
KC_INV_X1 T15375 ( .Y(T15375_Y), .A(T10391_Y));
KC_INV_X1 T6749 ( .Y(T6749_Y), .A(T5696_Y));
KC_INV_X1 T6468 ( .Y(T6468_Y), .A(T7010_Y));
KC_INV_X1 T403 ( .Y(T403_Y), .A(T7337_Y));
KC_INV_X1 T402 ( .Y(T402_Y), .A(T5701_Y));
KC_INV_X1 T401 ( .Y(T401_Y), .A(T7496_Y));
KC_INV_X1 T15676 ( .Y(T15676_Y), .A(T10373_Y));
KC_INV_X1 T15395 ( .Y(T15395_Y), .A(T5681_Y));
KC_INV_X1 T15393 ( .Y(T15393_Y), .A(T7703_Y));
KC_INV_X1 T589 ( .Y(T589_Y), .A(T7548_Y));
KC_INV_X1 T587 ( .Y(T587_Y), .A(T5695_Y));
KC_INV_X1 T853 ( .Y(T853_Y), .A(T7738_Y));
KC_INV_X1 T851 ( .Y(T851_Y), .A(T10338_Y));
KC_INV_X1 T827 ( .Y(T827_Y), .A(T7739_Y));
KC_INV_X1 T821 ( .Y(T821_Y), .A(T7717_Y));
KC_INV_X1 T15439 ( .Y(T15439_Y), .A(T9790_Y));
KC_INV_X1 T15436 ( .Y(T15436_Y), .A(T7711_Y));
KC_INV_X1 T16440 ( .Y(T16440_Y), .A(T10917_Y));
KC_INV_X1 T16399 ( .Y(T16399_Y), .A(T7991_Y));
KC_INV_X1 T1080 ( .Y(T1080_Y), .A(T7935_Y));
KC_INV_X1 T1058 ( .Y(T1058_Y), .A(T10907_Y));
KC_INV_X1 T1038 ( .Y(T1038_Y), .A(T10012_Y));
KC_INV_X1 T1035 ( .Y(T1035_Y), .A(T7934_Y));
KC_INV_X1 T1033 ( .Y(T1033_Y), .A(T9997_Y));
KC_INV_X1 T1027 ( .Y(T1027_Y), .A(T9999_Y));
KC_INV_X1 T15660 ( .Y(T15660_Y), .A(T11010_Y));
KC_INV_X1 T15468 ( .Y(T15468_Y), .A(T7928_Y));
KC_INV_X1 T1472 ( .Y(T1472_Y), .A(T10883_Y));
KC_INV_X1 T292 ( .Y(T292_Y), .A(T1521_Y));
KC_INV_X1 T15396 ( .Y(T15396_Y), .A(T5662_Y));
KC_INV_X1 T15392 ( .Y(T15392_Y), .A(T7320_Y));
KC_INV_X1 T6789 ( .Y(T6789_Y), .A(T5650_Y));
KC_INV_X1 T835 ( .Y(T835_Y), .A(T9781_Y));
KC_INV_X1 T15435 ( .Y(T15435_Y), .A(T3656_Y));
KC_INV_X1 T15462 ( .Y(T15462_Y), .A(T10239_Y));
KC_INV_X1 T16437 ( .Y(T16437_Y), .A(T10239_Y));
KC_INV_X1 T1079 ( .Y(T1079_Y), .A(T10310_Y));
KC_INV_X1 T1055 ( .Y(T1055_Y), .A(T16464_Q));
KC_INV_X1 T1054 ( .Y(T1054_Y), .A(T8004_Y));
KC_INV_X1 T1026 ( .Y(T1026_Y), .A(T9992_Y));
KC_INV_X1 T975 ( .Y(T975_Y), .A(T13082_Y));
KC_INV_X1 T15469 ( .Y(T15469_Y), .A(T16410_Q));
KC_INV_X1 T15467 ( .Y(T15467_Y), .A(T16409_Q));
KC_INV_X1 T1479 ( .Y(T1479_Y), .A(T8002_Y));
KC_INV_X1 T1471 ( .Y(T1471_Y), .A(T10906_Y));
KC_INV_X1 T1450 ( .Y(T1450_Y), .A(T11016_Y));
KC_INV_X1 T6462 ( .Y(T6462_Y), .A(T7334_Y));
KC_INV_X1 T6753 ( .Y(T6753_Y), .A(T14940_Q));
KC_INV_X1 T6752 ( .Y(T6752_Y), .A(T13732_Q));
KC_INV_X1 T6751 ( .Y(T6751_Y), .A(T14739_Q));
KC_INV_X1 T496 ( .Y(T496_Y), .A(T6989_Y));
KC_INV_X1 T494 ( .Y(T494_Y), .A(T14769_Q));
KC_INV_X1 T461 ( .Y(T461_Y), .A(T14773_Q));
KC_INV_X1 T458 ( .Y(T458_Y), .A(T13777_Q));
KC_INV_X1 T457 ( .Y(T457_Y), .A(T7185_Y));
KC_INV_X1 T417 ( .Y(T417_Y), .A(T10399_Y));
KC_INV_X1 T15693 ( .Y(T15693_Y), .A(T14941_Q));
KC_INV_X1 T15675 ( .Y(T15675_Y), .A(T6594_Q));
KC_INV_X1 T15401 ( .Y(T15401_Y), .A(T7347_Y));
KC_INV_X1 T16192 ( .Y(T16192_Y), .A(T1687_Y));
KC_INV_X1 T844 ( .Y(T844_Y), .A(T2539_Y));
KC_INV_X1 T809 ( .Y(T809_Y), .A(T1661_Q));
KC_INV_X1 T803 ( .Y(T803_Y), .A(T16231_Q));
KC_INV_X1 T16436 ( .Y(T16436_Y), .A(T16468_Q));
KC_INV_X1 T16374 ( .Y(T16374_Y), .A(T8877_Q));
KC_INV_X1 T16372 ( .Y(T16372_Y), .A(T1717_Q));
KC_INV_X1 T1192 ( .Y(T1192_Y), .A(T1707_Q));
KC_INV_X1 T1148 ( .Y(T1148_Y), .A(T16433_Q));
KC_INV_X1 T1107 ( .Y(T1107_Y), .A(T1690_Q));
KC_INV_X1 T1057 ( .Y(T1057_Y), .A(T4921_Y));
KC_INV_X1 T1456 ( .Y(T1456_Y), .A(T10905_Y));
KC_INV_X1 T15519 ( .Y(T15519_Y), .A(T5390_Q));
KC_INV_X1 T15515 ( .Y(T15515_Y), .A(T2051_Q));
KC_INV_X1 T4902 ( .Y(T4902_Y), .A(T12982_Y));
KC_INV_X1 T15531 ( .Y(T15531_Y), .A(T10918_Y));
KC_INV_X1 T15529 ( .Y(T15529_Y), .A(T13121_Y));
KC_INV_X1 T15858 ( .Y(T15858_Y), .A(T15809_Q));
KC_INV_X1 T15857 ( .Y(T15857_Y), .A(T16088_Q));
KC_INV_X1 T15856 ( .Y(T15856_Y), .A(T15808_Q));
KC_INV_X1 T15855 ( .Y(T15855_Y), .A(T15796_Q));
KC_INV_X1 T15854 ( .Y(T15854_Y), .A(T16299_Q));
KC_INV_X1 T16474 ( .Y(T16474_Y), .A(T15005_Y));
KC_INV_X1 T5814 ( .Y(T5814_Y), .A(T8335_Y));
KC_INV_X1 T5794 ( .Y(T5794_Y), .A(T10225_Y));
KC_INV_X1 T5945 ( .Y(T5945_Y), .A(T2150_Q));
KC_INV_X1 T5928 ( .Y(T5928_Y), .A(T11530_Y));
KC_INV_X1 T5911 ( .Y(T5911_Y), .A(T1770_Y));
KC_INV_X1 T5903 ( .Y(T5903_Y), .A(T5452_Q));
KC_INV_X1 T15989 ( .Y(T15989_Y), .A(T3415_Y));
KC_INV_X1 T5966 ( .Y(T5966_Y), .A(T1774_Q));
KC_INV_X1 T16017 ( .Y(T16017_Y), .A(T8352_Q));
KC_INV_X1 T6005 ( .Y(T6005_Y), .A(T1807_Q));
KC_INV_X1 T6164 ( .Y(T6164_Y), .A(T6121_Y));
KC_INV_X1 T6125 ( .Y(T6125_Y), .A(T1821_Q));
KC_INV_X1 T15618 ( .Y(T15618_Y), .A(T12269_Y));
KC_INV_X1 T6201 ( .Y(T6201_Y), .A(T2958_Y));
KC_INV_X1 T6199 ( .Y(T6199_Y), .A(T2399_Y));
KC_INV_X1 T15332 ( .Y(T15332_Y), .A(T11753_Y));
KC_INV_X1 T6543 ( .Y(T6543_Y), .A(T1857_Q));
KC_INV_X1 T6542 ( .Y(T6542_Y), .A(T11775_Y));
KC_INV_X1 T6498 ( .Y(T6498_Y), .A(T1856_Q));
KC_INV_X1 T6496 ( .Y(T6496_Y), .A(T8434_Y));
KC_INV_X1 T6495 ( .Y(T6495_Y), .A(T11047_Y));
KC_INV_X1 T6494 ( .Y(T6494_Y), .A(T2400_Y));
KC_INV_X1 T6459 ( .Y(T6459_Y), .A(T1621_Y));
KC_INV_X1 T6756 ( .Y(T6756_Y), .A(T14934_Q));
KC_INV_X1 T6593 ( .Y(T6593_Y), .A(T12569_Y));
KC_INV_X1 T6460 ( .Y(T6460_Y), .A(T1885_Y));
KC_INV_X1 T493 ( .Y(T493_Y), .A(T1628_Y));
KC_INV_X1 T491 ( .Y(T491_Y), .A(T13776_Q));
KC_INV_X1 T490 ( .Y(T490_Y), .A(T13774_Q));
KC_INV_X1 T487 ( .Y(T487_Y), .A(T1913_Y));
KC_INV_X1 T485 ( .Y(T485_Y), .A(T13758_Q));
KC_INV_X1 T484 ( .Y(T484_Y), .A(T1899_Y));
KC_INV_X1 T451 ( .Y(T451_Y), .A(T14939_Q));
KC_INV_X1 T448 ( .Y(T448_Y), .A(T10386_Y));
KC_INV_X1 T410 ( .Y(T410_Y), .A(T1892_Y));
KC_INV_X1 T409 ( .Y(T409_Y), .A(T14771_Q));
KC_INV_X1 T407 ( .Y(T407_Y), .A(T13746_Q));
KC_INV_X1 T15692 ( .Y(T15692_Y), .A(T14840_Q));
KC_INV_X1 T15405 ( .Y(T15405_Y), .A(T6980_Y));
KC_INV_X1 T15400 ( .Y(T15400_Y), .A(T13771_Q));
KC_INV_X1 T15399 ( .Y(T15399_Y), .A(T13775_Q));
KC_INV_X1 T15398 ( .Y(T15398_Y), .A(T4937_Y));
KC_INV_X1 T6783 ( .Y(T6783_Y), .A(T10352_Y));
KC_INV_X1 T6782 ( .Y(T6782_Y), .A(T13896_Q));
KC_INV_X1 T6781 ( .Y(T6781_Y), .A(T1941_Y));
KC_INV_X1 T6775 ( .Y(T6775_Y), .A(T14932_Q));
KC_INV_X1 T635 ( .Y(T635_Y), .A(T4983_Y));
KC_INV_X1 T629 ( .Y(T629_Y), .A(T10334_Y));
KC_INV_X1 T623 ( .Y(T623_Y), .A(T1645_Y));
KC_INV_X1 T15685 ( .Y(T15685_Y), .A(T7481_Y));
KC_INV_X1 T15684 ( .Y(T15684_Y), .A(T1939_Y));
KC_INV_X1 T15421 ( .Y(T15421_Y), .A(T1648_Y));
KC_INV_X1 T16169 ( .Y(T16169_Y), .A(T13020_Q));
KC_INV_X1 T868 ( .Y(T868_Y), .A(T2005_Q));
KC_INV_X1 T16406 ( .Y(T16406_Y), .A(T5320_Q));
KC_INV_X1 T16378 ( .Y(T16378_Y), .A(T2015_Q));
KC_INV_X1 T16369 ( .Y(T16369_Y), .A(T5367_Y));
KC_INV_X1 T16368 ( .Y(T16368_Y), .A(T5363_Q));
KC_INV_X1 T1162 ( .Y(T1162_Y), .A(T1998_Y));
KC_INV_X1 T1142 ( .Y(T1142_Y), .A(T2008_Q));
KC_INV_X1 T1124 ( .Y(T1124_Y), .A(T9949_Y));
KC_INV_X1 T1123 ( .Y(T1123_Y), .A(T2024_Y));
KC_INV_X1 T1119 ( .Y(T1119_Y), .A(T12330_Y));
KC_INV_X1 T1118 ( .Y(T1118_Y), .A(T10524_Y));
KC_INV_X1 T1117 ( .Y(T1117_Y), .A(T2028_Q));
KC_INV_X1 T1116 ( .Y(T1116_Y), .A(T2016_Q));
KC_INV_X1 T1106 ( .Y(T1106_Y), .A(T11949_Y));
KC_INV_X1 T15478 ( .Y(T15478_Y), .A(T2023_Q));
KC_INV_X1 T15474 ( .Y(T15474_Y), .A(T15154_Y));
KC_INV_X1 T16295 ( .Y(T16295_Y), .A(T2061_Y));
KC_INV_X1 T1548 ( .Y(T1548_Y), .A(T5389_Q));
KC_INV_X1 T1533 ( .Y(T1533_Y), .A(T5391_Q));
KC_INV_X1 T1532 ( .Y(T1532_Y), .A(T2012_Q));
KC_INV_X1 T1527 ( .Y(T1527_Y), .A(T5388_Q));
KC_INV_X1 T1519 ( .Y(T1519_Y), .A(T1735_Q));
KC_INV_X1 T1518 ( .Y(T1518_Y), .A(T16305_Y));
KC_INV_X1 T1517 ( .Y(T1517_Y), .A(T2053_Q));
KC_INV_X1 T1509 ( .Y(T1509_Y), .A(T2550_Y));
KC_INV_X1 T1506 ( .Y(T1506_Y), .A(T13042_Q));
KC_INV_X1 T1496 ( .Y(T1496_Y), .A(T2040_Y));
KC_INV_X1 T1495 ( .Y(T1495_Y), .A(T10068_Y));
KC_INV_X1 T1485 ( .Y(T1485_Y), .A(T8394_Y));
KC_INV_X1 T15512 ( .Y(T15512_Y), .A(T1736_Q));
KC_INV_X1 T15511 ( .Y(T15511_Y), .A(T2002_Q));
KC_INV_X1 T15506 ( .Y(T15506_Y), .A(T13032_Y));
KC_INV_X1 T16237 ( .Y(T16237_Y), .A(T12651_Y));
KC_INV_X1 T4868 ( .Y(T4868_Y), .A(T13131_Y));
KC_INV_X1 T15534 ( .Y(T15534_Y), .A(T2069_Y));
KC_INV_X1 T10245 ( .Y(T10245_Y), .A(T15804_Q));
KC_INV_X1 T5745 ( .Y(T5745_Y), .A(T5577_Q));
KC_INV_X1 T5731 ( .Y(T5731_Y), .A(T8484_Y));
KC_INV_X1 T5759 ( .Y(T5759_Y), .A(T15860_Q));
KC_INV_X1 T15882 ( .Y(T15882_Y), .A(T964_Q));
KC_INV_X1 T15881 ( .Y(T15881_Y), .A(T15797_Q));
KC_INV_X1 T5834 ( .Y(T5834_Y), .A(T15891_Q));
KC_INV_X1 T5833 ( .Y(T5833_Y), .A(T2114_Q));
KC_INV_X1 T5820 ( .Y(T5820_Y), .A(T12165_Y));
KC_INV_X1 T5793 ( .Y(T5793_Y), .A(T8448_Y));
KC_INV_X1 T15906 ( .Y(T15906_Y), .A(T4177_Y));
KC_INV_X1 T5848 ( .Y(T5848_Y), .A(T10933_Y));
KC_INV_X1 T15574 ( .Y(T15574_Y), .A(T11480_Y));
KC_INV_X1 T15942 ( .Y(T15942_Y), .A(T8238_Y));
KC_INV_X1 T5944 ( .Y(T5944_Y), .A(T11025_Y));
KC_INV_X1 T5943 ( .Y(T5943_Y), .A(T8316_Y));
KC_INV_X1 T5927 ( .Y(T5927_Y), .A(T15138_Q));
KC_INV_X1 T5926 ( .Y(T5926_Y), .A(T2183_Y));
KC_INV_X1 T5909 ( .Y(T5909_Y), .A(T10932_Y));
KC_INV_X1 T5908 ( .Y(T5908_Y), .A(T11499_Y));
KC_INV_X1 T5902 ( .Y(T5902_Y), .A(T15990_Q));
KC_INV_X1 T5898 ( .Y(T5898_Y), .A(T5461_Q));
KC_INV_X1 T5878 ( .Y(T5878_Y), .A(T16023_Q));
KC_INV_X1 T5991 ( .Y(T5991_Y), .A(T2275_Q));
KC_INV_X1 T5990 ( .Y(T5990_Y), .A(T2802_Y));
KC_INV_X1 T5983 ( .Y(T5983_Y), .A(T2809_Q));
KC_INV_X1 T5982 ( .Y(T5982_Y), .A(T16018_Q));
KC_INV_X1 T5967 ( .Y(T5967_Y), .A(T2217_Y));
KC_INV_X1 T16009 ( .Y(T16009_Y), .A(T11566_Y));
KC_INV_X1 T6028 ( .Y(T6028_Y), .A(T2316_Q));
KC_INV_X1 T6026 ( .Y(T6026_Y), .A(T2236_Q));
KC_INV_X1 T6004 ( .Y(T6004_Y), .A(T16007_Q));
KC_INV_X1 T6003 ( .Y(T6003_Y), .A(T5002_Y));
KC_INV_X1 T6000 ( .Y(T6000_Y), .A(T11727_Y));
KC_INV_X1 T15611 ( .Y(T15611_Y), .A(T2345_Q));
KC_INV_X1 T15608 ( .Y(T15608_Y), .A(T13152_Y));
KC_INV_X1 T16042 ( .Y(T16042_Y), .A(T5571_Q));
KC_INV_X1 T16041 ( .Y(T16041_Y), .A(T2278_Q));
KC_INV_X1 T6073 ( .Y(T6073_Y), .A(T11032_Y));
KC_INV_X1 T6040 ( .Y(T6040_Y), .A(T5481_Q));
KC_INV_X1 T6185 ( .Y(T6185_Y), .A(T4965_Y));
KC_INV_X1 T6162 ( .Y(T6162_Y), .A(T1285_Y));
KC_INV_X1 T6147 ( .Y(T6147_Y), .A(T3482_Y));
KC_INV_X1 T6101 ( .Y(T6101_Y), .A(T12102_Y));
KC_INV_X1 T16131 ( .Y(T16131_Y), .A(T12105_Y));
KC_INV_X1 T6571 ( .Y(T6571_Y), .A(T10573_Y));
KC_INV_X1 T4962 ( .Y(T4962_Y), .A(T6611_S));
KC_INV_X1 T6243 ( .Y(T6243_Y), .A(T10998_Y));
KC_INV_X1 T6232 ( .Y(T6232_Y), .A(T5517_Y));
KC_INV_X1 T6229 ( .Y(T6229_Y), .A(T10557_Y));
KC_INV_X1 T6227 ( .Y(T6227_Y), .A(T11766_Y));
KC_INV_X1 T6198 ( .Y(T6198_Y), .A(T5527_Q));
KC_INV_X1 T6197 ( .Y(T6197_Y), .A(T10997_Y));
KC_INV_X1 T291 ( .Y(T291_Y), .A(T5529_Q));
KC_INV_X1 T15712 ( .Y(T15712_Y), .A(T12108_Y));
KC_INV_X1 T15638 ( .Y(T15638_Y), .A(T2255_Y));
KC_INV_X1 T15633 ( .Y(T15633_Y), .A(T16270_Y));
KC_INV_X1 T15628 ( .Y(T15628_Y), .A(T2326_Y));
KC_INV_X1 T6541 ( .Y(T6541_Y), .A(T2388_Q));
KC_INV_X1 T6540 ( .Y(T6540_Y), .A(T6162_Y));
KC_INV_X1 T6502 ( .Y(T6502_Y), .A(T8432_Y));
KC_INV_X1 T6500 ( .Y(T6500_Y), .A(T2369_Y));
KC_INV_X1 T6499 ( .Y(T6499_Y), .A(T2338_Y));
KC_INV_X1 T6492 ( .Y(T6492_Y), .A(T11034_Y));
KC_INV_X1 T6491 ( .Y(T6491_Y), .A(T5489_Y));
KC_INV_X1 T15646 ( .Y(T15646_Y), .A(T15645_Y));
KC_INV_X1 T15645 ( .Y(T15645_Y), .A(T16473_Y));
KC_INV_X1 T6457 ( .Y(T6457_Y), .A(T13654_Q));
KC_INV_X1 T376 ( .Y(T376_Y), .A(T1620_Y));
KC_INV_X1 T375 ( .Y(T375_Y), .A(T3579_Y));
KC_INV_X1 T15384 ( .Y(T15384_Y), .A(T2973_Y));
KC_INV_X1 T6760 ( .Y(T6760_Y), .A(T2449_Y));
KC_INV_X1 T6758 ( .Y(T6758_Y), .A(T14935_Q));
KC_INV_X1 T6757 ( .Y(T6757_Y), .A(T14839_Q));
KC_INV_X1 T6592 ( .Y(T6592_Y), .A(T4937_Y));
KC_INV_X1 T6458 ( .Y(T6458_Y), .A(T13655_Q));
KC_INV_X1 T6456 ( .Y(T6456_Y), .A(T5033_Y));
KC_INV_X1 T488 ( .Y(T488_Y), .A(T5208_Y));
KC_INV_X1 T477 ( .Y(T477_Y), .A(T13770_Q));
KC_INV_X1 T444 ( .Y(T444_Y), .A(T13772_Q));
KC_INV_X1 T437 ( .Y(T437_Y), .A(T13773_Q));
KC_INV_X1 T418 ( .Y(T418_Y), .A(T13769_Q));
KC_INV_X1 T416 ( .Y(T416_Y), .A(T2447_Y));
KC_INV_X1 T414 ( .Y(T414_Y), .A(T2447_Y));
KC_INV_X1 T411 ( .Y(T411_Y), .A(T14928_Q));
KC_INV_X1 T406 ( .Y(T406_Y), .A(T13783_Q));
KC_INV_X1 T405 ( .Y(T405_Y), .A(T1914_Y));
KC_INV_X1 T404 ( .Y(T404_Y), .A(T14766_Q));
KC_INV_X1 T15691 ( .Y(T15691_Y), .A(T14933_Q));
KC_INV_X1 T15404 ( .Y(T15404_Y), .A(T1886_Y));
KC_INV_X1 T15902 ( .Y(T15902_Y), .A(T3614_Y));
KC_INV_X1 T6770 ( .Y(T6770_Y), .A(T14838_Q));
KC_INV_X1 T6768 ( .Y(T6768_Y), .A(T16079_Q));
KC_INV_X1 T6767 ( .Y(T6767_Y), .A(T16079_Q));
KC_INV_X1 T6765 ( .Y(T6765_Y), .A(T14984_Y));
KC_INV_X1 T6762 ( .Y(T6762_Y), .A(T10369_Y));
KC_INV_X1 T634 ( .Y(T634_Y), .A(T2454_Y));
KC_INV_X1 T633 ( .Y(T633_Y), .A(T2466_Y));
KC_INV_X1 T611 ( .Y(T611_Y), .A(T2478_Y));
KC_INV_X1 T610 ( .Y(T610_Y), .A(T2476_Y));
KC_INV_X1 T609 ( .Y(T609_Y), .A(T4252_Y));
KC_INV_X1 T15682 ( .Y(T15682_Y), .A(T16079_Q));
KC_INV_X1 T15681 ( .Y(T15681_Y), .A(T1535_Y));
KC_INV_X1 T15422 ( .Y(T15422_Y), .A(T16079_Q));
KC_INV_X1 T15419 ( .Y(T15419_Y), .A(T4986_Y));
KC_INV_X1 T16194 ( .Y(T16194_Y), .A(T3070_Y));
KC_INV_X1 T883 ( .Y(T883_Y), .A(T2861_Y));
KC_INV_X1 T882 ( .Y(T882_Y), .A(T5021_Y));
KC_INV_X1 T15447 ( .Y(T15447_Y), .A(T2529_Y));
KC_INV_X1 T15443 ( .Y(T15443_Y), .A(T2526_Q));
KC_INV_X1 T16412 ( .Y(T16412_Y), .A(T12735_Y));
KC_INV_X1 T1141 ( .Y(T1141_Y), .A(T2591_Q));
KC_INV_X1 T1138 ( .Y(T1138_Y), .A(T5322_Y));
KC_INV_X1 T1114 ( .Y(T1114_Y), .A(T14995_Y));
KC_INV_X1 T1103 ( .Y(T1103_Y), .A(T10509_Y));
KC_INV_X1 T1102 ( .Y(T1102_Y), .A(T2567_Y));
KC_INV_X1 T1101 ( .Y(T1101_Y), .A(T15476_Y));
KC_INV_X1 T1097 ( .Y(T1097_Y), .A(T3713_Y));
KC_INV_X1 T15477 ( .Y(T15477_Y), .A(T5869_Co));
KC_INV_X1 T15473 ( .Y(T15473_Y), .A(T3685_Y));
KC_INV_X1 T16411 ( .Y(T16411_Y), .A(T2551_Y));
KC_INV_X1 T1546 ( .Y(T1546_Y), .A(T14367_Q));
KC_INV_X1 T1544 ( .Y(T1544_Y), .A(T14342_Q));
KC_INV_X1 T1524 ( .Y(T1524_Y), .A(T3129_Y));
KC_INV_X1 T1508 ( .Y(T1508_Y), .A(T2627_Q));
KC_INV_X1 T1499 ( .Y(T1499_Y), .A(T2625_Q));
KC_INV_X1 T1482 ( .Y(T1482_Y), .A(T4291_Y));
KC_INV_X1 T15518 ( .Y(T15518_Y), .A(T12091_Y));
KC_INV_X1 T15503 ( .Y(T15503_Y), .A(T4982_Y));
KC_INV_X1 T15502 ( .Y(T15502_Y), .A(T2057_Y));
KC_INV_X1 T15501 ( .Y(T15501_Y), .A(T2604_Y));
KC_INV_X1 T16234 ( .Y(T16234_Y), .A(T14514_Q));
KC_INV_X1 T4898 ( .Y(T4898_Y), .A(T4981_Y));
KC_INV_X1 T4896 ( .Y(T4896_Y), .A(T10184_Y));
KC_INV_X1 T4895 ( .Y(T4895_Y), .A(T2062_Y));
KC_INV_X1 T4886 ( .Y(T4886_Y), .A(T3763_Y));
KC_INV_X1 T4883 ( .Y(T4883_Y), .A(T3166_Y));
KC_INV_X1 T4871 ( .Y(T4871_Y), .A(T3742_Y));
KC_INV_X1 T4867 ( .Y(T4867_Y), .A(T3161_Y));
KC_INV_X1 T4864 ( .Y(T4864_Y), .A(T3761_Y));
KC_INV_X1 T4852 ( .Y(T4852_Y), .A(T3739_Y));
KC_INV_X1 T15535 ( .Y(T15535_Y), .A(T2640_Q));
KC_INV_X1 T15533 ( .Y(T15533_Y), .A(T16079_Q));
KC_INV_X1 T15532 ( .Y(T15532_Y), .A(T10239_Y));
KC_INV_X1 T15552 ( .Y(T15552_Y), .A(T14984_Y));
KC_INV_X1 T16161 ( .Y(T16161_Y), .A(T10274_Y));
KC_INV_X1 T5754 ( .Y(T5754_Y), .A(T5576_Q));
KC_INV_X1 T5751 ( .Y(T5751_Y), .A(T5421_Q));
KC_INV_X1 T5750 ( .Y(T5750_Y), .A(T10273_Y));
KC_INV_X1 T5749 ( .Y(T5749_Y), .A(T2662_Y));
KC_INV_X1 T5741 ( .Y(T5741_Y), .A(T2468_Y));
KC_INV_X1 T5740 ( .Y(T5740_Y), .A(T2483_Y));
KC_INV_X1 T5738 ( .Y(T5738_Y), .A(T2484_Y));
KC_INV_X1 T5724 ( .Y(T5724_Y), .A(T11355_Y));
KC_INV_X1 T5717 ( .Y(T5717_Y), .A(T5424_Q));
KC_INV_X1 T5714 ( .Y(T5714_Y), .A(T2663_Y));
KC_INV_X1 T5710 ( .Y(T5710_Y), .A(T5425_Q));
KC_INV_X1 T15861 ( .Y(T15861_Y), .A(T11321_Y));
KC_INV_X1 T15754 ( .Y(T15754_Y), .A(T10270_Y));
KC_INV_X1 T15753 ( .Y(T15753_Y), .A(T11009_Y));
KC_INV_X1 T5786 ( .Y(T5786_Y), .A(T11362_Y));
KC_INV_X1 T5784 ( .Y(T5784_Y), .A(T11343_Y));
KC_INV_X1 T5776 ( .Y(T5776_Y), .A(T11963_Y));
KC_INV_X1 T5775 ( .Y(T5775_Y), .A(T11341_Y));
KC_INV_X1 T5773 ( .Y(T5773_Y), .A(T14535_Q));
KC_INV_X1 T5766 ( .Y(T5766_Y), .A(T14954_Q));
KC_INV_X1 T5758 ( .Y(T5758_Y), .A(T14528_Q));
KC_INV_X1 T15700 ( .Y(T15700_Y), .A(T15231_Y));
KC_INV_X1 T15696 ( .Y(T15696_Y), .A(T10281_Y));
KC_INV_X1 T5791 ( .Y(T5791_Y), .A(T10945_Y));
KC_INV_X1 T15895 ( .Y(T15895_Y), .A(T15803_Q));
KC_INV_X1 T5845 ( .Y(T5845_Y), .A(T3860_Y));
KC_INV_X1 T5819 ( .Y(T5819_Y), .A(T8198_Y));
KC_INV_X1 T5813 ( .Y(T5813_Y), .A(T15880_Q));
KC_INV_X1 T5812 ( .Y(T5812_Y), .A(T15879_Q));
KC_INV_X1 T15928 ( .Y(T15928_Y), .A(T10643_Y));
KC_INV_X1 T15912 ( .Y(T15912_Y), .A(T5380_Q));
KC_INV_X1 T5875 ( .Y(T5875_Y), .A(T12248_Y));
KC_INV_X1 T15566 ( .Y(T15566_Y), .A(T2752_Q));
KC_INV_X1 T5941 ( .Y(T5941_Y), .A(T3284_Y));
KC_INV_X1 T5925 ( .Y(T5925_Y), .A(T13128_Q));
KC_INV_X1 T5924 ( .Y(T5924_Y), .A(T4177_Y));
KC_INV_X1 T5896 ( .Y(T5896_Y), .A(T11604_Y));
KC_INV_X1 T5877 ( .Y(T5877_Y), .A(T2747_Y));
KC_INV_X1 T15582 ( .Y(T15582_Y), .A(T2754_Y));
KC_INV_X1 T15579 ( .Y(T15579_Y), .A(T10641_Y));
KC_INV_X1 T16003 ( .Y(T16003_Y), .A(T8338_Y));
KC_INV_X1 T15982 ( .Y(T15982_Y), .A(T11581_Y));
KC_INV_X1 T5978 ( .Y(T5978_Y), .A(T12460_Y));
KC_INV_X1 T15597 ( .Y(T15597_Y), .A(T2778_Y));
KC_INV_X1 T15596 ( .Y(T15596_Y), .A(T8492_Y));
KC_INV_X1 T16024 ( .Y(T16024_Y), .A(T11970_Y));
KC_INV_X1 T16015 ( .Y(T16015_Y), .A(T14563_Q));
KC_INV_X1 T6013 ( .Y(T6013_Y), .A(T8286_Y));
KC_INV_X1 T6011 ( .Y(T6011_Y), .A(T2723_Y));
KC_INV_X1 T6007 ( .Y(T6007_Y), .A(T5058_Y));
KC_INV_X1 T5999 ( .Y(T5999_Y), .A(T2756_Y));
KC_INV_X1 T15600 ( .Y(T15600_Y), .A(T3516_Y));
KC_INV_X1 T16101 ( .Y(T16101_Y), .A(T4748_Y));
KC_INV_X1 T16100 ( .Y(T16100_Y), .A(T2800_Y));
KC_INV_X1 T16099 ( .Y(T16099_Y), .A(T8261_Y));
KC_INV_X1 T16056 ( .Y(T16056_Y), .A(T16055_Y));
KC_INV_X1 T16055 ( .Y(T16055_Y), .A(T15038_Y));
KC_INV_X1 T6088 ( .Y(T6088_Y), .A(T5539_Y));
KC_INV_X1 T6085 ( .Y(T6085_Y), .A(T3379_Y));
KC_INV_X1 T6072 ( .Y(T6072_Y), .A(T16056_Y));
KC_INV_X1 T6070 ( .Y(T6070_Y), .A(T2854_Y));
KC_INV_X1 T6054 ( .Y(T6054_Y), .A(T2833_Q));
KC_INV_X1 T6039 ( .Y(T6039_Y), .A(T15234_Y));
KC_INV_X1 T15615 ( .Y(T15615_Y), .A(T11647_Y));
KC_INV_X1 T6183 ( .Y(T6183_Y), .A(T2874_Q));
KC_INV_X1 T6182 ( .Y(T6182_Y), .A(T3436_Y));
KC_INV_X1 T6181 ( .Y(T6181_Y), .A(T2876_Y));
KC_INV_X1 T6180 ( .Y(T6180_Y), .A(T11831_Y));
KC_INV_X1 T6161 ( .Y(T6161_Y), .A(T11743_Y));
KC_INV_X1 T6160 ( .Y(T6160_Y), .A(T11809_Y));
KC_INV_X1 T6159 ( .Y(T6159_Y), .A(T11739_Y));
KC_INV_X1 T6145 ( .Y(T6145_Y), .A(T12104_Y));
KC_INV_X1 T6144 ( .Y(T6144_Y), .A(T2870_Y));
KC_INV_X1 T6140 ( .Y(T6140_Y), .A(T12039_Y));
KC_INV_X1 T6124 ( .Y(T6124_Y), .A(T6511_Y));
KC_INV_X1 T6123 ( .Y(T6123_Y), .A(T10986_Y));
KC_INV_X1 T6100 ( .Y(T6100_Y), .A(T2882_Y));
KC_INV_X1 T15624 ( .Y(T15624_Y), .A(T2871_Y));
KC_INV_X1 T15622 ( .Y(T15622_Y), .A(T2860_Y));
KC_INV_X1 T15953 ( .Y(T15953_Y), .A(T2896_Y));
KC_INV_X1 T16132 ( .Y(T16132_Y), .A(T10555_Y));
KC_INV_X1 T6583 ( .Y(T6583_Y), .A(T10553_Y));
KC_INV_X1 T6582 ( .Y(T6582_Y), .A(T11741_Y));
KC_INV_X1 T6580 ( .Y(T6580_Y), .A(T6581_Y));
KC_INV_X1 T6578 ( .Y(T6578_Y), .A(T11742_Y));
KC_INV_X1 T6576 ( .Y(T6576_Y), .A(T5515_Y));
KC_INV_X1 T6573 ( .Y(T6573_Y), .A(T2887_Y));
KC_INV_X1 T6572 ( .Y(T6572_Y), .A(T10558_Y));
KC_INV_X1 T6559 ( .Y(T6559_Y), .A(T15255_Y));
KC_INV_X1 T6239 ( .Y(T6239_Y), .A(T2909_Y));
KC_INV_X1 T6237 ( .Y(T6237_Y), .A(T10985_Y));
KC_INV_X1 T6225 ( .Y(T6225_Y), .A(T12107_Y));
KC_INV_X1 T6224 ( .Y(T6224_Y), .A(T2900_Y));
KC_INV_X1 T6223 ( .Y(T6223_Y), .A(T10988_Y));
KC_INV_X1 T6222 ( .Y(T6222_Y), .A(T12106_Y));
KC_INV_X1 T6221 ( .Y(T6221_Y), .A(T2911_Y));
KC_INV_X1 T6214 ( .Y(T6214_Y), .A(T12064_Y));
KC_INV_X1 T6196 ( .Y(T6196_Y), .A(T3489_Y));
KC_INV_X1 T6195 ( .Y(T6195_Y), .A(T2952_Q));
KC_INV_X1 T6192 ( .Y(T6192_Y), .A(T11037_Y));
KC_INV_X1 T6190 ( .Y(T6190_Y), .A(T11744_Y));
KC_INV_X1 T290 ( .Y(T290_Y), .A(T4054_Y));
KC_INV_X1 T15632 ( .Y(T15632_Y), .A(T2926_Y));
KC_INV_X1 T15627 ( .Y(T15627_Y), .A(T2325_Y));
KC_INV_X1 T6539 ( .Y(T6539_Y), .A(T6538_Y));
KC_INV_X1 T6538 ( .Y(T6538_Y), .A(T12067_Y));
KC_INV_X1 T6537 ( .Y(T6537_Y), .A(T2959_Y));
KC_INV_X1 T6532 ( .Y(T6532_Y), .A(T11836_Y));
KC_INV_X1 T6531 ( .Y(T6531_Y), .A(T2941_Y));
KC_INV_X1 T6530 ( .Y(T6530_Y), .A(T4055_Y));
KC_INV_X1 T6509 ( .Y(T6509_Y), .A(T5536_Q));
KC_INV_X1 T6506 ( .Y(T6506_Y), .A(T11002_Y));
KC_INV_X1 T6488 ( .Y(T6488_Y), .A(T2943_Q));
KC_INV_X1 T15643 ( .Y(T15643_Y), .A(T5540_Y));
KC_INV_X1 T374 ( .Y(T374_Y), .A(T3001_Y));
KC_INV_X1 T15679 ( .Y(T15679_Y), .A(T2981_Y));
KC_INV_X1 T15383 ( .Y(T15383_Y), .A(T3565_Y));
KC_INV_X1 T6761 ( .Y(T6761_Y), .A(T14931_Q));
KC_INV_X1 T483 ( .Y(T483_Y), .A(T13781_Q));
KC_INV_X1 T478 ( .Y(T478_Y), .A(T2991_Y));
KC_INV_X1 T475 ( .Y(T475_Y), .A(T3014_Y));
KC_INV_X1 T431 ( .Y(T431_Y), .A(T2962_Y));
KC_INV_X1 T424 ( .Y(T424_Y), .A(T3587_Y));
KC_INV_X1 T423 ( .Y(T423_Y), .A(T3549_Y));
KC_INV_X1 T15403 ( .Y(T15403_Y), .A(T13767_Q));
KC_INV_X1 T15397 ( .Y(T15397_Y), .A(T3536_Y));
KC_INV_X1 T632 ( .Y(T632_Y), .A(T3037_Y));
KC_INV_X1 T602 ( .Y(T602_Y), .A(T3051_Y));
KC_INV_X1 T15683 ( .Y(T15683_Y), .A(T2467_Y));
KC_INV_X1 T15424 ( .Y(T15424_Y), .A(T5268_Y));
KC_INV_X1 T15420 ( .Y(T15420_Y), .A(T5270_Y));
KC_INV_X1 T884 ( .Y(T884_Y), .A(T3669_Y));
KC_INV_X1 T881 ( .Y(T881_Y), .A(T2525_Q));
KC_INV_X1 T880 ( .Y(T880_Y), .A(T3679_Y));
KC_INV_X1 T875 ( .Y(T875_Y), .A(T10239_Y));
KC_INV_X1 T874 ( .Y(T874_Y), .A(T3627_Y));
KC_INV_X1 T872 ( .Y(T872_Y), .A(T14082_Q));
KC_INV_X1 T871 ( .Y(T871_Y), .A(T4231_Y));
KC_INV_X1 T870 ( .Y(T870_Y), .A(T4250_Y));
KC_INV_X1 T866 ( .Y(T866_Y), .A(T5083_Y));
KC_INV_X1 T864 ( .Y(T864_Y), .A(T5825_S));
KC_INV_X1 T859 ( .Y(T859_Y), .A(T14032_Q));
KC_INV_X1 T15442 ( .Y(T15442_Y), .A(T2674_Y));
KC_INV_X1 T1136 ( .Y(T1136_Y), .A(T3137_Y));
KC_INV_X1 T1132 ( .Y(T1132_Y), .A(T2065_Y));
KC_INV_X1 T1109 ( .Y(T1109_Y), .A(T3082_Y));
KC_INV_X1 T1108 ( .Y(T1108_Y), .A(T12089_Y));
KC_INV_X1 T5748 ( .Y(T5748_Y), .A(T10241_Y));
KC_INV_X1 T5747 ( .Y(T5747_Y), .A(T10242_Y));
KC_INV_X1 T5736 ( .Y(T5736_Y), .A(T2516_Y));
KC_INV_X1 T5734 ( .Y(T5734_Y), .A(T2514_Y));
KC_INV_X1 T5729 ( .Y(T5729_Y), .A(T4987_Y));
KC_INV_X1 T5706 ( .Y(T5706_Y), .A(T2512_Y));
KC_INV_X1 T5704 ( .Y(T5704_Y), .A(T2509_Y));
KC_INV_X1 T5544 ( .Y(T5544_Y), .A(T2455_Y));
KC_INV_X1 T5405 ( .Y(T5405_Y), .A(T2461_Y));
KC_INV_X1 T15550 ( .Y(T15550_Y), .A(T2511_Y));
KC_INV_X1 T15549 ( .Y(T15549_Y), .A(T2515_Y));
KC_INV_X1 T15548 ( .Y(T15548_Y), .A(T2470_Y));
KC_INV_X1 T15546 ( .Y(T15546_Y), .A(T2513_Y));
KC_INV_X1 T15864 ( .Y(T15864_Y), .A(T14956_Q));
KC_INV_X1 T15832 ( .Y(T15832_Y), .A(T5425_Q));
KC_INV_X1 T15826 ( .Y(T15826_Y), .A(T5750_Y));
KC_INV_X1 T15821 ( .Y(T15821_Y), .A(T14529_Q));
KC_INV_X1 T15819 ( .Y(T15819_Y), .A(T3184_Y));
KC_INV_X1 T5783 ( .Y(T5783_Y), .A(T11394_Y));
KC_INV_X1 T5774 ( .Y(T5774_Y), .A(T16160_Y));
KC_INV_X1 T5765 ( .Y(T5765_Y), .A(T13069_Y));
KC_INV_X1 T5764 ( .Y(T5764_Y), .A(T14534_Q));
KC_INV_X1 T15694 ( .Y(T15694_Y), .A(T11335_Y));
KC_INV_X1 T15559 ( .Y(T15559_Y), .A(T5040_Y));
KC_INV_X1 T15929 ( .Y(T15929_Y), .A(T10642_Y));
KC_INV_X1 T15911 ( .Y(T15911_Y), .A(T8199_Y));
KC_INV_X1 T5871 ( .Y(T5871_Y), .A(T8223_Y));
KC_INV_X1 T5860 ( .Y(T5860_Y), .A(T5022_Y));
KC_INV_X1 T15960 ( .Y(T15960_Y), .A(T2777_Y));
KC_INV_X1 T5890 ( .Y(T5890_Y), .A(T13139_Y));
KC_INV_X1 T5942 ( .Y(T5942_Y), .A(T10630_Y));
KC_INV_X1 T5940 ( .Y(T5940_Y), .A(T11457_Y));
KC_INV_X1 T5939 ( .Y(T5939_Y), .A(T13104_Q));
KC_INV_X1 T5923 ( .Y(T5923_Y), .A(T3268_Y));
KC_INV_X1 T5922 ( .Y(T5922_Y), .A(T15981_Y));
KC_INV_X1 T5921 ( .Y(T5921_Y), .A(T5922_Y));
KC_INV_X1 T5894 ( .Y(T5894_Y), .A(T3295_Y));
KC_INV_X1 T5893 ( .Y(T5893_Y), .A(T11486_Y));
KC_INV_X1 T16002 ( .Y(T16002_Y), .A(T15855_Y));
KC_INV_X1 T16001 ( .Y(T16001_Y), .A(T3991_Y));
KC_INV_X1 T16000 ( .Y(T16000_Y), .A(T12215_Y));
KC_INV_X1 T15980 ( .Y(T15980_Y), .A(T3951_Y));
KC_INV_X1 T15978 ( .Y(T15978_Y), .A(T13139_Y));
KC_INV_X1 T15977 ( .Y(T15977_Y), .A(T12461_Y));
KC_INV_X1 T15976 ( .Y(T15976_Y), .A(T16083_Y));
KC_INV_X1 T5965 ( .Y(T5965_Y), .A(T12817_Y));
KC_INV_X1 T5964 ( .Y(T5964_Y), .A(T6278_Y));
KC_INV_X1 T15591 ( .Y(T15591_Y), .A(T10637_Y));
KC_INV_X1 T16014 ( .Y(T16014_Y), .A(T15960_Y));
KC_INV_X1 T6024 ( .Y(T6024_Y), .A(T11558_Y));
KC_INV_X1 T6006 ( .Y(T6006_Y), .A(T16302_Y));
KC_INV_X1 T5996 ( .Y(T5996_Y), .A(T2806_Y));
KC_INV_X1 T15607 ( .Y(T15607_Y), .A(T16022_Y));
KC_INV_X1 T15598 ( .Y(T15598_Y), .A(T12001_Y));
KC_INV_X1 T16105 ( .Y(T16105_Y), .A(T12043_Y));
KC_INV_X1 T16103 ( .Y(T16103_Y), .A(T10979_Y));
KC_INV_X1 T16102 ( .Y(T16102_Y), .A(T12322_Y));
KC_INV_X1 T16043 ( .Y(T16043_Y), .A(T3399_Y));
KC_INV_X1 T16036 ( .Y(T16036_Y), .A(T11996_Y));
KC_INV_X1 T6086 ( .Y(T6086_Y), .A(T12876_Y));
KC_INV_X1 T6084 ( .Y(T6084_Y), .A(T3362_Y));
KC_INV_X1 T6082 ( .Y(T6082_Y), .A(T4021_Y));
KC_INV_X1 T6081 ( .Y(T6081_Y), .A(T11677_Y));
KC_INV_X1 T6080 ( .Y(T6080_Y), .A(T10584_Y));
KC_INV_X1 T6069 ( .Y(T6069_Y), .A(T11769_Y));
KC_INV_X1 T6067 ( .Y(T6067_Y), .A(T12263_Y));
KC_INV_X1 T6065 ( .Y(T6065_Y), .A(T2841_Q));
KC_INV_X1 T6064 ( .Y(T6064_Y), .A(T3412_Q));
KC_INV_X1 T6052 ( .Y(T6052_Y), .A(T12829_Y));
KC_INV_X1 T6051 ( .Y(T6051_Y), .A(T10590_Y));
KC_INV_X1 T6050 ( .Y(T6050_Y), .A(T3396_Y));
KC_INV_X1 T6047 ( .Y(T6047_Y), .A(T3355_Y));
KC_INV_X1 T6046 ( .Y(T6046_Y), .A(T11642_Y));
KC_INV_X1 T6045 ( .Y(T6045_Y), .A(T10962_Y));
KC_INV_X1 T6036 ( .Y(T6036_Y), .A(T12249_Y));
KC_INV_X1 T15613 ( .Y(T15613_Y), .A(T11664_Y));
KC_INV_X1 T15612 ( .Y(T15612_Y), .A(T4031_Y));
KC_INV_X1 T8401 ( .Y(T8401_Y), .A(T3318_Y));
KC_INV_X1 T6179 ( .Y(T6179_Y), .A(T3530_Y));
KC_INV_X1 T6177 ( .Y(T6177_Y), .A(T12877_Y));
KC_INV_X1 T6158 ( .Y(T6158_Y), .A(T3394_Y));
KC_INV_X1 T6141 ( .Y(T6141_Y), .A(T3445_Y));
KC_INV_X1 T6139 ( .Y(T6139_Y), .A(T5046_Y));
KC_INV_X1 T6138 ( .Y(T6138_Y), .A(T3429_Y));
KC_INV_X1 T6120 ( .Y(T6120_Y), .A(T16148_Y));
KC_INV_X1 T6119 ( .Y(T6119_Y), .A(T12317_Y));
KC_INV_X1 T6098 ( .Y(T6098_Y), .A(T3490_Y));
KC_INV_X1 T6096 ( .Y(T6096_Y), .A(T3515_Y));
KC_INV_X1 T15616 ( .Y(T15616_Y), .A(T3443_Y));
KC_INV_X1 T16139 ( .Y(T16139_Y), .A(T6820_Y));
KC_INV_X1 T6585 ( .Y(T6585_Y), .A(T5522_Y));
KC_INV_X1 T6561 ( .Y(T6561_Y), .A(T2865_Y));
KC_INV_X1 T6236 ( .Y(T6236_Y), .A(T2906_Y));
KC_INV_X1 T6215 ( .Y(T6215_Y), .A(T10571_Y));
KC_INV_X1 T6213 ( .Y(T6213_Y), .A(T11765_Y));
KC_INV_X1 T6211 ( .Y(T6211_Y), .A(T5519_Y));
KC_INV_X1 T6209 ( .Y(T6209_Y), .A(T3528_Q));
KC_INV_X1 T6193 ( .Y(T6193_Y), .A(T3514_Y));
KC_INV_X1 T15711 ( .Y(T15711_Y), .A(T3526_Y));
KC_INV_X1 T15637 ( .Y(T15637_Y), .A(T3468_Y));
KC_INV_X1 T15636 ( .Y(T15636_Y), .A(T11746_Y));
KC_INV_X1 T6529 ( .Y(T6529_Y), .A(T4096_Y));
KC_INV_X1 T6516 ( .Y(T6516_Y), .A(T6469_Y));
KC_INV_X1 T6514 ( .Y(T6514_Y), .A(T3525_Q));
KC_INV_X1 T6512 ( .Y(T6512_Y), .A(T3521_Q));
KC_INV_X1 T6510 ( .Y(T6510_Y), .A(T8150_Y));
KC_INV_X1 T6490 ( .Y(T6490_Y), .A(T3519_Q));
KC_INV_X1 T6489 ( .Y(T6489_Y), .A(T3520_Q));
KC_INV_X1 T15641 ( .Y(T15641_Y), .A(T6614_S));
KC_INV_X1 T15640 ( .Y(T15640_Y), .A(T4164_Q));
KC_INV_X1 T15402 ( .Y(T15402_Y), .A(T3608_Y));
KC_INV_X1 T6846 ( .Y(T6846_Y), .A(T9733_Y));
KC_INV_X1 T6839 ( .Y(T6839_Y), .A(T3653_Y));
KC_INV_X1 T6802 ( .Y(T6802_Y), .A(T3650_Y));
KC_INV_X1 T622 ( .Y(T622_Y), .A(T5134_Y));
KC_INV_X1 T607 ( .Y(T607_Y), .A(T3621_Y));
KC_INV_X1 T16230 ( .Y(T16230_Y), .A(T14878_Q));
KC_INV_X1 T879 ( .Y(T879_Y), .A(T3666_Y));
KC_INV_X1 T857 ( .Y(T857_Y), .A(T3657_Y));
KC_INV_X1 T856 ( .Y(T856_Y), .A(T3667_Y));
KC_INV_X1 T16403 ( .Y(T16403_Y), .A(T3712_Y));
KC_INV_X1 T16402 ( .Y(T16402_Y), .A(T3069_Y));
KC_INV_X1 T5563 ( .Y(T5563_Y), .A(T2485_Y));
KC_INV_X1 T15870 ( .Y(T15870_Y), .A(T3795_Y));
KC_INV_X1 T15869 ( .Y(T15869_Y), .A(T11969_Y));
KC_INV_X1 T15867 ( .Y(T15867_Y), .A(T11985_Y));
KC_INV_X1 T15845 ( .Y(T15845_Y), .A(T3794_Y));
KC_INV_X1 T5781 ( .Y(T5781_Y), .A(T11389_Y));
KC_INV_X1 T5780 ( .Y(T5780_Y), .A(T11379_Y));
KC_INV_X1 T5772 ( .Y(T5772_Y), .A(T11336_Y));
KC_INV_X1 T5771 ( .Y(T5771_Y), .A(T3842_Y));
KC_INV_X1 T5770 ( .Y(T5770_Y), .A(T11353_Y));
KC_INV_X1 T5763 ( .Y(T5763_Y), .A(T5101_Y));
KC_INV_X1 T5756 ( .Y(T5756_Y), .A(T11983_Y));
KC_INV_X1 T15558 ( .Y(T15558_Y), .A(T3802_Y));
KC_INV_X1 T15896 ( .Y(T15896_Y), .A(T11419_Y));
KC_INV_X1 T15877 ( .Y(T15877_Y), .A(T3849_Y));
KC_INV_X1 T5843 ( .Y(T5843_Y), .A(T15186_Y));
KC_INV_X1 T5842 ( .Y(T5842_Y), .A(T11367_Y));
KC_INV_X1 T5840 ( .Y(T5840_Y), .A(T11426_Y));
KC_INV_X1 T5838 ( .Y(T5838_Y), .A(T15908_Y));
KC_INV_X1 T5837 ( .Y(T5837_Y), .A(T8188_Y));
KC_INV_X1 T5830 ( .Y(T5830_Y), .A(T3826_Y));
KC_INV_X1 T5827 ( .Y(T5827_Y), .A(T4438_Y));
KC_INV_X1 T5826 ( .Y(T5826_Y), .A(T3827_Y));
KC_INV_X1 T5816 ( .Y(T5816_Y), .A(T11365_Y));
KC_INV_X1 T5806 ( .Y(T5806_Y), .A(T11370_Y));
KC_INV_X1 T5803 ( .Y(T5803_Y), .A(T11427_Y));
KC_INV_X1 T5802 ( .Y(T5802_Y), .A(T11410_Y));
KC_INV_X1 T5801 ( .Y(T5801_Y), .A(T11428_Y));
KC_INV_X1 T5800 ( .Y(T5800_Y), .A(T15897_Y));
KC_INV_X1 T5790 ( .Y(T5790_Y), .A(T6068_Y));
KC_INV_X1 T5789 ( .Y(T5789_Y), .A(T4487_Q));
KC_INV_X1 T5788 ( .Y(T5788_Y), .A(T4465_Q));
KC_INV_X1 T15562 ( .Y(T15562_Y), .A(T5446_Y));
KC_INV_X1 T15940 ( .Y(T15940_Y), .A(T6797_Co));
KC_INV_X1 T15939 ( .Y(T15939_Y), .A(T3868_Y));
KC_INV_X1 T15919 ( .Y(T15919_Y), .A(T16152_Y));
KC_INV_X1 T15918 ( .Y(T15918_Y), .A(T10641_Y));
KC_INV_X1 T15917 ( .Y(T15917_Y), .A(T2787_Y));
KC_INV_X1 T5874 ( .Y(T5874_Y), .A(T3889_Q));
KC_INV_X1 T5870 ( .Y(T5870_Y), .A(T3890_Q));
KC_INV_X1 T5868 ( .Y(T5868_Y), .A(T4493_Q));
KC_INV_X1 T5859 ( .Y(T5859_Y), .A(T2077_Y));
KC_INV_X1 T5858 ( .Y(T5858_Y), .A(T3878_Q));
KC_INV_X1 T15571 ( .Y(T15571_Y), .A(T3873_Q));
KC_INV_X1 T15945 ( .Y(T15945_Y), .A(T11587_Y));
KC_INV_X1 T5937 ( .Y(T5937_Y), .A(T3904_Y));
KC_INV_X1 T5919 ( .Y(T5919_Y), .A(T15961_Y));
KC_INV_X1 T5907 ( .Y(T5907_Y), .A(T3936_Q));
KC_INV_X1 T5905 ( .Y(T5905_Y), .A(T5459_Y));
KC_INV_X1 T5892 ( .Y(T5892_Y), .A(T3935_Q));
KC_INV_X1 T15581 ( .Y(T15581_Y), .A(T3887_Y));
KC_INV_X1 T15580 ( .Y(T15580_Y), .A(T6219_Y));
KC_INV_X1 T15578 ( .Y(T15578_Y), .A(T8237_Y));
KC_INV_X1 T15576 ( .Y(T15576_Y), .A(T4473_Y));
KC_INV_X1 T15994 ( .Y(T15994_Y), .A(T16453_Q));
KC_INV_X1 T15985 ( .Y(T15985_Y), .A(T3883_Q));
KC_INV_X1 T5989 ( .Y(T5989_Y), .A(T11534_Y));
KC_INV_X1 T5986 ( .Y(T5986_Y), .A(T11555_Y));
KC_INV_X1 T5985 ( .Y(T5985_Y), .A(T4549_Y));
KC_INV_X1 T5981 ( .Y(T5981_Y), .A(T10937_Y));
KC_INV_X1 T5973 ( .Y(T5973_Y), .A(T3965_Q));
KC_INV_X1 T5972 ( .Y(T5972_Y), .A(T3970_Q));
KC_INV_X1 T5963 ( .Y(T5963_Y), .A(T3949_Y));
KC_INV_X1 T5958 ( .Y(T5958_Y), .A(T10944_Y));
KC_INV_X1 T5957 ( .Y(T5957_Y), .A(T3975_Y));
KC_INV_X1 T5956 ( .Y(T5956_Y), .A(T16167_Y));
KC_INV_X1 T15589 ( .Y(T15589_Y), .A(T3968_Q));
KC_INV_X1 T15588 ( .Y(T15588_Y), .A(T3947_Y));
KC_INV_X1 T15587 ( .Y(T15587_Y), .A(T3964_Q));
KC_INV_X1 T6025 ( .Y(T6025_Y), .A(T5479_Q));
KC_INV_X1 T6023 ( .Y(T6023_Y), .A(T5972_Y));
KC_INV_X1 T6020 ( .Y(T6020_Y), .A(T6352_Y));
KC_INV_X1 T5995 ( .Y(T5995_Y), .A(T12239_Y));
KC_INV_X1 T5992 ( .Y(T5992_Y), .A(T12957_Y));
KC_INV_X1 T15610 ( .Y(T15610_Y), .A(T8277_Y));
KC_INV_X1 T15606 ( .Y(T15606_Y), .A(T16457_Q));
KC_INV_X1 T15601 ( .Y(T15601_Y), .A(T3937_Q));
KC_INV_X1 T16108 ( .Y(T16108_Y), .A(T4046_Y));
KC_INV_X1 T6044 ( .Y(T6044_Y), .A(T15760_Q));
KC_INV_X1 T16031 ( .Y(T16031_Y), .A(T11671_Y));
KC_INV_X1 T16030 ( .Y(T16030_Y), .A(T5114_Y));
KC_INV_X1 T16029 ( .Y(T16029_Y), .A(T1820_Q));
KC_INV_X1 T16028 ( .Y(T16028_Y), .A(T5114_Y));
KC_INV_X1 T6083 ( .Y(T6083_Y), .A(T11641_Y));
KC_INV_X1 T6079 ( .Y(T6079_Y), .A(T4176_Q));
KC_INV_X1 T6078 ( .Y(T6078_Y), .A(T4589_Y));
KC_INV_X1 T6077 ( .Y(T6077_Y), .A(T5466_Y));
KC_INV_X1 T6076 ( .Y(T6076_Y), .A(T5498_Q));
KC_INV_X1 T6062 ( .Y(T6062_Y), .A(T4032_Y));
KC_INV_X1 T6060 ( .Y(T6060_Y), .A(T4051_Q));
KC_INV_X1 T6048 ( .Y(T6048_Y), .A(T5525_Q));
KC_INV_X1 T6043 ( .Y(T6043_Y), .A(T4179_Q));
KC_INV_X1 T6034 ( .Y(T6034_Y), .A(T5530_Q));
KC_INV_X1 T6033 ( .Y(T6033_Y), .A(T6841_S));
KC_INV_X1 T8382 ( .Y(T8382_Y), .A(T16133_Y));
KC_INV_X1 T16124 ( .Y(T16124_Y), .A(T8386_Y));
KC_INV_X1 T6176 ( .Y(T6176_Y), .A(T8503_Y));
KC_INV_X1 T6175 ( .Y(T6175_Y), .A(T4147_Q));
KC_INV_X1 T6174 ( .Y(T6174_Y), .A(T12279_Y));
KC_INV_X1 T6170 ( .Y(T6170_Y), .A(T5568_Q));
KC_INV_X1 T6157 ( .Y(T6157_Y), .A(T5135_Y));
KC_INV_X1 T6156 ( .Y(T6156_Y), .A(T4178_Q));
KC_INV_X1 T6155 ( .Y(T6155_Y), .A(T10581_Y));
KC_INV_X1 T6151 ( .Y(T6151_Y), .A(T5504_Y));
KC_INV_X1 T6137 ( .Y(T6137_Y), .A(T5510_Y));
KC_INV_X1 T6135 ( .Y(T6135_Y), .A(T4080_Y));
KC_INV_X1 T6134 ( .Y(T6134_Y), .A(T4081_Y));
KC_INV_X1 T6112 ( .Y(T6112_Y), .A(T10882_Y));
KC_INV_X1 T6111 ( .Y(T6111_Y), .A(T11658_Y));
KC_INV_X1 T6107 ( .Y(T6107_Y), .A(T10583_Y));
KC_INV_X1 T6106 ( .Y(T6106_Y), .A(T10617_Y));
KC_INV_X1 T6105 ( .Y(T6105_Y), .A(T10563_Y));
KC_INV_X1 T6094 ( .Y(T6094_Y), .A(T4083_Y));
KC_INV_X1 T15620 ( .Y(T15620_Y), .A(T4049_Y));
KC_INV_X1 T15619 ( .Y(T15619_Y), .A(T11715_Y));
KC_INV_X1 T16143 ( .Y(T16143_Y), .A(T4163_Q));
KC_INV_X1 T16142 ( .Y(T16142_Y), .A(T4085_Y));
KC_INV_X1 T6587 ( .Y(T6587_Y), .A(T5528_Q));
KC_INV_X1 T6586 ( .Y(T6586_Y), .A(T3427_Y));
KC_INV_X1 T6547 ( .Y(T6547_Y), .A(T2865_Y));
KC_INV_X1 T6210 ( .Y(T6210_Y), .A(T11796_Y));
KC_INV_X1 T6207 ( .Y(T6207_Y), .A(T5532_Q));
KC_INV_X1 T6205 ( .Y(T6205_Y), .A(T6208_Y));
KC_INV_X1 T6188 ( .Y(T6188_Y), .A(T4540_Y));
KC_INV_X1 T15631 ( .Y(T15631_Y), .A(T3481_Y));
KC_INV_X1 T6527 ( .Y(T6527_Y), .A(T4171_Q));
KC_INV_X1 T6524 ( .Y(T6524_Y), .A(T4169_Q));
KC_INV_X1 T6517 ( .Y(T6517_Y), .A(T4168_Q));
KC_INV_X1 T6438 ( .Y(T6438_Y), .A(T2964_Y));
KC_INV_X1 T15365 ( .Y(T15365_Y), .A(T15441_Y));
KC_INV_X1 T15441 ( .Y(T15441_Y), .A(T3073_Y));
KC_INV_X1 T16157 ( .Y(T16157_Y), .A(T14468_Q));
KC_INV_X1 T5746 ( .Y(T5746_Y), .A(T3793_Y));
KC_INV_X1 T15554 ( .Y(T15554_Y), .A(T16213_Y));
KC_INV_X1 T15553 ( .Y(T15553_Y), .A(T12950_Y));
KC_INV_X1 T15872 ( .Y(T15872_Y), .A(T11371_Y));
KC_INV_X1 T15871 ( .Y(T15871_Y), .A(T4383_Y));
KC_INV_X1 T15837 ( .Y(T15837_Y), .A(T4397_Y));
KC_INV_X1 T5778 ( .Y(T5778_Y), .A(T11378_Y));
KC_INV_X1 T5777 ( .Y(T5777_Y), .A(T4403_Y));
KC_INV_X1 T5767 ( .Y(T5767_Y), .A(T4394_Y));
KC_INV_X1 T5762 ( .Y(T5762_Y), .A(T4402_Y));
KC_INV_X1 T5761 ( .Y(T5761_Y), .A(T4401_Y));
KC_INV_X1 T5760 ( .Y(T5760_Y), .A(T14942_Q));
KC_INV_X1 T15557 ( .Y(T15557_Y), .A(T14523_Q));
KC_INV_X1 T15555 ( .Y(T15555_Y), .A(T4394_Y));
KC_INV_X1 T5835 ( .Y(T5835_Y), .A(T4464_Y));
KC_INV_X1 T5824 ( .Y(T5824_Y), .A(T11408_Y));
KC_INV_X1 T5823 ( .Y(T5823_Y), .A(T4439_Y));
KC_INV_X1 T5822 ( .Y(T5822_Y), .A(T4432_Y));
KC_INV_X1 T5821 ( .Y(T5821_Y), .A(T4445_Y));
KC_INV_X1 T5815 ( .Y(T5815_Y), .A(T4457_Y));
KC_INV_X1 T5799 ( .Y(T5799_Y), .A(T13085_Y));
KC_INV_X1 T5798 ( .Y(T5798_Y), .A(T3850_Y));
KC_INV_X1 T5787 ( .Y(T5787_Y), .A(T4463_Y));
KC_INV_X1 T15936 ( .Y(T15936_Y), .A(T10628_Y));
KC_INV_X1 T15935 ( .Y(T15935_Y), .A(T11520_Y));
KC_INV_X1 T5873 ( .Y(T5873_Y), .A(T4467_Y));
KC_INV_X1 T5867 ( .Y(T5867_Y), .A(T3258_Q));
KC_INV_X1 T5862 ( .Y(T5862_Y), .A(T4497_Y));
KC_INV_X1 T5857 ( .Y(T5857_Y), .A(T3222_Y));
KC_INV_X1 T5854 ( .Y(T5854_Y), .A(T14549_Q));
KC_INV_X1 T5853 ( .Y(T5853_Y), .A(T14548_Q));
KC_INV_X1 T5851 ( .Y(T5851_Y), .A(T8444_Y));
KC_INV_X1 T5846 ( .Y(T5846_Y), .A(T6127_Y));
KC_INV_X1 T15697 ( .Y(T15697_Y), .A(T14550_Q));
KC_INV_X1 T15572 ( .Y(T15572_Y), .A(T4496_Y));
KC_INV_X1 T15570 ( .Y(T15570_Y), .A(T4492_Q));
KC_INV_X1 T15569 ( .Y(T15569_Y), .A(T4484_Q));
KC_INV_X1 T8252 ( .Y(T8252_Y), .A(T12199_Y));
KC_INV_X1 T5934 ( .Y(T5934_Y), .A(T12197_Y));
KC_INV_X1 T5932 ( .Y(T5932_Y), .A(T4530_Y));
KC_INV_X1 T5930 ( .Y(T5930_Y), .A(T12182_Y));
KC_INV_X1 T5929 ( .Y(T5929_Y), .A(T4535_Y));
KC_INV_X1 T5917 ( .Y(T5917_Y), .A(T4527_Q));
KC_INV_X1 T5914 ( .Y(T5914_Y), .A(T4474_Y));
KC_INV_X1 T5889 ( .Y(T5889_Y), .A(T4534_Y));
KC_INV_X1 T5888 ( .Y(T5888_Y), .A(T15934_Y));
KC_INV_X1 T5885 ( .Y(T5885_Y), .A(T5888_Y));
KC_INV_X1 T5884 ( .Y(T5884_Y), .A(T5156_Y));
KC_INV_X1 T15577 ( .Y(T15577_Y), .A(T6194_Co));
KC_INV_X1 T15988 ( .Y(T15988_Y), .A(T3876_Y));
KC_INV_X1 T15987 ( .Y(T15987_Y), .A(T4552_Y));
KC_INV_X1 T15966 ( .Y(T15966_Y), .A(T3876_Y));
KC_INV_X1 T15965 ( .Y(T15965_Y), .A(T4543_Y));
KC_INV_X1 T5980 ( .Y(T5980_Y), .A(T4560_Y));
KC_INV_X1 T5971 ( .Y(T5971_Y), .A(T5149_Y));
KC_INV_X1 T5969 ( .Y(T5969_Y), .A(T4551_Y));
KC_INV_X1 T5955 ( .Y(T5955_Y), .A(T12212_Y));
KC_INV_X1 T5954 ( .Y(T5954_Y), .A(T4576_Q));
KC_INV_X1 T5953 ( .Y(T5953_Y), .A(T11538_Y));
KC_INV_X1 T5952 ( .Y(T5952_Y), .A(T4578_Q));
KC_INV_X1 T5947 ( .Y(T5947_Y), .A(T11540_Y));
KC_INV_X1 T5946 ( .Y(T5946_Y), .A(T2757_Y));
KC_INV_X1 T15586 ( .Y(T15586_Y), .A(T4561_Y));
KC_INV_X1 T15584 ( .Y(T15584_Y), .A(T4575_Q));
KC_INV_X1 T16021 ( .Y(T16021_Y), .A(T8265_Y));
KC_INV_X1 T16020 ( .Y(T16020_Y), .A(T15605_Y));
KC_INV_X1 T16019 ( .Y(T16019_Y), .A(T3281_Y));
KC_INV_X1 T6022 ( .Y(T6022_Y), .A(T4602_Q));
KC_INV_X1 T6021 ( .Y(T6021_Y), .A(T4608_Q));
KC_INV_X1 T6019 ( .Y(T6019_Y), .A(T4611_Y));
KC_INV_X1 T6018 ( .Y(T6018_Y), .A(T11605_Y));
KC_INV_X1 T6016 ( .Y(T6016_Y), .A(T5158_Q));
KC_INV_X1 T6012 ( .Y(T6012_Y), .A(T4594_Y));
KC_INV_X1 T6010 ( .Y(T6010_Y), .A(T16019_Y));
KC_INV_X1 T6009 ( .Y(T6009_Y), .A(T6327_Y));
KC_INV_X1 T6008 ( .Y(T6008_Y), .A(T16021_Y));
KC_INV_X1 T15609 ( .Y(T15609_Y), .A(T11608_Y));
KC_INV_X1 T15604 ( .Y(T15604_Y), .A(T5159_Q));
KC_INV_X1 T16112 ( .Y(T16112_Y), .A(T11681_Y));
KC_INV_X1 T16111 ( .Y(T16111_Y), .A(T4669_Q));
KC_INV_X1 T16110 ( .Y(T16110_Y), .A(T6448_Y));
KC_INV_X1 T16045 ( .Y(T16045_Y), .A(T4703_Y));
KC_INV_X1 T6075 ( .Y(T6075_Y), .A(T5499_Q));
KC_INV_X1 T6057 ( .Y(T6057_Y), .A(T11705_Y));
KC_INV_X1 T6042 ( .Y(T6042_Y), .A(T12034_Y));
KC_INV_X1 T6030 ( .Y(T6030_Y), .A(T12031_Y));
KC_INV_X1 T6029 ( .Y(T6029_Y), .A(T3451_Y));
KC_INV_X1 T16122 ( .Y(T16122_Y), .A(T6129_Y));
KC_INV_X1 T8498 ( .Y(T8498_Y), .A(T10601_Y));
KC_INV_X1 T6171 ( .Y(T6171_Y), .A(T4713_Q));
KC_INV_X1 T6169 ( .Y(T6169_Y), .A(T4719_Q));
KC_INV_X1 T6148 ( .Y(T6148_Y), .A(T12277_Y));
KC_INV_X1 T6129 ( .Y(T6129_Y), .A(T4718_Q));
KC_INV_X1 T6126 ( .Y(T6126_Y), .A(T11707_Y));
KC_INV_X1 T6104 ( .Y(T6104_Y), .A(T5464_Y));
KC_INV_X1 T6103 ( .Y(T6103_Y), .A(T16460_Q));
KC_INV_X1 T6102 ( .Y(T6102_Y), .A(T4722_Q));
KC_INV_X1 T6091 ( .Y(T6091_Y), .A(T4723_Q));
KC_INV_X1 T6090 ( .Y(T6090_Y), .A(T4738_Y));
KC_INV_X1 T16146 ( .Y(T16146_Y), .A(T4704_Y));
KC_INV_X1 T6244 ( .Y(T6244_Y), .A(T4739_Y));
KC_INV_X1 T6234 ( .Y(T6234_Y), .A(T12308_Y));
KC_INV_X1 T6203 ( .Y(T6203_Y), .A(T4756_Q));
KC_INV_X1 T6202 ( .Y(T6202_Y), .A(T4757_Q));
KC_INV_X1 T6187 ( .Y(T6187_Y), .A(T4749_Y));
KC_INV_X1 T286 ( .Y(T286_Y), .A(T4758_Q));
KC_INV_X1 T15634 ( .Y(T15634_Y), .A(T6589_Y));
KC_INV_X1 T15630 ( .Y(T15630_Y), .A(T4755_Q));
KC_INV_X1 T15629 ( .Y(T15629_Y), .A(T4759_Q));
KC_INV_X1 T15625 ( .Y(T15625_Y), .A(T4760_Q));
KC_INV_X1 T16317 ( .Y(T16317_Y), .A(T8705_Y));
KC_INV_X1 T16314 ( .Y(T16314_Y), .A(T16316_Y));
KC_INV_X1 T16285 ( .Y(T16285_Y), .A(T9085_Y));
KC_INV_X1 T16284 ( .Y(T16284_Y), .A(T9080_S));
KC_INV_X1 T16283 ( .Y(T16283_Y), .A(T9084_Y));
KC_INV_X1 T6727 ( .Y(T6727_Y), .A(T166_Q));
KC_INV_X1 T16334 ( .Y(T16334_Y), .A(T7820_Y));
KC_INV_X1 T16332 ( .Y(T16332_Y), .A(T7825_Y));
KC_INV_X1 T16328 ( .Y(T16328_Y), .A(T7816_Y));
KC_INV_X1 T16325 ( .Y(T16325_Y), .A(T7826_Y));
KC_INV_X1 T16318 ( .Y(T16318_Y), .A(T7697_Y));
KC_INV_X1 T16287 ( .Y(T16287_Y), .A(T9447_Y));
KC_INV_X1 T16286 ( .Y(T16286_Y), .A(T9014_Y));
KC_INV_X1 T6728 ( .Y(T6728_Y), .A(T5275_Q));
KC_INV_X1 T16333 ( .Y(T16333_Y), .A(T7688_Y));
KC_INV_X1 T16187 ( .Y(T16187_Y), .A(T9243_Y));
KC_INV_X1 T6266 ( .Y(T6266_Y), .A(T434_Q));
KC_INV_X1 T6264 ( .Y(T6264_Y), .A(T440_Q));
KC_INV_X1 T285 ( .Y(T285_Y), .A(T5221_Q));
KC_INV_X1 T6700 ( .Y(T6700_Y), .A(T4836_Q));
KC_INV_X1 T15658 ( .Y(T15658_Y), .A(T781_Q));
KC_INV_X1 T6694 ( .Y(T6694_Y), .A(T886_Y));
KC_INV_X1 T6693 ( .Y(T6693_Y), .A(T6826_Y));
KC_INV_X1 T6250 ( .Y(T6250_Y), .A(T6289_Y));
KC_INV_X1 T16277 ( .Y(T16277_Y), .A(T8112_Y));
KC_INV_X1 T16400 ( .Y(T16400_Y), .A(T9896_Y));
KC_INV_X1 T16276 ( .Y(T16276_Y), .A(T16159_Y));
KC_INV_X1 T16275 ( .Y(T16275_Y), .A(T10942_Y));
KC_INV_X1 T16274 ( .Y(T16274_Y), .A(T10880_Y));
KC_INV_X1 T15663 ( .Y(T15663_Y), .A(T9897_Y));
KC_INV_X1 T15667 ( .Y(T15667_Y), .A(T5680_Y));
KC_INV_X1 T16398 ( .Y(T16398_Y), .A(T9994_Y));
KC_INV_X1 T16397 ( .Y(T16397_Y), .A(T8011_Y));
KC_INV_X1 T16396 ( .Y(T16396_Y), .A(T10010_Y));
KC_INV_X1 T16395 ( .Y(T16395_Y), .A(T16079_Q));
KC_INV_X1 T6791 ( .Y(T6791_Y), .A(T5663_Y));
KC_INV_X1 T15662 ( .Y(T15662_Y), .A(T12937_Y));
KC_INV_X1 T16373 ( .Y(T16373_Y), .A(T1691_Q));
KC_INV_X1 T16271 ( .Y(T16271_Y), .A(T10884_Y));
KC_INV_X1 T15974 ( .Y(T15974_Y), .A(T16156_Y));
KC_INV_X1 T15973 ( .Y(T15973_Y), .A(T10224_Y));
KC_INV_X1 T15904 ( .Y(T15904_Y), .A(T3415_Y));
KC_INV_X1 T6787 ( .Y(T6787_Y), .A(T10353_Y));
KC_INV_X1 T6786 ( .Y(T6786_Y), .A(T10335_Y));
KC_INV_X1 T6784 ( .Y(T6784_Y), .A(T10333_Y));
KC_INV_X1 T15666 ( .Y(T15666_Y), .A(T10364_Y));
KC_INV_X1 T16489 ( .Y(T16489_Y), .A(T11551_Y));
KC_INV_X1 T16371 ( .Y(T16371_Y), .A(T10525_Y));
KC_INV_X1 T16367 ( .Y(T16367_Y), .A(T10526_Y));
KC_INV_X1 T16366 ( .Y(T16366_Y), .A(T2001_Q));
KC_INV_X1 T16365 ( .Y(T16365_Y), .A(T10519_Y));
KC_INV_X1 T16364 ( .Y(T16364_Y), .A(T5369_Y));
KC_INV_X1 T16269 ( .Y(T16269_Y), .A(T5397_Q));
KC_INV_X1 T10258 ( .Y(T10258_Y), .A(T12111_Y));
KC_INV_X1 T16130 ( .Y(T16130_Y), .A(T12103_Y));
KC_INV_X1 T16129 ( .Y(T16129_Y), .A(T15713_Y));
KC_INV_X1 T16008 ( .Y(T16008_Y), .A(T16452_Y));
KC_INV_X1 T15859 ( .Y(T15859_Y), .A(T2689_Q));
KC_INV_X1 T6778 ( .Y(T6778_Y), .A(T14938_Q));
KC_INV_X1 T6777 ( .Y(T6777_Y), .A(T14937_Q));
KC_INV_X1 T6774 ( .Y(T6774_Y), .A(T1950_Y));
KC_INV_X1 T15713 ( .Y(T15713_Y), .A(T2285_Y));
KC_INV_X1 T15701 ( .Y(T15701_Y), .A(T5574_Q));
KC_INV_X1 T16404 ( .Y(T16404_Y), .A(T9743_Y));
KC_INV_X1 T16363 ( .Y(T16363_Y), .A(T2583_Q));
KC_INV_X1 T16362 ( .Y(T16362_Y), .A(T10061_Y));
KC_INV_X1 T16264 ( .Y(T16264_Y), .A(T2632_Y));
KC_INV_X1 T16181 ( .Y(T16181_Y), .A(T5548_Y));
KC_INV_X1 T16039 ( .Y(T16039_Y), .A(T15802_Q));
KC_INV_X1 T16038 ( .Y(T16038_Y), .A(T16034_Y));
KC_INV_X1 T15752 ( .Y(T15752_Y), .A(T2661_Y));
KC_INV_X1 T6773 ( .Y(T6773_Y), .A(T1949_Y));
KC_INV_X1 T6771 ( .Y(T6771_Y), .A(T10239_Y));
KC_INV_X1 T6764 ( .Y(T6764_Y), .A(T3039_Y));
KC_INV_X1 T6763 ( .Y(T6763_Y), .A(T3038_Y));
KC_INV_X1 T6545 ( .Y(T6545_Y), .A(T11564_Y));
KC_INV_X1 T287 ( .Y(T287_Y), .A(T6545_Y));
KC_INV_X1 T15689 ( .Y(T15689_Y), .A(T16181_Y));
KC_INV_X1 T15686 ( .Y(T15686_Y), .A(T14936_Q));
KC_INV_X1 T16405 ( .Y(T16405_Y), .A(T14884_Q));
KC_INV_X1 T16138 ( .Y(T16138_Y), .A(T11818_Y));
KC_INV_X1 T16137 ( .Y(T16137_Y), .A(T10550_Y));
KC_INV_X1 T16136 ( .Y(T16136_Y), .A(T10548_Y));
KC_INV_X1 T16135 ( .Y(T16135_Y), .A(T11816_Y));
KC_INV_X1 T16104 ( .Y(T16104_Y), .A(T12046_Y));
KC_INV_X1 T16037 ( .Y(T16037_Y), .A(T10965_Y));
KC_INV_X1 T16035 ( .Y(T16035_Y), .A(T6555_Q));
KC_INV_X1 T15997 ( .Y(T15997_Y), .A(T3294_Y));
KC_INV_X1 T15863 ( .Y(T15863_Y), .A(T14543_Q));
KC_INV_X1 T15699 ( .Y(T15699_Y), .A(T14541_Q));
KC_INV_X1 T15688 ( .Y(T15688_Y), .A(T2469_Y));
KC_INV_X1 T16141 ( .Y(T16141_Y), .A(T11745_Y));
KC_INV_X1 T16140 ( .Y(T16140_Y), .A(T11683_Y));
KC_INV_X1 T16107 ( .Y(T16107_Y), .A(T4059_Y));
KC_INV_X1 T16106 ( .Y(T16106_Y), .A(T4015_Y));
KC_INV_X1 T15996 ( .Y(T15996_Y), .A(T15878_Y));
KC_INV_X1 T15995 ( .Y(T15995_Y), .A(T11616_Y));
KC_INV_X1 T15971 ( .Y(T15971_Y), .A(T3974_Q));
KC_INV_X1 T15907 ( .Y(T15907_Y), .A(T16153_Y));
KC_INV_X1 T15868 ( .Y(T15868_Y), .A(T3836_Y));
KC_INV_X1 T15709 ( .Y(T15709_Y), .A(T5116_Y));
KC_INV_X1 T15705 ( .Y(T15705_Y), .A(T6340_Y));
KC_INV_X1 T16444 ( .Y(T16444_Y), .A(T4312_Y));
KC_INV_X1 T16145 ( .Y(T16145_Y), .A(T4736_Y));
KC_INV_X1 T16144 ( .Y(T16144_Y), .A(T4735_Y));
KC_INV_X1 T15969 ( .Y(T15969_Y), .A(T11505_Y));
KC_INV_X1 T15968 ( .Y(T15968_Y), .A(T5141_Y));
KC_INV_X1 T15967 ( .Y(T15967_Y), .A(T11539_Y));
KC_INV_X1 T15964 ( .Y(T15964_Y), .A(T4568_Q));
KC_INV_X1 T15938 ( .Y(T15938_Y), .A(T12461_Y));
KC_INV_X1 T15824 ( .Y(T15824_Y), .A(T15555_Y));
KC_INV_X1 T15706 ( .Y(T15706_Y), .A(T4519_Y));
KC_INV_X1 T15704 ( .Y(T15704_Y), .A(T12833_Y));
KC_INV_X1 T15703 ( .Y(T15703_Y), .A(T4579_Q));
KC_INV_X1 T304 ( .Y(T304_Y), .A(T442_Q));
KC_INV_X1 T15351 ( .Y(T15351_Y), .A(T436_Q));
KC_INV_X1 T6595 ( .Y(T6595_Y), .A(T3071_Y));
KC_INV_X1 T6652 ( .Y(T6652_Y), .A(T7551_Y));
KC_INV_X1 T8713 ( .Y(T8713_Y), .A(T7593_Y));
KC_INV_X1 T730 ( .Y(T730_Y), .A(T8724_Y));
KC_INV_X1 T659 ( .Y(T659_Y), .A(T669_Q));
KC_INV_X1 T1081 ( .Y(T1081_Y), .A(T7945_Y));
KC_INV_X1 T969 ( .Y(T969_Y), .A(T11264_Y));
KC_INV_X1 T930 ( .Y(T930_Y), .A(T8794_Y));
KC_INV_X1 T1330 ( .Y(T1330_Y), .A(T613_Y));
KC_INV_X1 T1323 ( .Y(T1323_Y), .A(T751_Q));
KC_INV_X1 T15525 ( .Y(T15525_Y), .A(T9496_Y));
KC_INV_X1 T5735 ( .Y(T5735_Y), .A(T10536_Y));
KC_INV_X1 T5730 ( .Y(T5730_Y), .A(T10537_Y));
KC_INV_X1 T15865 ( .Y(T15865_Y), .A(T3840_Y));
KC_INV_X1 T15853 ( .Y(T15853_Y), .A(T15844_Q));
KC_INV_X1 T15886 ( .Y(T15886_Y), .A(T2741_Y));
KC_INV_X1 T5795 ( .Y(T5795_Y), .A(T4452_Y));
KC_INV_X1 T15916 ( .Y(T15916_Y), .A(T3411_Y));
KC_INV_X1 T5861 ( .Y(T5861_Y), .A(T2731_Y));
KC_INV_X1 T5852 ( .Y(T5852_Y), .A(T14551_Q));
KC_INV_X1 T15959 ( .Y(T15959_Y), .A(T11479_Y));
KC_INV_X1 T15943 ( .Y(T15943_Y), .A(T3411_Y));
KC_INV_X1 T5895 ( .Y(T5895_Y), .A(T11488_Y));
KC_INV_X1 T15970 ( .Y(T15970_Y), .A(T16202_Y));
KC_INV_X1 T15592 ( .Y(T15592_Y), .A(T11536_Y));
KC_INV_X1 T15590 ( .Y(T15590_Y), .A(T5480_Q));
KC_INV_X1 T6015 ( .Y(T6015_Y), .A(T10959_Y));
KC_INV_X1 T6087 ( .Y(T6087_Y), .A(T3517_Y));
KC_INV_X1 T6066 ( .Y(T6066_Y), .A(T5490_Y));
KC_INV_X1 T6055 ( .Y(T6055_Y), .A(T2843_Q));
KC_INV_X1 T6184 ( .Y(T6184_Y), .A(T12270_Y));
KC_INV_X1 T6178 ( .Y(T6178_Y), .A(T5056_Y));
KC_INV_X1 T15623 ( .Y(T15623_Y), .A(T15233_Y));
KC_INV_X1 T15621 ( .Y(T15621_Y), .A(T5523_Y));
KC_INV_X1 T6565 ( .Y(T6565_Y), .A(T1829_Q));
KC_INV_X1 T6560 ( .Y(T6560_Y), .A(T10999_Y));
KC_INV_X1 T6240 ( .Y(T6240_Y), .A(T12101_Y));
KC_INV_X1 T6238 ( .Y(T6238_Y), .A(T2888_Y));
KC_INV_X1 T6200 ( .Y(T6200_Y), .A(T1833_Q));
KC_INV_X1 T6257 ( .Y(T6257_Y), .A(T822_Q));
KC_XNOR2_X3 T15147 ( .Y(T15147_Y), .A(T2071_Y), .B(T9427_Y));
KC_XNOR2_X3 T15146 ( .Y(T15146_Y), .A(T8928_Y), .B(T9428_Y));
KC_XNOR2_X3 T15145 ( .Y(T15145_Y), .A(T8092_Y), .B(T9426_Y));
KC_XNOR2_X3 T15144 ( .Y(T15144_Y), .A(T8881_Y), .B(T9430_Y));
KC_XNOR2_X3 T15066 ( .Y(T15066_Y), .A(T7914_Y), .B(T8875_Y));
KC_XNOR2_X3 T15065 ( .Y(T15065_Y), .A(T8884_Y), .B(T8876_Y));
KC_XNOR2_X3 T15064 ( .Y(T15064_Y), .A(T8824_Y), .B(T8885_Y));
KC_XNOR2_X3 T15063 ( .Y(T15063_Y), .A(T8842_Y), .B(T8839_Y));
KC_XNOR2_X3 T15062 ( .Y(T15062_Y), .A(T8879_Y), .B(T8817_Y));
KC_XNOR2_X3 T15061 ( .Y(T15061_Y), .A(T8840_Y), .B(T8816_Y));
KC_XNOR2_X3 T15060 ( .Y(T15060_Y), .A(T7865_Y), .B(T8819_Y));
KC_XNOR2_X3 T15059 ( .Y(T15059_Y), .A(T7914_Y), .B(T8820_Y));
KC_XNOR2_X3 T15058 ( .Y(T15058_Y), .A(T7920_Y), .B(T8822_Y));
KC_XNOR2_X3 T15057 ( .Y(T15057_Y), .A(T7920_Y), .B(T8818_Y));
KC_XNOR2_X3 T16064 ( .Y(T16064_Y), .A(T8968_Y), .B(T8955_Y));
KC_XNOR2_X3 T15083 ( .Y(T15083_Y), .A(T8055_Y), .B(T8952_Y));
KC_XNOR2_X3 T15082 ( .Y(T15082_Y), .A(T8090_Y), .B(T8953_Y));
KC_XNOR2_X3 T15081 ( .Y(T15081_Y), .A(T8971_Y), .B(T8961_Y));
KC_XNOR2_X3 T15080 ( .Y(T15080_Y), .A(T8958_Y), .B(T8954_Y));
KC_XNOR2_X3 T15079 ( .Y(T15079_Y), .A(T7874_Y), .B(T8930_Y));
KC_XNOR2_X3 T15078 ( .Y(T15078_Y), .A(T8957_Y), .B(T8919_Y));
KC_XNOR2_X3 T15077 ( .Y(T15077_Y), .A(T15081_Y), .B(T8931_Y));
KC_XNOR2_X3 T15076 ( .Y(T15076_Y), .A(T2071_Y), .B(T8921_Y));
KC_XNOR2_X3 T15075 ( .Y(T15075_Y), .A(T2277_Y), .B(T8920_Y));
KC_XNOR2_X3 T15100 ( .Y(T15100_Y), .A(T1523_Y), .B(T9175_Y));
KC_XNOR2_X3 T15099 ( .Y(T15099_Y), .A(T9250_Y), .B(T9176_Y));
KC_XNOR2_X3 T15098 ( .Y(T15098_Y), .A(T5415_Y), .B(T9177_Y));
KC_XNOR2_X3 T15096 ( .Y(T15096_Y), .A(T15097_Y), .B(T9153_Y));
KC_XNOR2_X3 T15095 ( .Y(T15095_Y), .A(T9214_Y), .B(T9155_Y));
KC_XNOR2_X3 T15094 ( .Y(T15094_Y), .A(T9236_Y), .B(T9154_Y));
KC_XNOR2_X3 T15093 ( .Y(T15093_Y), .A(T1016_Y), .B(T9130_Y));
KC_XNOR2_X3 T15092 ( .Y(T15092_Y), .A(T9082_Y), .B(T9131_Y));
KC_XNOR2_X3 T15091 ( .Y(T15091_Y), .A(T1016_Y), .B(T9081_Y));
KC_XNOR2_X3 T15119 ( .Y(T15119_Y), .A(T591_Y), .B(T9246_Y));
KC_XNOR2_X3 T15118 ( .Y(T15118_Y), .A(T1167_Y), .B(T9247_Y));
KC_XNOR2_X3 T15117 ( .Y(T15117_Y), .A(T9203_Y), .B(T9245_Y));
KC_XNOR2_X3 T15115 ( .Y(T15115_Y), .A(T9201_Y), .B(T9235_Y));
KC_XNOR2_X3 T15114 ( .Y(T15114_Y), .A(T9212_Y), .B(T9231_Y));
KC_XNOR2_X3 T15113 ( .Y(T15113_Y), .A(T9207_Y), .B(T9234_Y));
KC_XNOR2_X3 T15112 ( .Y(T15112_Y), .A(T9205_Y), .B(T9233_Y));
KC_XNOR2_X3 T15111 ( .Y(T15111_Y), .A(T9204_Y), .B(T9232_Y));
KC_XNOR2_X3 T15107 ( .Y(T15107_Y), .A(T9236_Y), .B(T9200_Y));
KC_XNOR2_X3 T15143 ( .Y(T15143_Y), .A(T8923_Y), .B(T9429_Y));
KC_XNOR2_X3 T15056 ( .Y(T15056_Y), .A(T8869_Y), .B(T8821_Y));
KC_XNOR2_X3 T15074 ( .Y(T15074_Y), .A(T8972_Y), .B(T8918_Y));
KC_XNOR2_X3 T15151 ( .Y(T15151_Y), .A(T9492_Y), .B(T9480_Y));
KC_XNOR2_X3 T15150 ( .Y(T15150_Y), .A(T425_Y), .B(T9479_Y));
KC_XNOR2_X3 T15148 ( .Y(T15148_Y), .A(T9493_Y), .B(T9473_Y));
KC_XNOR2_X3 T15097 ( .Y(T15097_Y), .A(T9216_Y), .B(T9167_Y));
KC_XNOR2_X3 T15116 ( .Y(T15116_Y), .A(T426_Y), .B(T9244_Y));
KC_XNOR2_X3 T15110 ( .Y(T15110_Y), .A(T591_Y), .B(T9228_Y));
KC_XNOR2_X3 T15109 ( .Y(T15109_Y), .A(T425_Y), .B(T9229_Y));
KC_XNOR2_X3 T15108 ( .Y(T15108_Y), .A(T9197_Y), .B(T9230_Y));
KC_XNOR2_X3 T15106 ( .Y(T15106_Y), .A(T9215_Y), .B(T9195_Y));
KC_XNOR2_X3 T15105 ( .Y(T15105_Y), .A(T9214_Y), .B(T9196_Y));
KC_XNOR2_X3 T15104 ( .Y(T15104_Y), .A(T606_Q), .B(T9192_Y));
KC_XNOR2_X3 T15103 ( .Y(T15103_Y), .A(T606_Q), .B(T9189_Y));
KC_XNOR2_X3 T15102 ( .Y(T15102_Y), .A(T15891_Q), .B(T9191_Y));
KC_XNOR2_X3 T15046 ( .Y(T15046_Y), .A(T840_Y), .B(T8615_Y));
KC_XNOR2_X3 T15120 ( .Y(T15120_Y), .A(T2114_Q), .B(T10229_Y));
KC_XNOR2_X3 T15073 ( .Y(T15073_Y), .A(T10531_Y), .B(T9975_Y));
KC_XNOR2_X3 T15071 ( .Y(T15071_Y), .A(T5366_Q), .B(T9942_Y));
KC_XNOR2_X3 T15067 ( .Y(T15067_Y), .A(T1709_Y), .B(T9881_Y));
KC_XNOR2_X3 T15087 ( .Y(T15087_Y), .A(T15531_Y), .B(T10029_Y));
KC_XNOR2_X3 T15086 ( .Y(T15086_Y), .A(T16271_Y), .B(T10030_Y));
KC_XNOR2_X3 T15053 ( .Y(T15053_Y), .A(T13008_Q), .B(T9840_Y));
KC_XNOR2_X3 T15052 ( .Y(T15052_Y), .A(T5311_Q), .B(T9842_Y));
KC_XNOR2_X3 T15051 ( .Y(T15051_Y), .A(T13013_Q), .B(T9841_Y));
KC_XNOR2_X3 T15089 ( .Y(T15089_Y), .A(T10107_Y), .B(T10081_Y));
KC_XNOR2_X3 T15039 ( .Y(T15039_Y), .A(T12794_Y), .B(T8191_Y));
KC_XNOR2_X3 T15125 ( .Y(T15125_Y), .A(T11489_Y), .B(T8210_Y));
KC_XNOR2_X3 T15164 ( .Y(T15164_Y), .A(T15608_Y), .B(T8483_Y));
KC_XNOR2_X3 T15140 ( .Y(T15140_Y), .A(T8410_Y), .B(T8419_Y));
KC_XNOR2_X3 T15142 ( .Y(T15142_Y), .A(T6605_Y), .B(T8158_Y));
KC_XNOR2_X3 T15055 ( .Y(T15055_Y), .A(T5314_Y), .B(T9872_Y));
KC_XNOR2_X3 T15050 ( .Y(T15050_Y), .A(T9743_Y), .B(T9835_Y));
KC_XNOR2_X3 T15155 ( .Y(T15155_Y), .A(T6676_Y), .B(T10514_Y));
KC_XNOR2_X3 T15090 ( .Y(T15090_Y), .A(T14404_Q), .B(T10119_Y));
KC_XNOR2_X3 T15088 ( .Y(T15088_Y), .A(T14303_Q), .B(T10054_Y));
KC_XNOR2_X3 T15129 ( .Y(T15129_Y), .A(T3260_Y), .B(T8231_Y));
KC_XNOR2_X3 T15127 ( .Y(T15127_Y), .A(T3280_Y), .B(T8214_Y));
KC_XNOR2_X3 T15162 ( .Y(T15162_Y), .A(T3332_Y), .B(T8479_Y));
KC_XNOR2_X3 T15131 ( .Y(T15131_Y), .A(T8239_Y), .B(T8292_Y));
KC_XNOR2_X3 T15134 ( .Y(T15134_Y), .A(T3346_Y), .B(T8336_Y));
KC_XNOR2_X3 T15133 ( .Y(T15133_Y), .A(T6335_Y), .B(T8314_Y));
KC_XNOR2_X3 T15054 ( .Y(T15054_Y), .A(T13011_Y), .B(T9871_Y));
KC_XNOR2_X3 T15128 ( .Y(T15128_Y), .A(T3265_Y), .B(T8221_Y));
KC_XNOR2_X3 T15126 ( .Y(T15126_Y), .A(T5859_Y), .B(T8212_Y));
KC_XNOR2_X3 T15130 ( .Y(T15130_Y), .A(T3934_Y), .B(T8245_Y));
KC_XNOR2_X3 T15163 ( .Y(T15163_Y), .A(T16417_Y), .B(T8476_Y));
KC_XNOR2_X3 T15157 ( .Y(T15157_Y), .A(T3793_Y), .B(T8438_Y));
KC_XNOR2_X3 T15156 ( .Y(T15156_Y), .A(T5169_Y), .B(T8439_Y));
KC_XNOR2_X3 T15121 ( .Y(T15121_Y), .A(T15157_Y), .B(T8177_Y));
KC_XNOR2_X3 T15132 ( .Y(T15132_Y), .A(T4623_Y), .B(T8299_Y));
KC_XNOR2_X3 T15135 ( .Y(T15135_Y), .A(T6029_Y), .B(T8365_Y));
KC_XNOR2_X3 T15136 ( .Y(T15136_Y), .A(T13169_Y), .B(T8383_Y));
KC_XNOR2_X3 T15149 ( .Y(T15149_Y), .A(T9248_Y), .B(T9481_Y));
KC_XNOR2_X3 T15152 ( .Y(T15152_Y), .A(T13941_Q), .B(T10321_Y));
KC_XNOR2_X3 T15161 ( .Y(T15161_Y), .A(T15894_Q), .B(T8454_Y));
KC_XNOR2_X3 T15154 ( .Y(T15154_Y), .A(T4983_Y), .B(T10510_Y));
KC_XNOR2_X3 T15153 ( .Y(T15153_Y), .A(T5312_Y), .B(T10511_Y));
KC_XNOR2_X3 T15042 ( .Y(T15042_Y), .A(T11038_Y), .B(T8169_Y));
KC_XNOR2_X3 T15043 ( .Y(T15043_Y), .A(T11036_Y), .B(T8168_Y));
KC_XNOR2_X3 T15160 ( .Y(T15160_Y), .A(T6074_Y), .B(T8449_Y));
KC_XNOR2_X3 T15158 ( .Y(T15158_Y), .A(T16157_Y), .B(T8437_Y));
KC_XNOR2_X3 T15069 ( .Y(T15069_Y), .A(T15463_Y), .B(T9901_Y));
KC_XNOR2_X3 T15101 ( .Y(T15101_Y), .A(T15891_Q), .B(T9190_Y));
KC_XNOR2_X3 T15159 ( .Y(T15159_Y), .A(T3822_Y), .B(T8443_Y));
KC_TLAT_X1 T13332 ( .B(T15323_Y), .Q(T13332_Q), .CK(T14982_Y),     .A(T5622_Y));
KC_TLAT_X1 T13330 ( .B(T16490_Y), .Q(T13330_Q), .CK(T13288_Y),     .A(T8539_Y));
KC_TLAT_X1 T13440 ( .B(T15337_Y), .Q(T13440_Q), .CK(T4841_Y),     .A(T8568_Y));
KC_TLAT_X1 T13936 ( .B(T785_Y), .Q(T13936_Q), .CK(T16476_Y),     .A(T11886_Y));
KC_TLAT_X1 T13935 ( .B(T15651_Y), .Q(T13935_Q), .CK(T4849_Y),     .A(T9341_Y));
KC_TLAT_X1 T13934 ( .B(T785_Y), .Q(T13934_Q), .CK(T706_Y),     .A(T11217_Y));
KC_TLAT_X1 T13933 ( .B(T16175_Y), .Q(T13933_Q), .CK(T943_Y),     .A(T8733_Y));
KC_TLAT_X1 T13932 ( .B(T15651_Y), .Q(T13932_Q), .CK(T943_Y),     .A(T9342_Y));
KC_TLAT_X1 T14096 ( .B(T15456_Y), .Q(T14096_Q), .CK(T942_Y),     .A(T11887_Y));
KC_TLAT_X1 T14094 ( .B(T15456_Y), .Q(T14094_Q), .CK(T15175_Y),     .A(T11888_Y));
KC_TLAT_X1 T14588 ( .B(T643_Y), .Q(T14588_Q), .CK(T4849_Y),     .A(T12442_Y));
KC_TLAT_X1 T14097 ( .B(T16175_Y), .Q(T14097_Q), .CK(T4849_Y),     .A(T8734_Y));
KC_TLAT_X1 T14095 ( .B(T885_Y), .Q(T14095_Q), .CK(T942_Y),     .A(T7842_Y));
KC_TLAT_X1 T14203 ( .B(T16300_Y), .Q(T14203_Q), .CK(T13288_Y),     .A(T9000_Y));
KC_TLAT_X1 T14202 ( .B(T15481_Y), .Q(T14202_Q), .CK(T774_Y),     .A(T8892_Y));
KC_TLAT_X1 T14201 ( .B(T15482_Y), .Q(T14201_Q), .CK(T1105_Y),     .A(T11263_Y));
KC_TLAT_X1 T14200 ( .B(T15456_Y), .Q(T14200_Q), .CK(T15173_Y),     .A(T16463_Y));
KC_TLAT_X1 T14370 ( .B(T15521_Y), .Q(T14370_Q), .CK(T15185_Y),     .A(T12887_Y));
KC_TLAT_X1 T14369 ( .B(T15522_Y), .Q(T14369_Q), .CK(T991_Y),     .A(T1010_Y));
KC_TLAT_X1 T14137 ( .B(T15465_Y), .Q(T14137_Q), .CK(T16415_Y),     .A(T16431_Y));
KC_TLAT_X1 T14216 ( .B(T15521_Y), .Q(T14216_Q), .CK(T1137_Y),     .A(T12891_Y));
KC_TLAT_X1 T14199 ( .B(T15465_Y), .Q(T14199_Q), .CK(T16415_Y),     .A(T1099_Y));
KC_TLAT_X1 T13467 ( .B(T15340_Y), .Q(T13467_Q), .CK(T1325_Y),     .A(T1409_Y));
KC_TLAT_X1 T14643 ( .B(T15418_Y), .Q(T14643_Q), .CK(T5361_Y),     .A(T12577_Y));
KC_TLAT_X1 T14642 ( .B(T15418_Y), .Q(T14642_Q), .CK(T5361_Y),     .A(T595_Y));
KC_TLAT_X1 T13376 ( .B(T15343_Y), .Q(T13376_Q), .CK(T1403_Y),     .A(T312_Y));
KC_TLAT_X1 T13347 ( .B(T15343_Y), .Q(T13347_Q), .CK(T1324_Y),     .A(T12908_Y));
KC_TLAT_X1 T13346 ( .B(T15340_Y), .Q(T13346_Q), .CK(T1324_Y),     .A(T314_Y));
KC_TLAT_X1 T14693 ( .B(T15361_Y), .Q(T14693_Q), .CK(T1325_Y),     .A(T6441_Y));
KC_TLAT_X1 T13608 ( .B(T15360_Y), .Q(T13608_Q), .CK(T1963_Y),     .A(T1408_Y));
KC_TLAT_X1 T14638 ( .B(T588_Y), .Q(T14638_Q), .CK(T5361_Y),     .A(T6823_Y));
KC_TLAT_X1 T13858 ( .B(T15417_Y), .Q(T13858_Q), .CK(T5361_Y),     .A(T1347_Y));
KC_TLAT_X1 T13857 ( .B(T15417_Y), .Q(T13857_Q), .CK(T5361_Y),     .A(T6837_Y));
KC_TLAT_X1 T13856 ( .B(T15418_Y), .Q(T13856_Q), .CK(T5361_Y),     .A(T12586_Y));
KC_TLAT_X1 T13815 ( .B(T15418_Y), .Q(T13815_Q), .CK(T5361_Y),     .A(T1452_Y));
KC_TLAT_X1 T13793 ( .B(T15417_Y), .Q(T13793_Q), .CK(T5361_Y),     .A(T6836_Y));
KC_TLAT_X1 T13792 ( .B(T15417_Y), .Q(T13792_Q), .CK(T5361_Y),     .A(T1348_Y));
KC_TLAT_X1 T13791 ( .B(T15418_Y), .Q(T13791_Q), .CK(T5361_Y),     .A(T12585_Y));
KC_TLAT_X1 T14276 ( .B(T15493_Y), .Q(T14276_Q), .CK(T13261_Y),     .A(T12977_Y));
KC_TLAT_X1 T14227 ( .B(T15528_Y), .Q(T14227_Q), .CK(T1356_Y),     .A(T10131_Y));
KC_TLAT_X1 T14212 ( .B(T15530_Y), .Q(T14212_Q), .CK(T13261_Y),     .A(T12978_Y));
KC_TLAT_X1 T13345 ( .B(T15339_Y), .Q(T13345_Q), .CK(T1325_Y),     .A(T12482_Y));
KC_TLAT_X1 T14691 ( .B(T15360_Y), .Q(T14691_Q), .CK(T1963_Y),     .A(T12485_Y));
KC_TLAT_X1 T14690 ( .B(T15360_Y), .Q(T14690_Q), .CK(T1963_Y),     .A(T1407_Y));
KC_TLAT_X1 T14689 ( .B(T15360_Y), .Q(T14689_Q), .CK(T1324_Y),     .A(T1406_Y));
KC_TLAT_X1 T14688 ( .B(T15360_Y), .Q(T14688_Q), .CK(T1963_Y),     .A(T12483_Y));
KC_TLAT_X1 T13496 ( .B(T15339_Y), .Q(T13496_Q), .CK(T1325_Y),     .A(T12481_Y));
KC_TLAT_X1 T13495 ( .B(T15361_Y), .Q(T13495_Q), .CK(T1525_Y),     .A(T1404_Y));
KC_TLAT_X1 T13466 ( .B(T15361_Y), .Q(T13466_Q), .CK(T1324_Y),     .A(T6442_Y));
KC_TLAT_X1 T13448 ( .B(T15361_Y), .Q(T13448_Q), .CK(T1325_Y),     .A(T1410_Y));
KC_TLAT_X1 T14659 ( .B(T588_Y), .Q(T14659_Q), .CK(T5361_Y),     .A(T12579_Y));
KC_TLAT_X1 T14012 ( .B(T818_Y), .Q(T14012_Q), .CK(T1560_Y),     .A(T850_Y));
KC_TLAT_X1 T13957 ( .B(T818_Y), .Q(T13957_Q), .CK(T1560_Y),     .A(T12635_Y));
KC_TLAT_X1 T14270 ( .B(T15495_Y), .Q(T14270_Q), .CK(T13261_Y),     .A(T12730_Y));
KC_TLAT_X1 T14253 ( .B(T15495_Y), .Q(T14253_Q), .CK(T13261_Y),     .A(T1502_Y));
KC_TLAT_X1 T14252 ( .B(T15661_Y), .Q(T14252_Q), .CK(T13261_Y),     .A(T1500_Y));
KC_TLAT_X1 T14251 ( .B(T15495_Y), .Q(T14251_Q), .CK(T13261_Y),     .A(T12729_Y));
KC_TLAT_X1 T14250 ( .B(T15661_Y), .Q(T14250_Q), .CK(T13261_Y),     .A(T1501_Y));
KC_TLAT_X1 T14236 ( .B(T15495_Y), .Q(T14236_Q), .CK(T13261_Y),     .A(T16307_Y));
KC_TLAT_X1 T14225 ( .B(T15495_Y), .Q(T14225_Q), .CK(T13261_Y),     .A(T1504_Y));
KC_TLAT_X1 T14224 ( .B(T15493_Y), .Q(T14224_Q), .CK(T13261_Y),     .A(T1507_Y));
KC_TLAT_X1 T14210 ( .B(T15493_Y), .Q(T14210_Q), .CK(T1510_Y),     .A(T16298_Y));
KC_TLAT_X1 T14209 ( .B(T15494_Y), .Q(T14209_Q), .CK(T13261_Y),     .A(T16273_Y));
KC_TLAT_X1 T14591 ( .B(T15542_Y), .Q(T14591_Q), .CK(T13261_Y),     .A(T12727_Y));
KC_TLAT_X1 T13329 ( .B(T15542_Y), .Q(T13329_Q), .CK(T13261_Y),     .A(T16272_Y));
KC_TLAT_X1 T14677 ( .B(T15668_Y), .Q(T14677_Q), .CK(T1525_Y),     .A(T1520_Y));
KC_TLAT_X1 T13340 ( .B(T15668_Y), .Q(T13340_Q), .CK(T1525_Y),     .A(T1401_Y));
KC_TLAT_X1 T13492 ( .B(T15344_Y), .Q(T13492_Q), .CK(T1525_Y),     .A(T12907_Y));
KC_TLAT_X1 T13491 ( .B(T15341_Y), .Q(T13491_Q), .CK(T1525_Y),     .A(T12486_Y));
KC_TLAT_X1 T13490 ( .B(T15359_Y), .Q(T13490_Q), .CK(T1525_Y),     .A(T6439_Y));
KC_TLAT_X1 T13478 ( .B(T15339_Y), .Q(T13478_Q), .CK(T1525_Y),     .A(T12490_Y));
KC_TLAT_X1 T13464 ( .B(T15359_Y), .Q(T13464_Q), .CK(T1963_Y),     .A(T5218_Y));
KC_TLAT_X1 T13446 ( .B(T15359_Y), .Q(T13446_Q), .CK(T1963_Y),     .A(T12479_Y));
KC_TLAT_X1 T13445 ( .B(T15341_Y), .Q(T13445_Q), .CK(T1525_Y),     .A(T12488_Y));
KC_TLAT_X1 T13804 ( .B(T818_Y), .Q(T13804_Q), .CK(T1560_Y),     .A(T1459_Y));
KC_TLAT_X1 T14008 ( .B(T16180_Y), .Q(T14008_Q), .CK(T1560_Y),     .A(T12630_Y));
KC_TLAT_X1 T13953 ( .B(T15437_Y), .Q(T13953_Q), .CK(T1560_Y),     .A(T1552_Y));
KC_TLAT_X1 T13952 ( .B(T15437_Y), .Q(T13952_Q), .CK(T1560_Y),     .A(T12616_Y));
KC_TLAT_X1 T13940 ( .B(T849_Y), .Q(T13940_Q), .CK(T1560_Y),     .A(T12628_Y));
KC_TLAT_X1 T13939 ( .B(T849_Y), .Q(T13939_Q), .CK(T1560_Y),     .A(T1553_Y));
KC_TLAT_X1 T14683 ( .B(T15668_Y), .Q(T14683_Q), .CK(T1963_Y),     .A(T12487_Y));
KC_TLAT_X1 T14682 ( .B(T15344_Y), .Q(T14682_Q), .CK(T1963_Y),     .A(T5183_Y));
KC_TLAT_X1 T13642 ( .B(T15669_Y), .Q(T13642_Q), .CK(T1963_Y),     .A(T6445_Y));
KC_TLAT_X1 T14865 ( .B(T15437_Y), .Q(T14865_Q), .CK(T1560_Y),     .A(T1557_Y));
KC_TLAT_X1 T13951 ( .B(T15437_Y), .Q(T13951_Q), .CK(T1560_Y),     .A(T830_Y));
KC_TLAT_X1 T14554 ( .B(T15698_Y), .Q(T14554_Q), .CK(T2157_Y),     .A(T15038_Y));
KC_TLAT_X1 T13757 ( .B(T15669_Y), .Q(T13757_Q), .CK(T1963_Y),     .A(T1526_Y));
KC_TLAT_X1 T13745 ( .B(T15669_Y), .Q(T13745_Q), .CK(T1963_Y),     .A(T6446_Y));
KC_TLAT_X1 T14174 ( .B(T15479_Y), .Q(T14174_Q), .CK(T15188_Y),     .A(T2010_Y));
KC_TLAT_X1 T14173 ( .B(T15479_Y), .Q(T14173_Q), .CK(T5423_Y),     .A(T12092_Y));
KC_TLAT_X1 T14368 ( .B(T15690_Y), .Q(T14368_Q), .CK(T15174_Y),     .A(T10248_Y));
KC_TLAT_X1 T14326 ( .B(T1139_Y), .Q(T14326_Q), .CK(T16446_Q),     .A(T2567_Y));
KC_TLAT_X1 T14960 ( .B(T15575_Y), .Q(T14960_Q), .CK(T2156_Y),     .A(T13109_Y));
KC_TLAT_X1 T14557 ( .B(T15575_Y), .Q(T14557_Q), .CK(T13268_Y),     .A(T2155_Y));
KC_TLAT_X1 T14565 ( .B(T15583_Y), .Q(T14565_Q), .CK(T2157_Y),     .A(T2185_Y));
KC_TLAT_X1 T14564 ( .B(T15950_Y), .Q(T14564_Q), .CK(T2157_Y),     .A(T2176_Y));
KC_TLAT_X1 T14560 ( .B(T15950_Y), .Q(T14560_Q), .CK(T2157_Y),     .A(T11500_Y));
KC_TLAT_X1 T14559 ( .B(T15583_Y), .Q(T14559_Q), .CK(T2157_Y),     .A(T11517_Y));
KC_TLAT_X1 T14558 ( .B(T15583_Y), .Q(T14558_Q), .CK(T2157_Y),     .A(T8493_Y));
KC_TLAT_X1 T14577 ( .B(T6554_Y), .Q(T14577_Q), .CK(T15192_Y),     .A(T2327_Y));
KC_TLAT_X1 T14185 ( .B(T15475_Y), .Q(T14185_Q), .CK(T5423_Y),     .A(T2613_Y));
KC_TLAT_X1 T14304 ( .B(T15505_Y), .Q(T14304_Q), .CK(T15188_Y),     .A(T10056_Y));
KC_TLAT_X1 T14481 ( .B(T15547_Y), .Q(T14481_Q), .CK(T3217_Y),     .A(T12127_Y));
KC_TLAT_X1 T14566 ( .B(T16452_Y), .Q(T14566_Q), .CK(T2790_Y),     .A(T11563_Y));
KC_TLAT_X1 T14572 ( .B(T11548_Y), .Q(T14572_Q), .CK(VDD),     .A(T16456_Y));
KC_TLAT_X1 T14571 ( .B(T11548_Y), .Q(T14571_Q), .CK(VDD),     .A(T16452_Y));
KC_TLAT_X1 T14570 ( .B(T15603_Y), .Q(T14570_Q), .CK(T2813_Y),     .A(T2801_Y));
KC_TLAT_X1 T14961 ( .B(T15710_Y), .Q(T14961_Q), .CK(T15192_Y),     .A(T11030_Y));
KC_TLAT_X1 T14573 ( .B(T15614_Y), .Q(T14573_Q), .CK(T15192_Y),     .A(T11031_Y));
KC_TLAT_X1 T14581 ( .B(T15644_Y), .Q(T14581_Q), .CK(T15192_Y),     .A(T11685_Y));
KC_TLAT_X1 T14080 ( .B(T15449_Y), .Q(T14080_Q), .CK(T3075_Y),     .A(T12646_Y));
KC_TLAT_X1 T14079 ( .B(T15449_Y), .Q(T14079_Q), .CK(T3075_Y),     .A(T12667_Y));
KC_TLAT_X1 T14078 ( .B(T15446_Y), .Q(T14078_Q), .CK(T3075_Y),     .A(T12666_Y));
KC_TLAT_X1 T14077 ( .B(T15449_Y), .Q(T14077_Q), .CK(T3075_Y),     .A(T12645_Y));
KC_TLAT_X1 T14076 ( .B(T15449_Y), .Q(T14076_Q), .CK(T3075_Y),     .A(T12644_Y));
KC_TLAT_X1 T14031 ( .B(T15449_Y), .Q(T14031_Q), .CK(T3075_Y),     .A(T858_Y));
KC_TLAT_X1 T14519 ( .B(T15820_Y), .Q(T14519_Q), .CK(T3217_Y),     .A(T12333_Y));
KC_TLAT_X1 T14953 ( .B(T15820_Y), .Q(T14953_Q), .CK(T5715_Y),     .A(T11959_Y));
KC_TLAT_X1 T14532 ( .B(T15556_Y), .Q(T14532_Q), .CK(T3217_Y),     .A(T6035_Y));
KC_TLAT_X1 T14531 ( .B(T15822_Y), .Q(T14531_Q), .CK(T3215_Y),     .A(T6032_Y));
KC_TLAT_X1 T14524 ( .B(T5757_Y), .Q(T14524_Q), .CK(T3217_Y),     .A(T6058_Y));
KC_TLAT_X1 T14539 ( .B(T5757_Y), .Q(T14539_Q), .CK(T3217_Y),     .A(T11358_Y));
KC_TLAT_X1 T14552 ( .B(T15567_Y), .Q(T14552_Q), .CK(T3279_Y),     .A(T10636_Y));
KC_TLAT_X1 T14563 ( .B(T9227_Y), .Q(T14563_Q), .CK(T3288_Y),     .A(T13055_Y));
KC_TLAT_X1 T14575 ( .B(T15642_Y), .Q(T14575_Q), .CK(T13268_Y),     .A(T3438_Y));
KC_TLAT_X1 T14579 ( .B(T15719_Y), .Q(T14579_Q), .CK(T15192_Y),     .A(T3432_Y));
KC_TLAT_X1 T14580 ( .B(T15719_Y), .Q(T14580_Q), .CK(T15192_Y),     .A(T11683_Y));
KC_TLAT_X1 T13667 ( .B(T15385_Y), .Q(T13667_Q), .CK(T3584_Y),     .A(T12515_Y));
KC_TLAT_X1 T13926 ( .B(T6838_Y), .Q(T13926_Q), .CK(T3075_Y),     .A(T12665_Y));
KC_TLAT_X1 T14353 ( .B(T15516_Y), .Q(T14353_Q), .CK(T16253_Y),     .A(T16252_Y));
KC_TLAT_X1 T14352 ( .B(T15517_Y), .Q(T14352_Q), .CK(T16253_Y),     .A(T16257_Y));
KC_TLAT_X1 T14333 ( .B(T15514_Y), .Q(T14333_Q), .CK(T16253_Y),     .A(T12742_Y));
KC_TLAT_X1 T14331 ( .B(T15516_Y), .Q(T14331_Q), .CK(T16253_Y),     .A(T12741_Y));
KC_TLAT_X1 T14321 ( .B(T15514_Y), .Q(T14321_Q), .CK(T16253_Y),     .A(T1542_Y));
KC_TLAT_X1 T14394 ( .B(T15516_Y), .Q(T14394_Q), .CK(T16253_Y),     .A(T3773_Y));
KC_TLAT_X1 T14393 ( .B(T4870_Y), .Q(T14393_Q), .CK(T16253_Y),     .A(T16246_Y));
KC_TLAT_X1 T14545 ( .B(T15563_Y), .Q(T14545_Q), .CK(T3217_Y),     .A(T3813_Y));
KC_TLAT_X1 T14542 ( .B(T5757_Y), .Q(T14542_Q), .CK(T3215_Y),     .A(T11337_Y));
KC_TLAT_X1 T14556 ( .B(T15564_Y), .Q(T14556_Q), .CK(T5715_Y),     .A(T15878_Y));
KC_TLAT_X1 T14791 ( .B(T15363_Y), .Q(T14791_Q), .CK(T3584_Y),     .A(T6454_Y));
KC_TLAT_X1 T14790 ( .B(T15680_Y), .Q(T14790_Q), .CK(T3584_Y),     .A(T12517_Y));
KC_TLAT_X1 T13519 ( .B(T15363_Y), .Q(T13519_Q), .CK(T3584_Y),     .A(T12522_Y));
KC_TLAT_X1 T13665 ( .B(T15382_Y), .Q(T13665_Q), .CK(T3584_Y),     .A(T6453_Y));
KC_TLAT_X1 T13664 ( .B(T15382_Y), .Q(T13664_Q), .CK(T3584_Y),     .A(T12524_Y));
KC_TLAT_X1 T13663 ( .B(T15363_Y), .Q(T13663_Q), .CK(T3584_Y),     .A(T4214_Y));
KC_TLAT_X1 T13645 ( .B(T15382_Y), .Q(T13645_Q), .CK(T3584_Y),     .A(T12516_Y));
KC_TLAT_X1 T13644 ( .B(T15363_Y), .Q(T13644_Q), .CK(T3584_Y),     .A(T4215_Y));
KC_TLAT_X1 T13634 ( .B(T15382_Y), .Q(T13634_Q), .CK(T1525_Y),     .A(T4212_Y));
KC_TLAT_X1 T13633 ( .B(T15385_Y), .Q(T13633_Q), .CK(T3584_Y),     .A(T12514_Y));
KC_TLAT_X1 T13621 ( .B(T15363_Y), .Q(T13621_Q), .CK(T3584_Y),     .A(T4210_Y));
KC_TLAT_X1 T13620 ( .B(T15680_Y), .Q(T13620_Q), .CK(T3584_Y),     .A(T4216_Y));
KC_TLAT_X1 T13619 ( .B(T15680_Y), .Q(T13619_Q), .CK(T3584_Y),     .A(T6447_Y));
KC_TLAT_X1 T13618 ( .B(T15385_Y), .Q(T13618_Q), .CK(T3584_Y),     .A(T4211_Y));
KC_TLAT_X1 T13617 ( .B(T15680_Y), .Q(T13617_Q), .CK(T3584_Y),     .A(T12523_Y));
KC_TLAT_X1 T14084 ( .B(T15450_Y), .Q(T14084_Q), .CK(T4282_Y),     .A(T4286_Y));
KC_TLAT_X1 T14062 ( .B(T15445_Y), .Q(T14062_Q), .CK(T4282_Y),     .A(T4274_Y));
KC_TLAT_X1 T14036 ( .B(T15445_Y), .Q(T14036_Q), .CK(T4282_Y),     .A(T12655_Y));
KC_TLAT_X1 T14035 ( .B(T15445_Y), .Q(T14035_Q), .CK(T4282_Y),     .A(T4278_Y));
KC_TLAT_X1 T14034 ( .B(T15445_Y), .Q(T14034_Q), .CK(T4282_Y),     .A(T12660_Y));
KC_TLAT_X1 T14033 ( .B(T16173_Y), .Q(T14033_Q), .CK(T4282_Y),     .A(T877_Y));
KC_TLAT_X1 T14026 ( .B(T16173_Y), .Q(T14026_Q), .CK(T4282_Y),     .A(T876_Y));
KC_TLAT_X1 T14025 ( .B(T15448_Y), .Q(T14025_Q), .CK(T4282_Y),     .A(T4280_Y));
KC_TLAT_X1 T14154 ( .B(T16173_Y), .Q(T14154_Q), .CK(T4282_Y),     .A(T12643_Y));
KC_TLAT_X1 T14153 ( .B(T16173_Y), .Q(T14153_Q), .CK(T4282_Y),     .A(T12663_Y));
KC_TLAT_X1 T14347 ( .B(T15513_Y), .Q(T14347_Q), .CK(T16253_Y),     .A(T12754_Y));
KC_TLAT_X1 T14346 ( .B(T15513_Y), .Q(T14346_Q), .CK(T16253_Y),     .A(T12746_Y));
KC_TLAT_X1 T14327 ( .B(T15513_Y), .Q(T14327_Q), .CK(T16253_Y),     .A(T1522_Y));
KC_TLAT_X1 T14406 ( .B(T4870_Y), .Q(T14406_Q), .CK(T16253_Y),     .A(T12753_Y));
KC_TLAT_X1 T14405 ( .B(T4870_Y), .Q(T14405_Q), .CK(T16253_Y),     .A(T12756_Y));
KC_TLAT_X1 T14389 ( .B(T4870_Y), .Q(T14389_Q), .CK(T16253_Y),     .A(T12755_Y));
KC_TLAT_X1 T14555 ( .B(T15573_Y), .Q(T14555_Q), .CK(T5351_Y),     .A(T12805_Y));
KC_TLAT_X1 T14561 ( .B(T5880_Y), .Q(T14561_Q), .CK(T5351_Y),     .A(T12811_Y));
KC_TLAT_X1 T14958 ( .B(T15585_Y), .Q(T14958_Q), .CK(T5351_Y),     .A(T12348_Y));
KC_TLAT_X1 T14569 ( .B(T15593_Y), .Q(T14569_Q), .CK(T5351_Y),     .A(T4520_Y));
KC_TLAT_X1 T14568 ( .B(T15593_Y), .Q(T14568_Q), .CK(T5351_Y),     .A(T12825_Y));
KC_TLAT_X1 T14567 ( .B(T15593_Y), .Q(T14567_Q), .CK(T5351_Y),     .A(T5467_Y));
KC_TLAT_X1 T14962 ( .B(T15635_Y), .Q(T14962_Q), .CK(T15192_Y),     .A(T4729_Y));
KC_TLAT_X1 T14578 ( .B(T15635_Y), .Q(T14578_Q), .CK(T15192_Y),     .A(T11784_Y));
KC_TLAT_X1 T14589 ( .B(T15652_Y), .Q(T14589_Q), .CK(T13288_Y),     .A(T16177_Y));
KC_TLAT_X1 T14666 ( .B(T15394_Y), .Q(T14666_Q), .CK(T5361_Y),     .A(T579_Y));
KC_TLAT_X1 T14637 ( .B(T15418_Y), .Q(T14637_Q), .CK(T5361_Y),     .A(T12584_Y));
KC_TLAT_X1 T14864 ( .B(T15437_Y), .Q(T14864_Q), .CK(T1560_Y),     .A(T16179_Y));
KC_TLAT_X1 T14702 ( .B(T15669_Y), .Q(T14702_Q), .CK(T1963_Y),     .A(T368_Y));
KC_TLAT_X1 T14625 ( .B(T15437_Y), .Q(T14625_Q), .CK(T1560_Y),     .A(T12633_Y));
KC_TLAT_X1 T14767 ( .B(T15668_Y), .Q(T14767_Q), .CK(T1963_Y),     .A(T5217_Y));
KC_TLAT_X1 T14944 ( .B(T15822_Y), .Q(T14944_Q), .CK(T5715_Y),     .A(T6720_Y));
KC_TLAT_X1 T14867 ( .B(T15450_Y), .Q(T14867_Q), .CK(T4282_Y),     .A(T4281_Y));
KC_TLAT_X1 T14866 ( .B(T15450_Y), .Q(T14866_Q), .CK(T4282_Y),     .A(T4285_Y));
KC_TLAT_X1 T14843 ( .B(T15445_Y), .Q(T14843_Q), .CK(T4282_Y),     .A(T4276_Y));
KC_TLAT_X1 T14842 ( .B(T16173_Y), .Q(T14842_Q), .CK(T4282_Y),     .A(T12656_Y));
KC_TLAT_X1 T14775 ( .B(T15680_Y), .Q(T14775_Q), .CK(T3584_Y),     .A(T4213_Y));
KC_TLAT_X1 T14678 ( .B(T15340_Y), .Q(T14678_Q), .CK(T1324_Y),     .A(T12489_Y));
KC_TLAT_X1 T13331 ( .B(T15323_Y), .Q(T13331_Q), .CK(T13288_Y),     .A(T5607_Y));
KC_TLAT_X1 T13497 ( .B(T15361_Y), .Q(T13497_Q), .CK(T1324_Y),     .A(T12480_Y));
KC_TLAT_X1 T13682 ( .B(T15359_Y), .Q(T13682_Q), .CK(T1963_Y),     .A(T12484_Y));
KC_TLAT_X1 T13666 ( .B(T15385_Y), .Q(T13666_Q), .CK(T3584_Y),     .A(T12975_Y));
KC_TLAT_X1 T13630 ( .B(T15669_Y), .Q(T13630_Q), .CK(T1963_Y),     .A(T6444_Y));
KC_TLAT_X1 T14745 ( .B(T588_Y), .Q(T14745_Q), .CK(T5361_Y),     .A(T1451_Y));
KC_TLAT_X1 T13720 ( .B(T15394_Y), .Q(T13720_Q), .CK(T5361_Y),     .A(T12920_Y));
KC_TLAT_X1 T13719 ( .B(T15394_Y), .Q(T13719_Q), .CK(T5361_Y),     .A(T12582_Y));
KC_TLAT_X1 T14664 ( .B(T588_Y), .Q(T14664_Q), .CK(T5361_Y),     .A(T12581_Y));
KC_TLAT_X1 T13927 ( .B(T6838_Y), .Q(T13927_Q), .CK(T3075_Y),     .A(T12669_Y));
KC_TLAT_X1 T13849 ( .B(T15438_Y), .Q(T13849_Q), .CK(T1560_Y),     .A(T12621_Y));
KC_TLAT_X1 T14067 ( .B(T15446_Y), .Q(T14067_Q), .CK(T3075_Y),     .A(T12668_Y));
KC_TLAT_X1 T14061 ( .B(T16058_Y), .Q(T14061_Q), .CK(T4282_Y),     .A(T12662_Y));
KC_TLAT_X1 T14040 ( .B(T16058_Y), .Q(T14040_Q), .CK(T4282_Y),     .A(T4279_Y));
KC_TLAT_X1 T14028 ( .B(T15448_Y), .Q(T14028_Q), .CK(T4282_Y),     .A(T12661_Y));
KC_TLAT_X1 T14010 ( .B(T818_Y), .Q(T14010_Q), .CK(T1560_Y),     .A(T12632_Y));
KC_TLAT_X1 T14009 ( .B(T818_Y), .Q(T14009_Q), .CK(T1560_Y),     .A(T1559_Y));
KC_TLAT_X1 T13950 ( .B(T15437_Y), .Q(T13950_Q), .CK(T1560_Y),     .A(T1556_Y));
KC_TLAT_X1 T13938 ( .B(T849_Y), .Q(T13938_Q), .CK(T1560_Y),     .A(T4892_Y));
KC_TLAT_X1 T13937 ( .B(T16180_Y), .Q(T13937_Q), .CK(T1560_Y),     .A(T12631_Y));
KC_TLAT_X1 T14184 ( .B(T15475_Y), .Q(T14184_Q), .CK(T5423_Y),     .A(T11284_Y));
KC_TLAT_X1 T14138 ( .B(T15465_Y), .Q(T14138_Q), .CK(T15172_Y),     .A(T1090_Y));
KC_TLAT_X1 T14113 ( .B(T15465_Y), .Q(T14113_Q), .CK(T1105_Y),     .A(T1104_Y));
KC_TLAT_X1 T14355 ( .B(T15516_Y), .Q(T14355_Q), .CK(T16253_Y),     .A(T16292_Y));
KC_TLAT_X1 T14354 ( .B(T15516_Y), .Q(T14354_Q), .CK(T16253_Y),     .A(T4326_Y));
KC_TLAT_X1 T14332 ( .B(T15516_Y), .Q(T14332_Q), .CK(T16253_Y),     .A(T12745_Y));
KC_TLAT_X1 T14255 ( .B(T15661_Y), .Q(T14255_Q), .CK(T13261_Y),     .A(T1503_Y));
KC_TLAT_X1 T14237 ( .B(T15661_Y), .Q(T14237_Q), .CK(T13261_Y),     .A(T12725_Y));
KC_TLAT_X1 T14211 ( .B(T15494_Y), .Q(T14211_Q), .CK(T13261_Y),     .A(T12726_Y));
KC_TLAT_X1 T14412 ( .B(T4870_Y), .Q(T14412_Q), .CK(T16253_Y),     .A(T5410_Y));
KC_TLAT_X1 T14392 ( .B(T4870_Y), .Q(T14392_Q), .CK(T16253_Y),     .A(T16247_Y));
KC_TLAT_X1 T14374 ( .B(T15526_Y), .Q(T14374_Q), .CK(T13261_Y),     .A(T12728_Y));
KC_TLAT_X1 T14497 ( .B(T15547_Y), .Q(T14497_Q), .CK(T3217_Y),     .A(T5724_Y));
KC_TLAT_X1 T14452 ( .B(T15541_Y), .Q(T14452_Q), .CK(T991_Y),     .A(T955_Y));
KC_TLAT_X1 T14451 ( .B(T15539_Y), .Q(T14451_Q), .CK(T774_Y),     .A(T9161_Y));
KC_TLAT_X1 T14948 ( .B(T15695_Y), .Q(T14948_Q), .CK(T3217_Y),     .A(T6722_Y));
KC_TLAT_X1 T14538 ( .B(T15708_Y), .Q(T14538_Q), .CK(T2157_Y),     .A(T13143_Y));
KC_TLAT_X1 T14955 ( .B(T15568_Y), .Q(T14955_Q), .CK(T2157_Y),     .A(T13122_Y));
KC_TLAT_X1 T14553 ( .B(T15568_Y), .Q(T14553_Q), .CK(T2157_Y),     .A(T2154_Y));
KC_TLAT_X1 T14562 ( .B(T15948_Y), .Q(T14562_Q), .CK(T5351_Y),     .A(T10950_Y));
KC_TLAT_X1 T14574 ( .B(T15617_Y), .Q(T14574_Q), .CK(T13268_Y),     .A(T2872_Y));
KC_TLAT_X1 T14576 ( .B(T15714_Y), .Q(T14576_Q), .CK(T16134_Y),     .A(T15137_Y));
KC_TLAT_X1 T14963 ( .B(T15715_Y), .Q(T14963_Q), .CK(T13268_Y),     .A(T12067_Y));
KC_TLAT_X1 T14582 ( .B(T15715_Y), .Q(T14582_Q), .CK(T5423_Y),     .A(T8151_Y));
KC_TLAT_X1 T14959 ( .B(T15635_Y), .Q(T14959_Q), .CK(T13268_Y),     .A(T4744_Y));
KC_TLAT_X1 T14703 ( .B(T15359_Y), .Q(T14703_Q), .CK(T1963_Y),     .A(T5219_Y));
KC_TLAT_X1 T14665 ( .B(T588_Y), .Q(T14665_Q), .CK(T5361_Y),     .A(T5273_Y));
KC_DFFHQ_X1 T13337 ( .Q(T13337_Q), .CK(T13345_Q), .D(T15242_Y));
KC_DFFHQ_X1 T13334 ( .Q(T13334_Q), .CK(T13346_Q), .D(T15242_Y));
KC_DFFHQ_X1 T14586 ( .Q(T14586_Q), .CK(T13467_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13438 ( .Q(T13438_Q), .CK(T13345_Q), .D(T15243_Y));
KC_DFFHQ_X1 T13436 ( .Q(T13436_Q), .CK(T13467_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13435 ( .Q(T13435_Q), .CK(T13345_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13433 ( .Q(T13433_Q), .CK(T14678_Q), .D(T15242_Y));
KC_DFFHQ_X1 T13432 ( .Q(T13432_Q), .CK(T13345_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13565 ( .Q(T13565_Q), .CK(T13496_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13386 ( .Q(T13386_Q), .CK(T14678_Q), .D(T15210_Y));
KC_DFFHQ_X1 T13383 ( .Q(T13383_Q), .CK(T13346_Q), .D(T15236_Y));
KC_DFFHQ_X1 T13382 ( .Q(T13382_Q), .CK(T13346_Q), .D(T15210_Y));
KC_DFFHQ_X1 T13369 ( .Q(T13369_Q), .CK(T13346_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13368 ( .Q(T13368_Q), .CK(T13346_Q), .D(T15241_Y));
KC_DFFHQ_X1 T13357 ( .Q(T13357_Q), .CK(T14678_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13354 ( .Q(T13354_Q), .CK(T14678_Q), .D(T15241_Y));
KC_DFFHQ_X1 T13352 ( .Q(T13352_Q), .CK(T13345_Q), .D(T15236_Y));
KC_DFFHQ_X1 T14701 ( .Q(T14701_Q), .CK(T13478_Q), .D(T15243_Y));
KC_DFFHQ_X1 T13486 ( .Q(T13486_Q), .CK(T14693_Q), .D(T15243_Y));
KC_DFFHQ_X1 T13485 ( .Q(T13485_Q), .CK(T13495_Q), .D(T15243_Y));
KC_DFFHQ_X1 T13472 ( .Q(T13472_Q), .CK(T13448_Q), .D(T15241_Y));
KC_DFFHQ_X1 T13469 ( .Q(T13469_Q), .CK(T13495_Q), .D(T15241_Y));
KC_DFFHQ_X1 T13462 ( .Q(T13462_Q), .CK(T14693_Q), .D(T15241_Y));
KC_DFFHQ_X1 T13458 ( .Q(T13458_Q), .CK(T13478_Q), .D(T15241_Y));
KC_DFFHQ_X1 T5753 ( .Q(T5753_Q), .CK(T13448_Q), .D(T15210_Y));
KC_DFFHQ_X1 T1262 ( .Q(T1262_Q), .CK(T13448_Q), .D(T15239_Y));
KC_DFFHQ_X1 T14738 ( .Q(T14738_Q), .CK(T13495_Q), .D(T15238_Y));
KC_DFFHQ_X1 T14736 ( .Q(T14736_Q), .CK(T14693_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13616 ( .Q(T13616_Q), .CK(T14693_Q), .D(T15242_Y));
KC_DFFHQ_X1 T13594 ( .Q(T13594_Q), .CK(T13448_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13593 ( .Q(T13593_Q), .CK(T13495_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13592 ( .Q(T13592_Q), .CK(T14693_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13578 ( .Q(T13578_Q), .CK(T13478_Q), .D(T15242_Y));
KC_DFFHQ_X1 T13567 ( .Q(T13567_Q), .CK(T13478_Q), .D(T15210_Y));
KC_DFFHQ_X1 T6745 ( .Q(T6745_Q), .CK(T14666_Q), .D(T9699_Y));
KC_DFFHQ_X1 T5768 ( .Q(T5768_Q), .CK(T13495_Q), .D(T15210_Y));
KC_DFFHQ_X1 T14755 ( .Q(T14755_Q), .CK(T13719_Q), .D(T9699_Y));
KC_DFFHQ_X1 T14753 ( .Q(T14753_Q), .CK(T14659_Q), .D(T10416_Y));
KC_DFFHQ_X1 T13744 ( .Q(T13744_Q), .CK(T13448_Q), .D(T15242_Y));
KC_DFFHQ_X1 T13743 ( .Q(T13743_Q), .CK(T14693_Q), .D(T15210_Y));
KC_DFFHQ_X1 T13740 ( .Q(T13740_Q), .CK(T13720_Q), .D(T15193_Y));
KC_DFFHQ_X1 T13730 ( .Q(T13730_Q), .CK(T14666_Q), .D(T15206_Y));
KC_DFFHQ_X1 T13729 ( .Q(T13729_Q), .CK(T13720_Q), .D(T10416_Y));
KC_DFFHQ_X1 T13727 ( .Q(T13727_Q), .CK(T13720_Q), .D(T15206_Y));
KC_DFFHQ_X1 T13709 ( .Q(T13709_Q), .CK(T14666_Q), .D(T15193_Y));
KC_DFFHQ_X1 T13708 ( .Q(T13708_Q), .CK(T13719_Q), .D(T15193_Y));
KC_DFFHQ_X1 T13707 ( .Q(T13707_Q), .CK(T13719_Q), .D(T15206_Y));
KC_DFFHQ_X1 T13706 ( .Q(T13706_Q), .CK(T13719_Q), .D(T10416_Y));
KC_DFFHQ_X1 T13702 ( .Q(T13702_Q), .CK(T14666_Q), .D(T10416_Y));
KC_DFFHQ_X1 T6794 ( .Q(T6794_Q), .CK(T14665_Q), .D(T9699_Y));
KC_DFFHQ_X1 T14672 ( .Q(T14672_Q), .CK(T14659_Q), .D(T15193_Y));
KC_DFFHQ_X1 T14670 ( .Q(T14670_Q), .CK(T14659_Q), .D(T15206_Y));
KC_DFFHQ_X1 T14652 ( .Q(T14652_Q), .CK(T14642_Q), .D(T9788_Y));
KC_DFFHQ_X1 T13869 ( .Q(T13869_Q), .CK(T14643_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13868 ( .Q(T13868_Q), .CK(T14642_Q), .D(T9789_Y));
KC_DFFHQ_X1 T13843 ( .Q(T13843_Q), .CK(T14638_Q), .D(T9699_Y));
KC_DFFHQ_X1 T13842 ( .Q(T13842_Q), .CK(T14638_Q), .D(T15206_Y));
KC_DFFHQ_X1 T13840 ( .Q(T13840_Q), .CK(T13720_Q), .D(T9699_Y));
KC_DFFHQ_X1 T13830 ( .Q(T13830_Q), .CK(T14659_Q), .D(T9699_Y));
KC_DFFHQ_X1 T13826 ( .Q(T13826_Q), .CK(T14642_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13797 ( .Q(T13797_Q), .CK(T14643_Q), .D(T9789_Y));
KC_DFFHQ_X1 T14006 ( .Q(T14006_Q), .CK(T14642_Q), .D(T9811_Y));
KC_DFFHQ_X1 T14003 ( .Q(T14003_Q), .CK(T14643_Q), .D(T9811_Y));
KC_DFFHQ_X1 T14681 ( .Q(T14681_Q), .CK(T13497_Q), .D(T10401_Y));
KC_DFFHQ_X1 T14680 ( .Q(T14680_Q), .CK(T13497_Q), .D(T15209_Y));
KC_DFFHQ_X1 T13384 ( .Q(T13384_Q), .CK(T13376_Q), .D(T9608_Y));
KC_DFFHQ_X1 T13381 ( .Q(T13381_Q), .CK(T13347_Q), .D(T15209_Y));
KC_DFFHQ_X1 T13379 ( .Q(T13379_Q), .CK(T13376_Q), .D(T15240_Y));
KC_DFFHQ_X1 T13378 ( .Q(T13378_Q), .CK(T13347_Q), .D(T10401_Y));
KC_DFFHQ_X1 T13367 ( .Q(T13367_Q), .CK(T13376_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13365 ( .Q(T13365_Q), .CK(T13376_Q), .D(T10401_Y));
KC_DFFHQ_X1 T13363 ( .Q(T13363_Q), .CK(T13376_Q), .D(T15209_Y));
KC_DFFHQ_X1 T13355 ( .Q(T13355_Q), .CK(T13347_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13353 ( .Q(T13353_Q), .CK(T13347_Q), .D(T9608_Y));
KC_DFFHQ_X1 T13351 ( .Q(T13351_Q), .CK(T13347_Q), .D(T15240_Y));
KC_DFFHQ_X1 T13350 ( .Q(T13350_Q), .CK(T13497_Q), .D(T15240_Y));
KC_DFFHQ_X1 T14700 ( .Q(T14700_Q), .CK(T13496_Q), .D(T15236_Y));
KC_DFFHQ_X1 T14699 ( .Q(T14699_Q), .CK(T14691_Q), .D(T15240_Y));
KC_DFFHQ_X1 T14698 ( .Q(T14698_Q), .CK(T14691_Q), .D(T10401_Y));
KC_DFFHQ_X1 T13503 ( .Q(T13503_Q), .CK(T13497_Q), .D(T9608_Y));
KC_DFFHQ_X1 T13501 ( .Q(T13501_Q), .CK(T13497_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13500 ( .Q(T13500_Q), .CK(T13608_Q), .D(T10401_Y));
KC_DFFHQ_X1 T13484 ( .Q(T13484_Q), .CK(T14689_Q), .D(T10401_Y));
KC_DFFHQ_X1 T13483 ( .Q(T13483_Q), .CK(T14689_Q), .D(T15240_Y));
KC_DFFHQ_X1 T13471 ( .Q(T13471_Q), .CK(T13448_Q), .D(T15236_Y));
KC_DFFHQ_X1 T13468 ( .Q(T13468_Q), .CK(T13466_Q), .D(T15240_Y));
KC_DFFHQ_X1 T13461 ( .Q(T13461_Q), .CK(T14693_Q), .D(T15236_Y));
KC_DFFHQ_X1 T13460 ( .Q(T13460_Q), .CK(T13495_Q), .D(T15236_Y));
KC_DFFHQ_X1 T13457 ( .Q(T13457_Q), .CK(T13608_Q), .D(T15240_Y));
KC_DFFHQ_X1 T13455 ( .Q(T13455_Q), .CK(T13466_Q), .D(T10401_Y));
KC_DFFHQ_X1 T14737 ( .Q(T14737_Q), .CK(T13608_Q), .D(T9608_Y));
KC_DFFHQ_X1 T14735 ( .Q(T14735_Q), .CK(T14689_Q), .D(T9608_Y));
KC_DFFHQ_X1 T14732 ( .Q(T14732_Q), .CK(T13608_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13615 ( .Q(T13615_Q), .CK(T13466_Q), .D(T15203_Y));
KC_DFFHQ_X1 T13614 ( .Q(T13614_Q), .CK(T13466_Q), .D(T15209_Y));
KC_DFFHQ_X1 T13612 ( .Q(T13612_Q), .CK(T13466_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13590 ( .Q(T13590_Q), .CK(T13608_Q), .D(T15209_Y));
KC_DFFHQ_X1 T13589 ( .Q(T13589_Q), .CK(T14689_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13588 ( .Q(T13588_Q), .CK(T14689_Q), .D(T15209_Y));
KC_DFFHQ_X1 T13577 ( .Q(T13577_Q), .CK(T14689_Q), .D(T15203_Y));
KC_DFFHQ_X1 T14751 ( .Q(T14751_Q), .CK(T14745_Q), .D(T9713_Y));
KC_DFFHQ_X1 T14749 ( .Q(T14749_Q), .CK(T13815_Q), .D(T9713_Y));
KC_DFFHQ_X1 T13741 ( .Q(T13741_Q), .CK(T14690_Q), .D(T15203_Y));
KC_DFFHQ_X1 T13739 ( .Q(T13739_Q), .CK(T14745_Q), .D(T15206_Y));
KC_DFFHQ_X1 T13737 ( .Q(T13737_Q), .CK(T14665_Q), .D(T9713_Y));
KC_DFFHQ_X1 T13728 ( .Q(T13728_Q), .CK(T14664_Q), .D(T15193_Y));
KC_DFFHQ_X1 T13726 ( .Q(T13726_Q), .CK(T14745_Q), .D(T15193_Y));
KC_DFFHQ_X1 T13725 ( .Q(T13725_Q), .CK(T14664_Q), .D(T10416_Y));
KC_DFFHQ_X1 T13724 ( .Q(T13724_Q), .CK(T13720_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13723 ( .Q(T13723_Q), .CK(T13720_Q), .D(T9713_Y));
KC_DFFHQ_X1 T13705 ( .Q(T13705_Q), .CK(T14665_Q), .D(T15193_Y));
KC_DFFHQ_X1 T13704 ( .Q(T13704_Q), .CK(T14745_Q), .D(T10416_Y));
KC_DFFHQ_X1 T13701 ( .Q(T13701_Q), .CK(T13719_Q), .D(T9713_Y));
KC_DFFHQ_X1 T13699 ( .Q(T13699_Q), .CK(T14666_Q), .D(T9713_Y));
KC_DFFHQ_X1 T14671 ( .Q(T14671_Q), .CK(T13815_Q), .D(T15193_Y));
KC_DFFHQ_X1 T14669 ( .Q(T14669_Q), .CK(T14664_Q), .D(T15206_Y));
KC_DFFHQ_X1 T14667 ( .Q(T14667_Q), .CK(T14664_Q), .D(T9713_Y));
KC_DFFHQ_X1 T14651 ( .Q(T14651_Q), .CK(T13858_Q), .D(T9789_Y));
KC_DFFHQ_X1 T14647 ( .Q(T14647_Q), .CK(T13792_Q), .D(T9789_Y));
KC_DFFHQ_X1 T13871 ( .Q(T13871_Q), .CK(T13856_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13867 ( .Q(T13867_Q), .CK(T13793_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13863 ( .Q(T13863_Q), .CK(T13792_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13861 ( .Q(T13861_Q), .CK(T13791_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13860 ( .Q(T13860_Q), .CK(T13857_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13841 ( .Q(T13841_Q), .CK(T13815_Q), .D(T15206_Y));
KC_DFFHQ_X1 T13839 ( .Q(T13839_Q), .CK(T14638_Q), .D(T9713_Y));
KC_DFFHQ_X1 T13829 ( .Q(T13829_Q), .CK(T14664_Q), .D(T9699_Y));
KC_DFFHQ_X1 T13828 ( .Q(T13828_Q), .CK(T13815_Q), .D(T9699_Y));
KC_DFFHQ_X1 T13827 ( .Q(T13827_Q), .CK(T13858_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13825 ( .Q(T13825_Q), .CK(T14659_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13823 ( .Q(T13823_Q), .CK(T14638_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13821 ( .Q(T13821_Q), .CK(T14659_Q), .D(T9713_Y));
KC_DFFHQ_X1 T13796 ( .Q(T13796_Q), .CK(T13793_Q), .D(T9789_Y));
KC_DFFHQ_X1 T13795 ( .Q(T13795_Q), .CK(T13856_Q), .D(T9789_Y));
KC_DFFHQ_X1 T14023 ( .Q(T14023_Q), .CK(T13858_Q), .D(T9812_Y));
KC_DFFHQ_X1 T14022 ( .Q(T14022_Q), .CK(T13858_Q), .D(T9811_Y));
KC_DFFHQ_X1 T14021 ( .Q(T14021_Q), .CK(T13857_Q), .D(T9811_Y));
KC_DFFHQ_X1 T14020 ( .Q(T14020_Q), .CK(T13791_Q), .D(T9811_Y));
KC_DFFHQ_X1 T14018 ( .Q(T14018_Q), .CK(T13792_Q), .D(T9811_Y));
KC_DFFHQ_X1 T14005 ( .Q(T14005_Q), .CK(T13856_Q), .D(T9788_Y));
KC_DFFHQ_X1 T14000 ( .Q(T14000_Q), .CK(T13793_Q), .D(T9788_Y));
KC_DFFHQ_X1 T13983 ( .Q(T13983_Q), .CK(T13856_Q), .D(T9811_Y));
KC_DFFHQ_X1 T13971 ( .Q(T13971_Q), .CK(T13793_Q), .D(T9811_Y));
KC_DFFHQ_X1 T13968 ( .Q(T13968_Q), .CK(T13791_Q), .D(T9788_Y));
KC_DFFHQ_X1 T13967 ( .Q(T13967_Q), .CK(T13857_Q), .D(T9788_Y));
KC_DFFHQ_X1 T13964 ( .Q(T13964_Q), .CK(T13791_Q), .D(T9789_Y));
KC_DFFHQ_X1 T13963 ( .Q(T13963_Q), .CK(T13857_Q), .D(T9789_Y));
KC_DFFHQ_X1 T13948 ( .Q(T13948_Q), .CK(T13857_Q), .D(T9812_Y));
KC_DFFHQ_X1 T14133 ( .Q(T14133_Q), .CK(T14255_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14111 ( .Q(T14111_Q), .CK(T14252_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14262 ( .Q(T14262_Q), .CK(T14255_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14261 ( .Q(T14261_Q), .CK(T14255_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14679 ( .Q(T14679_Q), .CK(T13497_Q), .D(T15208_Y));
KC_DFFHQ_X1 T13380 ( .Q(T13380_Q), .CK(T13376_Q), .D(T15208_Y));
KC_DFFHQ_X1 T13377 ( .Q(T13377_Q), .CK(T13376_Q), .D(T10394_Y));
KC_DFFHQ_X1 T13364 ( .Q(T13364_Q), .CK(T13347_Q), .D(T15208_Y));
KC_DFFHQ_X1 T13362 ( .Q(T13362_Q), .CK(T13347_Q), .D(T10394_Y));
KC_DFFHQ_X1 T13349 ( .Q(T13349_Q), .CK(T14678_Q), .D(T10402_Y));
KC_DFFHQ_X1 T13348 ( .Q(T13348_Q), .CK(T13346_Q), .D(T10402_Y));
KC_DFFHQ_X1 T14696 ( .Q(T14696_Q), .CK(T14690_Q), .D(T10394_Y));
KC_DFFHQ_X1 T14695 ( .Q(T14695_Q), .CK(T14691_Q), .D(T10394_Y));
KC_DFFHQ_X1 T14694 ( .Q(T14694_Q), .CK(T13466_Q), .D(T15208_Y));
KC_DFFHQ_X1 T13499 ( .Q(T13499_Q), .CK(T13345_Q), .D(T10402_Y));
KC_DFFHQ_X1 T13498 ( .Q(T13498_Q), .CK(T13497_Q), .D(T10394_Y));
KC_DFFHQ_X1 T13456 ( .Q(T13456_Q), .CK(T14693_Q), .D(T10402_Y));
KC_DFFHQ_X1 T13454 ( .Q(T13454_Q), .CK(T13467_Q), .D(T10402_Y));
KC_DFFHQ_X1 T13453 ( .Q(T13453_Q), .CK(T13495_Q), .D(T10402_Y));
KC_DFFHQ_X1 T13451 ( .Q(T13451_Q), .CK(T13496_Q), .D(T10402_Y));
KC_DFFHQ_X1 T13450 ( .Q(T13450_Q), .CK(T13478_Q), .D(T10402_Y));
KC_DFFHQ_X1 T13449 ( .Q(T13449_Q), .CK(T13448_Q), .D(T10402_Y));
KC_DFFHQ_X1 T14734 ( .Q(T14734_Q), .CK(T14690_Q), .D(T15209_Y));
KC_DFFHQ_X1 T13611 ( .Q(T13611_Q), .CK(T14688_Q), .D(T15240_Y));
KC_DFFHQ_X1 T13610 ( .Q(T13610_Q), .CK(T14691_Q), .D(T15208_Y));
KC_DFFHQ_X1 T13597 ( .Q(T13597_Q), .CK(T1651_Y), .D(T12509_Y));
KC_DFFHQ_X1 T13587 ( .Q(T13587_Q), .CK(T14688_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13575 ( .Q(T13575_Q), .CK(T1651_Y), .D(T12498_Y));
KC_DFFHQ_X1 T14750 ( .Q(T14750_Q), .CK(T14745_Q), .D(T9698_Y));
KC_DFFHQ_X1 T14748 ( .Q(T14748_Q), .CK(T14665_Q), .D(T9698_Y));
KC_DFFHQ_X1 T14747 ( .Q(T14747_Q), .CK(T14745_Q), .D(T9700_Y));
KC_DFFHQ_X1 T14746 ( .Q(T14746_Q), .CK(T14665_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13722 ( .Q(T13722_Q), .CK(T14666_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13721 ( .Q(T13721_Q), .CK(T13720_Q), .D(T9698_Y));
KC_DFFHQ_X1 T13697 ( .Q(T13697_Q), .CK(T13719_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13696 ( .Q(T13696_Q), .CK(T14666_Q), .D(T9698_Y));
KC_DFFHQ_X1 T13695 ( .Q(T13695_Q), .CK(T13720_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13694 ( .Q(T13694_Q), .CK(T13719_Q), .D(T9698_Y));
KC_DFFHQ_X1 T14641 ( .Q(T14641_Q), .CK(T14643_Q), .D(T9792_Y));
KC_DFFHQ_X1 T13865 ( .Q(T13865_Q), .CK(T13791_Q), .D(T9793_Y));
KC_DFFHQ_X1 T13859 ( .Q(T13859_Q), .CK(T13857_Q), .D(T9793_Y));
KC_DFFHQ_X1 T13837 ( .Q(T13837_Q), .CK(T14664_Q), .D(T9698_Y));
KC_DFFHQ_X1 T13836 ( .Q(T13836_Q), .CK(T14664_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13820 ( .Q(T13820_Q), .CK(T14659_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13819 ( .Q(T13819_Q), .CK(T13815_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13818 ( .Q(T13818_Q), .CK(T13815_Q), .D(T9698_Y));
KC_DFFHQ_X1 T13817 ( .Q(T13817_Q), .CK(T14638_Q), .D(T9700_Y));
KC_DFFHQ_X1 T13816 ( .Q(T13816_Q), .CK(T14638_Q), .D(T9698_Y));
KC_DFFHQ_X1 T14024 ( .Q(T14024_Q), .CK(T13858_Q), .D(T9696_Y));
KC_DFFHQ_X1 T14017 ( .Q(T14017_Q), .CK(T13791_Q), .D(T9792_Y));
KC_DFFHQ_X1 T14016 ( .Q(T14016_Q), .CK(T13858_Q), .D(T9792_Y));
KC_DFFHQ_X1 T14015 ( .Q(T14015_Q), .CK(T13857_Q), .D(T9792_Y));
KC_DFFHQ_X1 T14014 ( .Q(T14014_Q), .CK(T13857_Q), .D(T9696_Y));
KC_DFFHQ_X1 T14001 ( .Q(T14001_Q), .CK(T14637_Q), .D(T9696_Y));
KC_DFFHQ_X1 T13999 ( .Q(T13999_Q), .CK(T14642_Q), .D(T9792_Y));
KC_DFFHQ_X1 T13998 ( .Q(T13998_Q), .CK(T14643_Q), .D(T9696_Y));
KC_DFFHQ_X1 T13997 ( .Q(T13997_Q), .CK(T14637_Q), .D(T9792_Y));
KC_DFFHQ_X1 T13969 ( .Q(T13969_Q), .CK(T13793_Q), .D(T9696_Y));
KC_DFFHQ_X1 T13966 ( .Q(T13966_Q), .CK(T13856_Q), .D(T9696_Y));
KC_DFFHQ_X1 T13962 ( .Q(T13962_Q), .CK(T13856_Q), .D(T9792_Y));
KC_DFFHQ_X1 T13961 ( .Q(T13961_Q), .CK(T13793_Q), .D(T9792_Y));
KC_DFFHQ_X1 T13947 ( .Q(T13947_Q), .CK(T13791_Q), .D(T9696_Y));
KC_DFFHQ_X1 T13946 ( .Q(T13946_Q), .CK(T1549_Y), .D(T12638_Y));
KC_DFFHQ_X1 T13945 ( .Q(T13945_Q), .CK(T13792_Q), .D(T9792_Y));
KC_DFFHQ_X1 T13944 ( .Q(T13944_Q), .CK(T13792_Q), .D(T9696_Y));
KC_DFFHQ_X1 T14619 ( .Q(T14619_Q), .CK(T14224_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14618 ( .Q(T14618_Q), .CK(T14237_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14617 ( .Q(T14617_Q), .CK(T14250_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14605 ( .Q(T14605_Q), .CK(T14252_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14603 ( .Q(T14603_Q), .CK(T14237_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14135 ( .Q(T14135_Q), .CK(T14276_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14132 ( .Q(T14132_Q), .CK(T14224_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14131 ( .Q(T14131_Q), .CK(T14237_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14130 ( .Q(T14130_Q), .CK(T14250_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14122 ( .Q(T14122_Q), .CK(T14211_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14120 ( .Q(T14120_Q), .CK(T14224_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14118 ( .Q(T14118_Q), .CK(T14237_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14112 ( .Q(T14112_Q), .CK(T14252_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14110 ( .Q(T14110_Q), .CK(T14211_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14109 ( .Q(T14109_Q), .CK(T14209_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14108 ( .Q(T14108_Q), .CK(T14250_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14106 ( .Q(T14106_Q), .CK(T14276_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14282 ( .Q(T14282_Q), .CK(T14211_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14281 ( .Q(T14281_Q), .CK(T14255_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14279 ( .Q(T14279_Q), .CK(T14224_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14278 ( .Q(T14278_Q), .CK(T14250_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14277 ( .Q(T14277_Q), .CK(T14212_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14259 ( .Q(T14259_Q), .CK(T14237_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14258 ( .Q(T14258_Q), .CK(T14211_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14257 ( .Q(T14257_Q), .CK(T14250_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14256 ( .Q(T14256_Q), .CK(T14252_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14240 ( .Q(T14240_Q), .CK(T14209_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14239 ( .Q(T14239_Q), .CK(T14250_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14238 ( .Q(T14238_Q), .CK(T14237_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14230 ( .Q(T14230_Q), .CK(T14252_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14229 ( .Q(T14229_Q), .CK(T14276_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14228 ( .Q(T14228_Q), .CK(T14224_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14214 ( .Q(T14214_Q), .CK(T14224_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14213 ( .Q(T14213_Q), .CK(T14209_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14387 ( .Q(T14387_Q), .CK(T14209_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14386 ( .Q(T14386_Q), .CK(T14211_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14382 ( .Q(T14382_Q), .CK(T14212_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14381 ( .Q(T14381_Q), .CK(T14209_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14375 ( .Q(T14375_Q), .CK(T14212_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14692 ( .Q(T14692_Q), .CK(T14688_Q), .D(T10394_Y));
KC_DFFHQ_X1 T13481 ( .Q(T13481_Q), .CK(T13608_Q), .D(T10394_Y));
KC_DFFHQ_X1 T14728 ( .Q(T14728_Q), .CK(T1651_Y), .D(T12909_Y));
KC_DFFHQ_X1 T13607 ( .Q(T13607_Q), .CK(T1651_Y), .D(T12512_Y));
KC_DFFHQ_X1 T13606 ( .Q(T13606_Q), .CK(T1651_Y), .D(T12510_Y));
KC_DFFHQ_X1 T13585 ( .Q(T13585_Q), .CK(T1651_Y), .D(T12507_Y));
KC_DFFHQ_X1 T13584 ( .Q(T13584_Q), .CK(T1651_Y), .D(T12508_Y));
KC_DFFHQ_X1 T13583 ( .Q(T13583_Q), .CK(T1651_Y), .D(T12504_Y));
KC_DFFHQ_X1 T14744 ( .Q(T14744_Q), .CK(T13804_Q), .D(T10351_Y));
KC_DFFHQ_X1 T14743 ( .Q(T14743_Q), .CK(T13849_Q), .D(T10351_Y));
KC_DFFHQ_X1 T14741 ( .Q(T14741_Q), .CK(T13804_Q), .D(T9618_Y));
KC_DFFHQ_X1 T13736 ( .Q(T13736_Q), .CK(T13938_Q), .D(T10351_Y));
KC_DFFHQ_X1 T13718 ( .Q(T13718_Q), .CK(T14009_Q), .D(T9618_Y));
KC_DFFHQ_X1 T13717 ( .Q(T13717_Q), .CK(T1650_Y), .D(T12919_Y));
KC_DFFHQ_X1 T13716 ( .Q(T13716_Q), .CK(T1650_Y), .D(T12536_Y));
KC_DFFHQ_X1 T13693 ( .Q(T13693_Q), .CK(T14009_Q), .D(T10351_Y));
KC_DFFHQ_X1 T13692 ( .Q(T13692_Q), .CK(T1650_Y), .D(T12542_Y));
KC_DFFHQ_X1 T13691 ( .Q(T13691_Q), .CK(T1650_Y), .D(T12541_Y));
KC_DFFHQ_X1 T14661 ( .Q(T14661_Q), .CK(T1650_Y), .D(T12921_Y));
KC_DFFHQ_X1 T14660 ( .Q(T14660_Q), .CK(T13957_Q), .D(T10351_Y));
KC_DFFHQ_X1 T14636 ( .Q(T14636_Q), .CK(T14010_Q), .D(T10348_Y));
KC_DFFHQ_X1 T14635 ( .Q(T14635_Q), .CK(T13957_Q), .D(T10348_Y));
KC_DFFHQ_X1 T13855 ( .Q(T13855_Q), .CK(T14010_Q), .D(T9617_Y));
KC_DFFHQ_X1 T13854 ( .Q(T13854_Q), .CK(T14012_Q), .D(T9618_Y));
KC_DFFHQ_X1 T13835 ( .Q(T13835_Q), .CK(T1650_Y), .D(T12906_Y));
KC_DFFHQ_X1 T13834 ( .Q(T13834_Q), .CK(T13957_Q), .D(T9617_Y));
KC_DFFHQ_X1 T13814 ( .Q(T13814_Q), .CK(T13957_Q), .D(T9618_Y));
KC_DFFHQ_X1 T13813 ( .Q(T13813_Q), .CK(T14012_Q), .D(T10351_Y));
KC_DFFHQ_X1 T13812 ( .Q(T13812_Q), .CK(T1650_Y), .D(T12578_Y));
KC_DFFHQ_X1 T13811 ( .Q(T13811_Q), .CK(T14012_Q), .D(T9617_Y));
KC_DFFHQ_X1 T13810 ( .Q(T13810_Q), .CK(T14010_Q), .D(T10351_Y));
KC_DFFHQ_X1 T13790 ( .Q(T13790_Q), .CK(T14010_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13789 ( .Q(T13789_Q), .CK(T14010_Q), .D(T9618_Y));
KC_DFFHQ_X1 T14013 ( .Q(T14013_Q), .CK(T1549_Y), .D(T12637_Y));
KC_DFFHQ_X1 T13996 ( .Q(T13996_Q), .CK(T13849_Q), .D(T10348_Y));
KC_DFFHQ_X1 T13995 ( .Q(T13995_Q), .CK(T14012_Q), .D(T10350_Y));
KC_DFFHQ_X1 T13994 ( .Q(T13994_Q), .CK(T13957_Q), .D(T10350_Y));
KC_DFFHQ_X1 T13981 ( .Q(T13981_Q), .CK(T14010_Q), .D(T10350_Y));
KC_DFFHQ_X1 T13980 ( .Q(T13980_Q), .CK(T14010_Q), .D(T10409_Y));
KC_DFFHQ_X1 T13979 ( .Q(T13979_Q), .CK(T14012_Q), .D(T10409_Y));
KC_DFFHQ_X1 T13978 ( .Q(T13978_Q), .CK(T1549_Y), .D(T12622_Y));
KC_DFFHQ_X1 T13960 ( .Q(T13960_Q), .CK(T1549_Y), .D(T12623_Y));
KC_DFFHQ_X1 T13959 ( .Q(T13959_Q), .CK(T1549_Y), .D(T12636_Y));
KC_DFFHQ_X1 T13958 ( .Q(T13958_Q), .CK(T1549_Y), .D(T12634_Y));
KC_DFFHQ_X1 T13943 ( .Q(T13943_Q), .CK(T1549_Y), .D(T12618_Y));
KC_DFFHQ_X1 T13942 ( .Q(T13942_Q), .CK(T4900_Y), .D(T12893_Y));
KC_DFFHQ_X1 T13941 ( .Q(T13941_Q), .CK(T1549_Y), .D(T12895_Y));
KC_DFFHQ_X1 T14614 ( .Q(T14614_Q), .CK(T1549_Y), .D(T12699_Y));
KC_DFFHQ_X1 T14613 ( .Q(T14613_Q), .CK(T1549_Y), .D(T13026_Y));
KC_DFFHQ_X1 T14602 ( .Q(T14602_Q), .CK(T14253_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14601 ( .Q(T14601_Q), .CK(T14253_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14129 ( .Q(T14129_Q), .CK(T4900_Y), .D(T12694_Y));
KC_DFFHQ_X1 T14128 ( .Q(T14128_Q), .CK(T1549_Y), .D(T12700_Y));
KC_DFFHQ_X1 T14127 ( .Q(T14127_Q), .CK(T1549_Y), .D(T12702_Y));
KC_DFFHQ_X1 T14126 ( .Q(T14126_Q), .CK(T1549_Y), .D(T12701_Y));
KC_DFFHQ_X1 T14117 ( .Q(T14117_Q), .CK(T14270_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14116 ( .Q(T14116_Q), .CK(T14270_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14115 ( .Q(T14115_Q), .CK(T14224_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14105 ( .Q(T14105_Q), .CK(T14210_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14104 ( .Q(T14104_Q), .CK(T14210_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14103 ( .Q(T14103_Q), .CK(T14251_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14102 ( .Q(T14102_Q), .CK(T14251_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14099 ( .Q(T14099_Q), .CK(T14270_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14275 ( .Q(T14275_Q), .CK(T14236_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14273 ( .Q(T14273_Q), .CK(T14209_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14272 ( .Q(T14272_Q), .CK(T14225_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14271 ( .Q(T14271_Q), .CK(T14211_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14265 ( .Q(T14265_Q), .CK(T14225_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14235 ( .Q(T14235_Q), .CK(T14236_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14226 ( .Q(T14226_Q), .CK(T14225_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14223 ( .Q(T14223_Q), .CK(T14253_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14208 ( .Q(T14208_Q), .CK(T14210_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14385 ( .Q(T14385_Q), .CK(T14374_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14380 ( .Q(T14380_Q), .CK(T14374_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14379 ( .Q(T14379_Q), .CK(T14591_Q), .D(T9905_Y));
KC_DFFHQ_X1 T14373 ( .Q(T14373_Q), .CK(T13329_Q), .D(T9905_Y));
KC_DFFHQ_X1 T13375 ( .Q(T13375_Q), .CK(T14702_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13374 ( .Q(T13374_Q), .CK(T13445_Q), .D(T15249_Y));
KC_DFFHQ_X1 T13370 ( .Q(T13370_Q), .CK(T13745_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13344 ( .Q(T13344_Q), .CK(T14683_Q), .D(T15249_Y));
KC_DFFHQ_X1 T13343 ( .Q(T13343_Q), .CK(T13491_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13342 ( .Q(T13342_Q), .CK(T13492_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13341 ( .Q(T13341_Q), .CK(T13745_Q), .D(T15249_Y));
KC_DFFHQ_X1 T14687 ( .Q(T14687_Q), .CK(T14683_Q), .D(T10444_Y));
KC_DFFHQ_X1 T14686 ( .Q(T14686_Q), .CK(T13464_Q), .D(T10444_Y));
KC_DFFHQ_X1 T14685 ( .Q(T14685_Q), .CK(T13490_Q), .D(T10444_Y));
KC_DFFHQ_X1 T13494 ( .Q(T13494_Q), .CK(T14682_Q), .D(T15249_Y));
KC_DFFHQ_X1 T13493 ( .Q(T13493_Q), .CK(T13340_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13487 ( .Q(T13487_Q), .CK(T13490_Q), .D(T15249_Y));
KC_DFFHQ_X1 T13480 ( .Q(T13480_Q), .CK(T13630_Q), .D(T10444_Y));
KC_DFFHQ_X1 T13479 ( .Q(T13479_Q), .CK(T14682_Q), .D(T10444_Y));
KC_DFFHQ_X1 T13473 ( .Q(T13473_Q), .CK(T13682_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13465 ( .Q(T13465_Q), .CK(T13630_Q), .D(T15249_Y));
KC_DFFHQ_X1 T13463 ( .Q(T13463_Q), .CK(T14703_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13447 ( .Q(T13447_Q), .CK(T13464_Q), .D(T15249_Y));
KC_DFFHQ_X1 T13444 ( .Q(T13444_Q), .CK(T13446_Q), .D(T15249_Y));
KC_DFFHQ_X1 T14724 ( .Q(T14724_Q), .CK(T13491_Q), .D(T9687_Y));
KC_DFFHQ_X1 T14723 ( .Q(T14723_Q), .CK(T14702_Q), .D(T9606_Y));
KC_DFFHQ_X1 T13605 ( .Q(T13605_Q), .CK(T13745_Q), .D(T10445_Y));
KC_DFFHQ_X1 T13604 ( .Q(T13604_Q), .CK(T13445_Q), .D(T10445_Y));
KC_DFFHQ_X1 T13598 ( .Q(T13598_Q), .CK(T13682_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13596 ( .Q(T13596_Q), .CK(T13491_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13582 ( .Q(T13582_Q), .CK(T14702_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13580 ( .Q(T13580_Q), .CK(T13492_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13574 ( .Q(T13574_Q), .CK(T14702_Q), .D(T9687_Y));
KC_DFFHQ_X1 T14742 ( .Q(T14742_Q), .CK(T13938_Q), .D(T9609_Y));
KC_DFFHQ_X1 T14740 ( .Q(T14740_Q), .CK(T13938_Q), .D(T9617_Y));
KC_DFFHQ_X1 T13735 ( .Q(T13735_Q), .CK(T13939_Q), .D(T9609_Y));
KC_DFFHQ_X1 T13734 ( .Q(T13734_Q), .CK(T13940_Q), .D(T9617_Y));
KC_DFFHQ_X1 T13733 ( .Q(T13733_Q), .CK(T13940_Q), .D(T9618_Y));
KC_DFFHQ_X1 T13731 ( .Q(T13731_Q), .CK(T13940_Q), .D(T9609_Y));
KC_DFFHQ_X1 T13714 ( .Q(T13714_Q), .CK(T13939_Q), .D(T9617_Y));
KC_DFFHQ_X1 T13713 ( .Q(T13713_Q), .CK(T14009_Q), .D(T9617_Y));
KC_DFFHQ_X1 T13710 ( .Q(T13710_Q), .CK(T1638_Y), .D(T12544_Y));
KC_DFFHQ_X1 T13690 ( .Q(T13690_Q), .CK(T13940_Q), .D(T10351_Y));
KC_DFFHQ_X1 T13689 ( .Q(T13689_Q), .CK(T13492_Q), .D(T9606_Y));
KC_DFFHQ_X1 T13686 ( .Q(T13686_Q), .CK(T13340_Q), .D(T9687_Y));
KC_DFFHQ_X1 T14658 ( .Q(T14658_Q), .CK(T13804_Q), .D(T9617_Y));
KC_DFFHQ_X1 T14629 ( .Q(T14629_Q), .CK(T14008_Q), .D(T8533_Y));
KC_DFFHQ_X1 T13853 ( .Q(T13853_Q), .CK(T13804_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13852 ( .Q(T13852_Q), .CK(T14012_Q), .D(T9609_Y));
KC_DFFHQ_X1 T13851 ( .Q(T13851_Q), .CK(T13804_Q), .D(T10409_Y));
KC_DFFHQ_X1 T13850 ( .Q(T13850_Q), .CK(T13940_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13846 ( .Q(T13846_Q), .CK(T14625_Q), .D(T8533_Y));
KC_DFFHQ_X1 T13833 ( .Q(T13833_Q), .CK(T13804_Q), .D(T9609_Y));
KC_DFFHQ_X1 T13809 ( .Q(T13809_Q), .CK(T13849_Q), .D(T9609_Y));
KC_DFFHQ_X1 T13808 ( .Q(T13808_Q), .CK(T14009_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13805 ( .Q(T13805_Q), .CK(T13957_Q), .D(T9609_Y));
KC_DFFHQ_X1 T13803 ( .Q(T13803_Q), .CK(T13939_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13799 ( .Q(T13799_Q), .CK(T14625_Q), .D(T6716_Y));
KC_DFFHQ_X1 T13787 ( .Q(T13787_Q), .CK(T13938_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13786 ( .Q(T13786_Q), .CK(T14010_Q), .D(T9609_Y));
KC_DFFHQ_X1 T13785 ( .Q(T13785_Q), .CK(T13849_Q), .D(T10409_Y));
KC_DFFHQ_X1 T13784 ( .Q(T13784_Q), .CK(T13952_Q), .D(T8533_Y));
KC_DFFHQ_X1 T16178 ( .Q(T16178_Q), .CK(T13938_Q), .D(T10409_Y));
KC_DFFHQ_X1 T9784 ( .Q(T9784_Q), .CK(T14009_Q), .D(T10348_Y));
KC_DFFHQ_X1 T15049 ( .Q(T15049_Q), .CK(T13940_Q), .D(T10348_Y));
KC_DFFHQ_X1 T14011 ( .Q(T14011_Q), .CK(T13939_Q), .D(T10409_Y));
KC_DFFHQ_X1 T13993 ( .Q(T13993_Q), .CK(T13940_Q), .D(T10350_Y));
KC_DFFHQ_X1 T13991 ( .Q(T13991_Q), .CK(T13938_Q), .D(T10350_Y));
KC_DFFHQ_X1 T13987 ( .Q(T13987_Q), .CK(T14625_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13977 ( .Q(T13977_Q), .CK(T13938_Q), .D(T10348_Y));
KC_DFFHQ_X1 T13976 ( .Q(T13976_Q), .CK(T13804_Q), .D(T10348_Y));
KC_DFFHQ_X1 T13975 ( .Q(T13975_Q), .CK(T13939_Q), .D(T10348_Y));
KC_DFFHQ_X1 T13974 ( .Q(T13974_Q), .CK(T13939_Q), .D(T10350_Y));
KC_DFFHQ_X1 T13955 ( .Q(T13955_Q), .CK(T13940_Q), .D(T10409_Y));
KC_DFFHQ_X1 T13954 ( .Q(T13954_Q), .CK(T14009_Q), .D(T10409_Y));
KC_DFFHQ_X1 T14611 ( .Q(T14611_Q), .CK(T4900_Y), .D(T12692_Y));
KC_DFFHQ_X1 T14610 ( .Q(T14610_Q), .CK(T4900_Y), .D(T12892_Y));
KC_DFFHQ_X1 T14609 ( .Q(T14609_Q), .CK(T4900_Y), .D(T12696_Y));
KC_DFFHQ_X1 T14600 ( .Q(T14600_Q), .CK(T14253_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14125 ( .Q(T14125_Q), .CK(T4900_Y), .D(T12697_Y));
KC_DFFHQ_X1 T14124 ( .Q(T14124_Q), .CK(T4900_Y), .D(T12693_Y));
KC_DFFHQ_X1 T14100 ( .Q(T14100_Q), .CK(T14251_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14098 ( .Q(T14098_Q), .CK(T14210_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14269 ( .Q(T14269_Q), .CK(T14253_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14268 ( .Q(T14268_Q), .CK(T14210_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14267 ( .Q(T14267_Q), .CK(T14270_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14248 ( .Q(T14248_Q), .CK(T14270_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14247 ( .Q(T14247_Q), .CK(T14251_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14246 ( .Q(T14246_Q), .CK(T14225_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14245 ( .Q(T14245_Q), .CK(T14270_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14243 ( .Q(T14243_Q), .CK(T14225_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14234 ( .Q(T14234_Q), .CK(T14253_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14233 ( .Q(T14233_Q), .CK(T14270_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14222 ( .Q(T14222_Q), .CK(T14253_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14221 ( .Q(T14221_Q), .CK(T14251_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14220 ( .Q(T14220_Q), .CK(T14251_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14217 ( .Q(T14217_Q), .CK(T14225_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14207 ( .Q(T14207_Q), .CK(T14210_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14206 ( .Q(T14206_Q), .CK(T14210_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14204 ( .Q(T14204_Q), .CK(T14225_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14384 ( .Q(T14384_Q), .CK(T14374_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14378 ( .Q(T14378_Q), .CK(T14374_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14377 ( .Q(T14377_Q), .CK(T14374_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14372 ( .Q(T14372_Q), .CK(T14374_Q), .D(T15225_Y));
KC_DFFHQ_X1 T13328 ( .Q(T13328_Q), .CK(T14591_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14458 ( .Q(T14458_Q), .CK(T14591_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14457 ( .Q(T14457_Q), .CK(T13329_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14456 ( .Q(T14456_Q), .CK(T14591_Q), .D(T9906_Y));
KC_DFFHQ_X1 T15045 ( .Q(T15045_Q), .CK(T13491_Q), .D(T10453_Y));
KC_DFFHQ_X1 T14819 ( .Q(T14819_Q), .CK(T14677_Q), .D(T10453_Y));
KC_DFFHQ_X1 T14676 ( .Q(T14676_Q), .CK(T13492_Q), .D(T10443_Y));
KC_DFFHQ_X1 T13431 ( .Q(T13431_Q), .CK(T13492_Q), .D(T10453_Y));
KC_DFFHQ_X1 T13416 ( .Q(T13416_Q), .CK(T14702_Q), .D(T10453_Y));
KC_DFFHQ_X1 T13372 ( .Q(T13372_Q), .CK(T13491_Q), .D(T10443_Y));
KC_DFFHQ_X1 T13371 ( .Q(T13371_Q), .CK(T14683_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13360 ( .Q(T13360_Q), .CK(T13745_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13359 ( .Q(T13359_Q), .CK(T14702_Q), .D(T10443_Y));
KC_DFFHQ_X1 T14809 ( .Q(T14809_Q), .CK(T13464_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13563 ( .Q(T13563_Q), .CK(T14767_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13537 ( .Q(T13537_Q), .CK(T13464_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13518 ( .Q(T13518_Q), .CK(T13490_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13489 ( .Q(T13489_Q), .CK(T13490_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13488 ( .Q(T13488_Q), .CK(T14682_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13477 ( .Q(T13477_Q), .CK(T13630_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13476 ( .Q(T13476_Q), .CK(T13642_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13475 ( .Q(T13475_Q), .CK(T13446_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13443 ( .Q(T13443_Q), .CK(T14767_Q), .D(T15250_Y));
KC_DFFHQ_X1 T14774 ( .Q(T14774_Q), .CK(T13642_Q), .D(T9687_Y));
KC_DFFHQ_X1 T14719 ( .Q(T14719_Q), .CK(T14703_Q), .D(T9606_Y));
KC_DFFHQ_X1 T13684 ( .Q(T13684_Q), .CK(T13446_Q), .D(T10445_Y));
KC_DFFHQ_X1 T13683 ( .Q(T13683_Q), .CK(T13490_Q), .D(T10445_Y));
KC_DFFHQ_X1 T13662 ( .Q(T13662_Q), .CK(T13757_Q), .D(T9687_Y));
KC_DFFHQ_X1 T13632 ( .Q(T13632_Q), .CK(T14767_Q), .D(T10445_Y));
KC_DFFHQ_X1 T13601 ( .Q(T13601_Q), .CK(T13446_Q), .D(T10444_Y));
KC_DFFHQ_X1 T13600 ( .Q(T13600_Q), .CK(T14677_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13599 ( .Q(T13599_Q), .CK(T14767_Q), .D(T10444_Y));
KC_DFFHQ_X1 T13581 ( .Q(T13581_Q), .CK(T13642_Q), .D(T9606_Y));
KC_DFFHQ_X1 T13572 ( .Q(T13572_Q), .CK(T13757_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13570 ( .Q(T13570_Q), .CK(T13642_Q), .D(T9605_Y));
KC_DFFHQ_X1 T6594 ( .Q(T6594_Q), .CK(T1638_Y), .D(T11921_Y));
KC_DFFHQ_X1 T14941 ( .Q(T14941_Q), .CK(T1638_Y), .D(T11956_Y));
KC_DFFHQ_X1 T14739 ( .Q(T14739_Q), .CK(T1638_Y), .D(T12326_Y));
KC_DFFHQ_X1 T13732 ( .Q(T13732_Q), .CK(T1638_Y), .D(T11919_Y));
KC_DFFHQ_X1 T13711 ( .Q(T13711_Q), .CK(T14677_Q), .D(T9687_Y));
KC_DFFHQ_X1 T13687 ( .Q(T13687_Q), .CK(T14677_Q), .D(T9606_Y));
KC_DFFHQ_X1 T13685 ( .Q(T13685_Q), .CK(T13340_Q), .D(T9606_Y));
KC_DFFHQ_X1 T6785 ( .Q(T6785_Q), .CK(T14865_Q), .D(T6716_Y));
KC_DFFHQ_X1 T14841 ( .Q(T14841_Q), .CK(T14865_Q), .D(T8533_Y));
KC_DFFHQ_X1 T14654 ( .Q(T14654_Q), .CK(T14864_Q), .D(T8533_Y));
KC_DFFHQ_X1 T14653 ( .Q(T14653_Q), .CK(T13950_Q), .D(T6716_Y));
KC_DFFHQ_X1 T14631 ( .Q(T14631_Q), .CK(T13951_Q), .D(T6716_Y));
KC_DFFHQ_X1 T14630 ( .Q(T14630_Q), .CK(T14008_Q), .D(T6716_Y));
KC_DFFHQ_X1 T13931 ( .Q(T13931_Q), .CK(T13952_Q), .D(T6716_Y));
KC_DFFHQ_X1 T13922 ( .Q(T13922_Q), .CK(T14865_Q), .D(T9757_Y));
KC_DFFHQ_X1 T13887 ( .Q(T13887_Q), .CK(T14865_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13848 ( .Q(T13848_Q), .CK(T13950_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13847 ( .Q(T13847_Q), .CK(T13953_Q), .D(T9757_Y));
KC_DFFHQ_X1 T13845 ( .Q(T13845_Q), .CK(T14864_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13832 ( .Q(T13832_Q), .CK(T13950_Q), .D(T8533_Y));
KC_DFFHQ_X1 T13802 ( .Q(T13802_Q), .CK(T14864_Q), .D(T9757_Y));
KC_DFFHQ_X1 T13800 ( .Q(T13800_Q), .CK(T13950_Q), .D(T9757_Y));
KC_DFFHQ_X1 T10247 ( .Q(T10247_Q), .CK(T13951_Q), .D(T9749_Y));
KC_DFFHQ_X1 T14075 ( .Q(T14075_Q), .CK(T14008_Q), .D(T9749_Y));
KC_DFFHQ_X1 T14060 ( .Q(T14060_Q), .CK(T13951_Q), .D(T9758_Y));
KC_DFFHQ_X1 T14058 ( .Q(T14058_Q), .CK(T14008_Q), .D(T9758_Y));
KC_DFFHQ_X1 T13990 ( .Q(T13990_Q), .CK(T13951_Q), .D(T9759_Y));
KC_DFFHQ_X1 T13988 ( .Q(T13988_Q), .CK(T13951_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13986 ( .Q(T13986_Q), .CK(T13952_Q), .D(T9759_Y));
KC_DFFHQ_X1 T13985 ( .Q(T13985_Q), .CK(T14008_Q), .D(T9759_Y));
KC_DFFHQ_X1 T13973 ( .Q(T13973_Q), .CK(T13952_Q), .D(T9808_Y));
KC_DFFHQ_X1 T14205 ( .Q(T14205_Q), .CK(T14236_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14383 ( .Q(T14383_Q), .CK(T13329_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14376 ( .Q(T14376_Q), .CK(T14591_Q), .D(T9904_Y));
KC_DFFHQ_X1 T14371 ( .Q(T14371_Q), .CK(T14591_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14818 ( .Q(T14818_Q), .CK(T14677_Q), .D(T10448_Y));
KC_DFFHQ_X1 T14817 ( .Q(T14817_Q), .CK(T14677_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13430 ( .Q(T13430_Q), .CK(T13492_Q), .D(T10448_Y));
KC_DFFHQ_X1 T13414 ( .Q(T13414_Q), .CK(T13491_Q), .D(T10448_Y));
KC_DFFHQ_X1 T13400 ( .Q(T13400_Q), .CK(T14702_Q), .D(T10448_Y));
KC_DFFHQ_X1 T14808 ( .Q(T14808_Q), .CK(T14682_Q), .D(T9601_Y));
KC_DFFHQ_X1 T14807 ( .Q(T14807_Q), .CK(T14682_Q), .D(T9600_Y));
KC_DFFHQ_X1 T14806 ( .Q(T14806_Q), .CK(T13630_Q), .D(T9600_Y));
KC_DFFHQ_X1 T14805 ( .Q(T14805_Q), .CK(T13642_Q), .D(T10443_Y));
KC_DFFHQ_X1 T13562 ( .Q(T13562_Q), .CK(T13682_Q), .D(T10453_Y));
KC_DFFHQ_X1 T13561 ( .Q(T13561_Q), .CK(T13682_Q), .D(T10443_Y));
KC_DFFHQ_X1 T13560 ( .Q(T13560_Q), .CK(T14703_Q), .D(T10453_Y));
KC_DFFHQ_X1 T13559 ( .Q(T13559_Q), .CK(T14703_Q), .D(T10443_Y));
KC_DFFHQ_X1 T13536 ( .Q(T13536_Q), .CK(T13446_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13535 ( .Q(T13535_Q), .CK(T13642_Q), .D(T10453_Y));
KC_DFFHQ_X1 T13534 ( .Q(T13534_Q), .CK(T13757_Q), .D(T10453_Y));
KC_DFFHQ_X1 T13533 ( .Q(T13533_Q), .CK(T13757_Q), .D(T10443_Y));
KC_DFFHQ_X1 T13516 ( .Q(T13516_Q), .CK(T13340_Q), .D(T10443_Y));
KC_DFFHQ_X1 T13515 ( .Q(T13515_Q), .CK(T13340_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13514 ( .Q(T13514_Q), .CK(T13340_Q), .D(T10453_Y));
KC_DFFHQ_X1 T13513 ( .Q(T13513_Q), .CK(T14677_Q), .D(T10443_Y));
KC_DFFHQ_X1 T14772 ( .Q(T14772_Q), .CK(T13445_Q), .D(T9600_Y));
KC_DFFHQ_X1 T14771 ( .Q(T14771_Q), .CK(T4977_Y), .D(T11926_Y));
KC_DFFHQ_X1 T13681 ( .Q(T13681_Q), .CK(T14767_Q), .D(T9601_Y));
KC_DFFHQ_X1 T13680 ( .Q(T13680_Q), .CK(T13490_Q), .D(T9601_Y));
KC_DFFHQ_X1 T13660 ( .Q(T13660_Q), .CK(T13745_Q), .D(T9600_Y));
KC_DFFHQ_X1 T13659 ( .Q(T13659_Q), .CK(T14683_Q), .D(T9599_Y));
KC_DFFHQ_X1 T13658 ( .Q(T13658_Q), .CK(T13745_Q), .D(T9599_Y));
KC_DFFHQ_X1 T13641 ( .Q(T13641_Q), .CK(T14683_Q), .D(T9600_Y));
KC_DFFHQ_X1 T13631 ( .Q(T13631_Q), .CK(T13446_Q), .D(T9601_Y));
KC_DFFHQ_X1 T14939 ( .Q(T14939_Q), .CK(T1638_Y), .D(T6755_Y));
KC_DFFHQ_X1 T14938 ( .Q(T14938_Q), .CK(T1638_Y), .D(T11936_Y));
KC_DFFHQ_X1 T14937 ( .Q(T14937_Q), .CK(T4977_Y), .D(T11933_Y));
KC_DFFHQ_X1 T14934 ( .Q(T14934_Q), .CK(T4977_Y), .D(T11955_Y));
KC_DFFHQ_X1 T14932 ( .Q(T14932_Q), .CK(T4977_Y), .D(T11939_Y));
KC_DFFHQ_X1 T13776 ( .Q(T13776_Q), .CK(T1638_Y), .D(T11122_Y));
KC_DFFHQ_X1 T13775 ( .Q(T13775_Q), .CK(T4977_Y), .D(T11123_Y));
KC_DFFHQ_X1 T13774 ( .Q(T13774_Q), .CK(T1638_Y), .D(T11126_Y));
KC_DFFHQ_X1 T13758 ( .Q(T13758_Q), .CK(T4977_Y), .D(T11133_Y));
KC_DFFHQ_X1 T13746 ( .Q(T13746_Q), .CK(T1638_Y), .D(T11135_Y));
KC_DFFHQ_X1 T14863 ( .Q(T14863_Q), .CK(T14864_Q), .D(T9758_Y));
KC_DFFHQ_X1 T13921 ( .Q(T13921_Q), .CK(T13937_Q), .D(T9757_Y));
KC_DFFHQ_X1 T13920 ( .Q(T13920_Q), .CK(T13937_Q), .D(T9758_Y));
KC_DFFHQ_X1 T13919 ( .Q(T13919_Q), .CK(T14865_Q), .D(T9760_Y));
KC_DFFHQ_X1 T13918 ( .Q(T13918_Q), .CK(T13937_Q), .D(T9759_Y));
KC_DFFHQ_X1 T13917 ( .Q(T13917_Q), .CK(T14865_Q), .D(T9759_Y));
KC_DFFHQ_X1 T13916 ( .Q(T13916_Q), .CK(T14865_Q), .D(T9758_Y));
KC_DFFHQ_X1 T13897 ( .Q(T13897_Q), .CK(T13937_Q), .D(T9760_Y));
KC_DFFHQ_X1 T13896 ( .Q(T13896_Q), .CK(T1638_Y), .D(T11943_Y));
KC_DFFHQ_X1 T13885 ( .Q(T13885_Q), .CK(T13950_Q), .D(T9749_Y));
KC_DFFHQ_X1 T13884 ( .Q(T13884_Q), .CK(T13950_Q), .D(T9760_Y));
KC_DFFHQ_X1 T13882 ( .Q(T13882_Q), .CK(T13950_Q), .D(T9758_Y));
KC_DFFHQ_X1 T14074 ( .Q(T14074_Q), .CK(T13952_Q), .D(T9749_Y));
KC_DFFHQ_X1 T14073 ( .Q(T14073_Q), .CK(T14625_Q), .D(T9760_Y));
KC_DFFHQ_X1 T14072 ( .Q(T14072_Q), .CK(T14625_Q), .D(T9749_Y));
KC_DFFHQ_X1 T14070 ( .Q(T14070_Q), .CK(T13953_Q), .D(T9749_Y));
KC_DFFHQ_X1 T14057 ( .Q(T14057_Q), .CK(T13953_Q), .D(T9759_Y));
KC_DFFHQ_X1 T14056 ( .Q(T14056_Q), .CK(T13953_Q), .D(T9758_Y));
KC_DFFHQ_X1 T14055 ( .Q(T14055_Q), .CK(T14625_Q), .D(T9759_Y));
KC_DFFHQ_X1 T14054 ( .Q(T14054_Q), .CK(T14625_Q), .D(T9758_Y));
KC_DFFHQ_X1 T14053 ( .Q(T14053_Q), .CK(T13952_Q), .D(T9760_Y));
KC_DFFHQ_X1 T14052 ( .Q(T14052_Q), .CK(T13953_Q), .D(T9760_Y));
KC_DFFHQ_X1 T14816 ( .Q(T14816_Q), .CK(T13663_Q), .D(T10456_Y));
KC_DFFHQ_X1 T14815 ( .Q(T14815_Q), .CK(T13663_Q), .D(T10447_Y));
KC_DFFHQ_X1 T13428 ( .Q(T13428_Q), .CK(T13634_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13427 ( .Q(T13427_Q), .CK(T13340_Q), .D(T10448_Y));
KC_DFFHQ_X1 T13413 ( .Q(T13413_Q), .CK(T13644_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13410 ( .Q(T13410_Q), .CK(T13644_Q), .D(T10456_Y));
KC_DFFHQ_X1 T13399 ( .Q(T13399_Q), .CK(T13663_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13398 ( .Q(T13398_Q), .CK(T13634_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13394 ( .Q(T13394_Q), .CK(T13634_Q), .D(T10456_Y));
KC_DFFHQ_X1 T14803 ( .Q(T14803_Q), .CK(T13642_Q), .D(T10446_Y));
KC_DFFHQ_X1 T14800 ( .Q(T14800_Q), .CK(T13664_Q), .D(T10447_Y));
KC_DFFHQ_X1 T14798 ( .Q(T14798_Q), .CK(T13664_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13558 ( .Q(T13558_Q), .CK(T13664_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13557 ( .Q(T13557_Q), .CK(T14703_Q), .D(T10448_Y));
KC_DFFHQ_X1 T13556 ( .Q(T13556_Q), .CK(T13621_Q), .D(T10447_Y));
KC_DFFHQ_X1 T13544 ( .Q(T13544_Q), .CK(T14703_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13543 ( .Q(T13543_Q), .CK(T13621_Q), .D(T10456_Y));
KC_DFFHQ_X1 T13531 ( .Q(T13531_Q), .CK(T13757_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13530 ( .Q(T13530_Q), .CK(T13757_Q), .D(T10448_Y));
KC_DFFHQ_X1 T13528 ( .Q(T13528_Q), .CK(T13664_Q), .D(T10456_Y));
KC_DFFHQ_X1 T13512 ( .Q(T13512_Q), .CK(T13682_Q), .D(T10448_Y));
KC_DFFHQ_X1 T13511 ( .Q(T13511_Q), .CK(T13621_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13509 ( .Q(T13509_Q), .CK(T13663_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13679 ( .Q(T13679_Q), .CK(T14767_Q), .D(T9599_Y));
KC_DFFHQ_X1 T13657 ( .Q(T13657_Q), .CK(T2495_Y), .D(T12520_Y));
KC_DFFHQ_X1 T13656 ( .Q(T13656_Q), .CK(T2495_Y), .D(T12521_Y));
KC_DFFHQ_X1 T13654 ( .Q(T13654_Q), .CK(T4977_Y), .D(T11924_Y));
KC_DFFHQ_X1 T13640 ( .Q(T13640_Q), .CK(T13490_Q), .D(T9599_Y));
KC_DFFHQ_X1 T13629 ( .Q(T13629_Q), .CK(T13446_Q), .D(T9599_Y));
KC_DFFHQ_X1 T14936 ( .Q(T14936_Q), .CK(T2495_Y), .D(T11953_Y));
KC_DFFHQ_X1 T14935 ( .Q(T14935_Q), .CK(T2495_Y), .D(T11116_Y));
KC_DFFHQ_X1 T14933 ( .Q(T14933_Q), .CK(T2495_Y), .D(T11952_Y));
KC_DFFHQ_X1 T14928 ( .Q(T14928_Q), .CK(T2495_Y), .D(T6759_Y));
KC_DFFHQ_X1 T13783 ( .Q(T13783_Q), .CK(T2495_Y), .D(T11130_Y));
KC_DFFHQ_X1 T13782 ( .Q(T13782_Q), .CK(T2495_Y), .D(T13003_Y));
KC_DFFHQ_X1 T13773 ( .Q(T13773_Q), .CK(T2495_Y), .D(T11131_Y));
KC_DFFHQ_X1 T13772 ( .Q(T13772_Q), .CK(T4977_Y), .D(T11132_Y));
KC_DFFHQ_X1 T13770 ( .Q(T13770_Q), .CK(T2495_Y), .D(T13001_Y));
KC_DFFHQ_X1 T13769 ( .Q(T13769_Q), .CK(T2495_Y), .D(T13002_Y));
KC_DFFHQ_X1 T14859 ( .Q(T14859_Q), .CK(T5315_Y), .D(T12587_Y));
KC_DFFHQ_X1 T14838 ( .Q(T14838_Q), .CK(T2495_Y), .D(T11940_Y));
KC_DFFHQ_X1 T13895 ( .Q(T13895_Q), .CK(T2495_Y), .D(T12591_Y));
KC_DFFHQ_X1 T13894 ( .Q(T13894_Q), .CK(T2495_Y), .D(T12933_Y));
KC_DFFHQ_X1 T14093 ( .Q(T14093_Q), .CK(T5315_Y), .D(T1110_Y));
KC_DFFHQ_X1 T14082 ( .Q(T14082_Q), .CK(T5315_Y), .D(T12672_Y));
KC_DFFHQ_X1 T14032 ( .Q(T14032_Q), .CK(T5315_Y), .D(T12676_Y));
KC_DFFHQ_X1 T14882 ( .Q(T14882_Q), .CK(T5315_Y), .D(T13209_Y));
KC_DFFHQ_X1 T14367 ( .Q(T14367_Q), .CK(T2047_Y), .D(T12757_Y));
KC_DFFHQ_X1 T14427 ( .Q(T14427_Q), .CK(T2047_Y), .D(T12763_Y));
KC_DFFHQ_X1 T14426 ( .Q(T14426_Q), .CK(T2047_Y), .D(T12768_Y));
KC_DFFHQ_X1 T14425 ( .Q(T14425_Q), .CK(T2047_Y), .D(T12762_Y));
KC_DFFHQ_X1 T14404 ( .Q(T14404_Q), .CK(T2047_Y), .D(T12758_Y));
KC_DFFHQ_X1 T14403 ( .Q(T14403_Q), .CK(T2047_Y), .D(T16263_Y));
KC_DFFHQ_X1 T14501 ( .Q(T14501_Q), .CK(T14481_Q), .D(T12142_Y));
KC_DFFHQ_X1 T14500 ( .Q(T14500_Q), .CK(T14481_Q), .D(T11359_Y));
KC_DFFHQ_X1 T14499 ( .Q(T14499_Q), .CK(T14481_Q), .D(T13072_Y));
KC_DFFHQ_X1 T14498 ( .Q(T14498_Q), .CK(T14481_Q), .D(T15848_Y));
KC_DFFHQ_X1 T14495 ( .Q(T14495_Q), .CK(T2047_Y), .D(T5994_Y));
KC_DFFHQ_X1 T14494 ( .Q(T14494_Q), .CK(T2047_Y), .D(T5993_Y));
KC_DFFHQ_X1 T14957 ( .Q(T14957_Q), .CK(T14532_Q), .D(T2684_Y));
KC_DFFHQ_X1 T14954 ( .Q(T14954_Q), .CK(T14532_Q), .D(T2694_Y));
KC_DFFHQ_X1 T14537 ( .Q(T14537_Q), .CK(T14532_Q), .D(T10896_Y));
KC_DFFHQ_X1 T14535 ( .Q(T14535_Q), .CK(T14532_Q), .D(T2697_Y));
KC_DFFHQ_X1 T14533 ( .Q(T14533_Q), .CK(T14532_Q), .D(T2680_Y));
KC_DFFHQ_X1 T14528 ( .Q(T14528_Q), .CK(T14532_Q), .D(T5785_Y));
KC_DFFHQ_X1 T14527 ( .Q(T14527_Q), .CK(T14532_Q), .D(T10897_Y));
KC_DFFHQ_X1 T14525 ( .Q(T14525_Q), .CK(T14532_Q), .D(T11340_Y));
KC_DFFHQ_X1 T14814 ( .Q(T14814_Q), .CK(T14791_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13425 ( .Q(T13425_Q), .CK(T13667_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13424 ( .Q(T13424_Q), .CK(T14790_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13423 ( .Q(T13423_Q), .CK(T13519_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13411 ( .Q(T13411_Q), .CK(T13667_Q), .D(T10456_Y));
KC_DFFHQ_X1 T13409 ( .Q(T13409_Q), .CK(T13519_Q), .D(T10456_Y));
KC_DFFHQ_X1 T13407 ( .Q(T13407_Q), .CK(T14790_Q), .D(T10456_Y));
KC_DFFHQ_X1 T13397 ( .Q(T13397_Q), .CK(T13667_Q), .D(T10447_Y));
KC_DFFHQ_X1 T13396 ( .Q(T13396_Q), .CK(T13634_Q), .D(T10447_Y));
KC_DFFHQ_X1 T13392 ( .Q(T13392_Q), .CK(T13519_Q), .D(T10447_Y));
KC_DFFHQ_X1 T13391 ( .Q(T13391_Q), .CK(T14790_Q), .D(T10447_Y));
KC_DFFHQ_X1 T14801 ( .Q(T14801_Q), .CK(T13644_Q), .D(T9592_Y));
KC_DFFHQ_X1 T14799 ( .Q(T14799_Q), .CK(T13663_Q), .D(T9592_Y));
KC_DFFHQ_X1 T14797 ( .Q(T14797_Q), .CK(T14791_Q), .D(T9593_Y));
KC_DFFHQ_X1 T14796 ( .Q(T14796_Q), .CK(T14790_Q), .D(T9593_Y));
KC_DFFHQ_X1 T13555 ( .Q(T13555_Q), .CK(T13667_Q), .D(T9589_Y));
KC_DFFHQ_X1 T13554 ( .Q(T13554_Q), .CK(T13634_Q), .D(T9589_Y));
KC_DFFHQ_X1 T13553 ( .Q(T13553_Q), .CK(T13519_Q), .D(T9589_Y));
KC_DFFHQ_X1 T13551 ( .Q(T13551_Q), .CK(T14791_Q), .D(T9592_Y));
KC_DFFHQ_X1 T13542 ( .Q(T13542_Q), .CK(T14790_Q), .D(T9589_Y));
KC_DFFHQ_X1 T13526 ( .Q(T13526_Q), .CK(T13519_Q), .D(T9592_Y));
KC_DFFHQ_X1 T13525 ( .Q(T13525_Q), .CK(T14790_Q), .D(T9592_Y));
KC_DFFHQ_X1 T13524 ( .Q(T13524_Q), .CK(T13519_Q), .D(T9593_Y));
KC_DFFHQ_X1 T13508 ( .Q(T13508_Q), .CK(T14790_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13507 ( .Q(T13507_Q), .CK(T14791_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13506 ( .Q(T13506_Q), .CK(T13519_Q), .D(T10454_Y));
KC_DFFHQ_X1 T14764 ( .Q(T14764_Q), .CK(T13619_Q), .D(T9644_Y));
KC_DFFHQ_X1 T13677 ( .Q(T13677_Q), .CK(T13667_Q), .D(T9592_Y));
KC_DFFHQ_X1 T13676 ( .Q(T13676_Q), .CK(T13634_Q), .D(T9592_Y));
KC_DFFHQ_X1 T13674 ( .Q(T13674_Q), .CK(T13664_Q), .D(T9593_Y));
KC_DFFHQ_X1 T13672 ( .Q(T13672_Q), .CK(T13634_Q), .D(T9593_Y));
KC_DFFHQ_X1 T13653 ( .Q(T13653_Q), .CK(T3026_Y), .D(T12519_Y));
KC_DFFHQ_X1 T13651 ( .Q(T13651_Q), .CK(T13617_Q), .D(T9644_Y));
KC_DFFHQ_X1 T13639 ( .Q(T13639_Q), .CK(T3026_Y), .D(T12518_Y));
KC_DFFHQ_X1 T13637 ( .Q(T13637_Q), .CK(T13620_Q), .D(T9644_Y));
KC_DFFHQ_X1 T13626 ( .Q(T13626_Q), .CK(T13621_Q), .D(T9592_Y));
KC_DFFHQ_X1 T13624 ( .Q(T13624_Q), .CK(T13621_Q), .D(T9593_Y));
KC_DFFHQ_X1 T14931 ( .Q(T14931_Q), .CK(T2495_Y), .D(T12945_Y));
KC_DFFHQ_X1 T14929 ( .Q(T14929_Q), .CK(T13927_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14926 ( .Q(T14926_Q), .CK(T14067_Q), .D(T9740_Y));
KC_DFFHQ_X1 T14925 ( .Q(T14925_Q), .CK(T13927_Q), .D(T9740_Y));
KC_DFFHQ_X1 T14924 ( .Q(T14924_Q), .CK(T14067_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14922 ( .Q(T14922_Q), .CK(T13926_Q), .D(T9740_Y));
KC_DFFHQ_X1 T13781 ( .Q(T13781_Q), .CK(T3026_Y), .D(T12547_Y));
KC_DFFHQ_X1 T13767 ( .Q(T13767_Q), .CK(T3026_Y), .D(T13000_Y));
KC_DFFHQ_X1 T13755 ( .Q(T13755_Q), .CK(T3026_Y), .D(T12998_Y));
KC_DFFHQ_X1 T14858 ( .Q(T14858_Q), .CK(T14077_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14854 ( .Q(T14854_Q), .CK(T14079_Q), .D(T9741_Y));
KC_DFFHQ_X1 T14835 ( .Q(T14835_Q), .CK(T14076_Q), .D(T9844_Y));
KC_DFFHQ_X1 T14829 ( .Q(T14829_Q), .CK(T13927_Q), .D(T9741_Y));
KC_DFFHQ_X1 T13929 ( .Q(T13929_Q), .CK(T14080_Q), .D(T9742_Y));
KC_DFFHQ_X1 T13928 ( .Q(T13928_Q), .CK(T14079_Q), .D(T9740_Y));
KC_DFFHQ_X1 T13913 ( .Q(T13913_Q), .CK(T14080_Q), .D(T9844_Y));
KC_DFFHQ_X1 T13912 ( .Q(T13912_Q), .CK(T14080_Q), .D(T9740_Y));
KC_DFFHQ_X1 T13911 ( .Q(T13911_Q), .CK(T14076_Q), .D(T9741_Y));
KC_DFFHQ_X1 T13910 ( .Q(T13910_Q), .CK(T14077_Q), .D(T9740_Y));
KC_DFFHQ_X1 T13893 ( .Q(T13893_Q), .CK(T14076_Q), .D(T9740_Y));
KC_DFFHQ_X1 T13881 ( .Q(T13881_Q), .CK(T14077_Q), .D(T9844_Y));
KC_DFFHQ_X1 T13880 ( .Q(T13880_Q), .CK(T14077_Q), .D(T9741_Y));
KC_DFFHQ_X1 T13879 ( .Q(T13879_Q), .CK(T14080_Q), .D(T9741_Y));
KC_DFFHQ_X1 T14091 ( .Q(T14091_Q), .CK(T14353_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14090 ( .Q(T14090_Q), .CK(T14355_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14083 ( .Q(T14083_Q), .CK(T5315_Y), .D(T12671_Y));
KC_DFFHQ_X1 T14081 ( .Q(T14081_Q), .CK(T5315_Y), .D(T12675_Y));
KC_DFFHQ_X1 T14069 ( .Q(T14069_Q), .CK(T5315_Y), .D(T12657_Y));
KC_DFFHQ_X1 T14068 ( .Q(T14068_Q), .CK(T14031_Q), .D(T9844_Y));
KC_DFFHQ_X1 T14050 ( .Q(T14050_Q), .CK(T14079_Q), .D(T9844_Y));
KC_DFFHQ_X1 T14049 ( .Q(T14049_Q), .CK(T14031_Q), .D(T9741_Y));
KC_DFFHQ_X1 T14047 ( .Q(T14047_Q), .CK(T14078_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14046 ( .Q(T14046_Q), .CK(T14031_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14045 ( .Q(T14045_Q), .CK(T14078_Q), .D(T9741_Y));
KC_DFFHQ_X1 T14044 ( .Q(T14044_Q), .CK(T14078_Q), .D(T9844_Y));
KC_DFFHQ_X1 T14030 ( .Q(T14030_Q), .CK(T14346_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14893 ( .Q(T14893_Q), .CK(T3122_Y), .D(T12716_Y));
KC_DFFHQ_X1 T14890 ( .Q(T14890_Q), .CK(T14354_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14198 ( .Q(T14198_Q), .CK(T3122_Y), .D(T12942_Y));
KC_DFFHQ_X1 T14197 ( .Q(T14197_Q), .CK(T14331_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14194 ( .Q(T14194_Q), .CK(T14354_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14193 ( .Q(T14193_Q), .CK(T14355_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14192 ( .Q(T14192_Q), .CK(T14353_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14183 ( .Q(T14183_Q), .CK(T14331_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14181 ( .Q(T14181_Q), .CK(T14352_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14172 ( .Q(T14172_Q), .CK(T3122_Y), .D(T12714_Y));
KC_DFFHQ_X1 T14169 ( .Q(T14169_Q), .CK(T14331_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14168 ( .Q(T14168_Q), .CK(T14352_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14151 ( .Q(T14151_Q), .CK(T3122_Y), .D(T12717_Y));
KC_DFFHQ_X1 T14150 ( .Q(T14150_Q), .CK(T14354_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14148 ( .Q(T14148_Q), .CK(T14352_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14147 ( .Q(T14147_Q), .CK(T14331_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14365 ( .Q(T14365_Q), .CK(T14331_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14364 ( .Q(T14364_Q), .CK(T14354_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14362 ( .Q(T14362_Q), .CK(T14352_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14360 ( .Q(T14360_Q), .CK(T14355_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14359 ( .Q(T14359_Q), .CK(T14353_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14357 ( .Q(T14357_Q), .CK(T14352_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14344 ( .Q(T14344_Q), .CK(T14354_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14343 ( .Q(T14343_Q), .CK(T14331_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14341 ( .Q(T14341_Q), .CK(T14352_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14339 ( .Q(T14339_Q), .CK(T14353_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14323 ( .Q(T14323_Q), .CK(T14355_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14318 ( .Q(T14318_Q), .CK(T14354_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14317 ( .Q(T14317_Q), .CK(T14355_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14316 ( .Q(T14316_Q), .CK(T14331_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14315 ( .Q(T14315_Q), .CK(T14353_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14313 ( .Q(T14313_Q), .CK(T14346_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14300 ( .Q(T14300_Q), .CK(T14353_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14299 ( .Q(T14299_Q), .CK(T14352_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14298 ( .Q(T14298_Q), .CK(T14355_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14296 ( .Q(T14296_Q), .CK(T14352_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14909 ( .Q(T14909_Q), .CK(T14412_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14907 ( .Q(T14907_Q), .CK(T14394_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14450 ( .Q(T14450_Q), .CK(T14392_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14449 ( .Q(T14449_Q), .CK(T14406_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14447 ( .Q(T14447_Q), .CK(T14412_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14446 ( .Q(T14446_Q), .CK(T14393_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14444 ( .Q(T14444_Q), .CK(T14405_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14433 ( .Q(T14433_Q), .CK(T14393_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14432 ( .Q(T14432_Q), .CK(T14412_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14424 ( .Q(T14424_Q), .CK(T14406_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14423 ( .Q(T14423_Q), .CK(T14392_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14421 ( .Q(T14421_Q), .CK(T14405_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14420 ( .Q(T14420_Q), .CK(T14394_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14419 ( .Q(T14419_Q), .CK(T14405_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14402 ( .Q(T14402_Q), .CK(T14406_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14401 ( .Q(T14401_Q), .CK(T14392_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14400 ( .Q(T14400_Q), .CK(T14394_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14399 ( .Q(T14399_Q), .CK(T14412_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14396 ( .Q(T14396_Q), .CK(T14393_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14521 ( .Q(T14521_Q), .CK(T14519_Q), .D(T5469_Y));
KC_DFFHQ_X1 T14520 ( .Q(T14520_Q), .CK(T3199_Y), .D(T12126_Y));
KC_DFFHQ_X1 T14516 ( .Q(T14516_Q), .CK(T3198_Y), .D(T3186_Y));
KC_DFFHQ_X1 T14515 ( .Q(T14515_Q), .CK(T3198_Y), .D(T10267_Y));
KC_DFFHQ_X1 T14496 ( .Q(T14496_Q), .CK(T3199_Y), .D(T12784_Y));
KC_DFFHQ_X1 T14491 ( .Q(T14491_Q), .CK(T3198_Y), .D(T12783_Y));
KC_DFFHQ_X1 T14490 ( .Q(T14490_Q), .CK(T3198_Y), .D(T12779_Y));
KC_DFFHQ_X1 T14479 ( .Q(T14479_Q), .CK(T3199_Y), .D(T12778_Y));
KC_DFFHQ_X1 T14478 ( .Q(T14478_Q), .CK(T3199_Y), .D(T12772_Y));
KC_DFFHQ_X1 T14476 ( .Q(T14476_Q), .CK(T3198_Y), .D(T12776_Y));
KC_DFFHQ_X1 T14474 ( .Q(T14474_Q), .CK(T3199_Y), .D(T12773_Y));
KC_DFFHQ_X1 T14464 ( .Q(T14464_Q), .CK(T3198_Y), .D(T12775_Y));
KC_DFFHQ_X1 T14462 ( .Q(T14462_Q), .CK(T3199_Y), .D(T12774_Y));
KC_DFFHQ_X1 T14956 ( .Q(T14956_Q), .CK(T14524_Q), .D(T15866_Y));
KC_DFFHQ_X1 T14949 ( .Q(T14949_Q), .CK(T3199_Y), .D(T11958_Y));
KC_DFFHQ_X1 T14534 ( .Q(T14534_Q), .CK(T14524_Q), .D(T11314_Y));
KC_DFFHQ_X1 T14530 ( .Q(T14530_Q), .CK(T14524_Q), .D(T3220_Y));
KC_DFFHQ_X1 T14529 ( .Q(T14529_Q), .CK(T14524_Q), .D(T11333_Y));
KC_DFFHQ_X1 T14543 ( .Q(T14543_Q), .CK(T14539_Q), .D(T11403_Y));
KC_DFFHQ_X1 T14541 ( .Q(T14541_Q), .CK(T14539_Q), .D(T11382_Y));
KC_DFFHQ_X1 T14813 ( .Q(T14813_Q), .CK(T13619_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13422 ( .Q(T13422_Q), .CK(T14775_Q), .D(T15199_Y));
KC_DFFHQ_X1 T13420 ( .Q(T13420_Q), .CK(T13666_Q), .D(T15199_Y));
KC_DFFHQ_X1 T13419 ( .Q(T13419_Q), .CK(T13619_Q), .D(T15199_Y));
KC_DFFHQ_X1 T13405 ( .Q(T13405_Q), .CK(T13645_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13404 ( .Q(T13404_Q), .CK(T13666_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13403 ( .Q(T13403_Q), .CK(T13618_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13390 ( .Q(T13390_Q), .CK(T14775_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13389 ( .Q(T13389_Q), .CK(T13633_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13388 ( .Q(T13388_Q), .CK(T13618_Q), .D(T15199_Y));
KC_DFFHQ_X1 T14794 ( .Q(T14794_Q), .CK(T13663_Q), .D(T9591_Y));
KC_DFFHQ_X1 T14793 ( .Q(T14793_Q), .CK(T14790_Q), .D(T9591_Y));
KC_DFFHQ_X1 T13550 ( .Q(T13550_Q), .CK(T13617_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13548 ( .Q(T13548_Q), .CK(T13620_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13547 ( .Q(T13547_Q), .CK(T13620_Q), .D(T15199_Y));
KC_DFFHQ_X1 T13540 ( .Q(T13540_Q), .CK(T13617_Q), .D(T15199_Y));
KC_DFFHQ_X1 T13522 ( .Q(T13522_Q), .CK(T13519_Q), .D(T9591_Y));
KC_DFFHQ_X1 T13505 ( .Q(T13505_Q), .CK(T13618_Q), .D(T6443_Y));
KC_DFFHQ_X1 T14760 ( .Q(T14760_Q), .CK(T14775_Q), .D(T9648_Y));
KC_DFFHQ_X1 T14759 ( .Q(T14759_Q), .CK(T14775_Q), .D(T15252_Y));
KC_DFFHQ_X1 T14758 ( .Q(T14758_Q), .CK(T13645_Q), .D(T9644_Y));
KC_DFFHQ_X1 T13673 ( .Q(T13673_Q), .CK(T13617_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13671 ( .Q(T13671_Q), .CK(T13667_Q), .D(T9591_Y));
KC_DFFHQ_X1 T13669 ( .Q(T13669_Q), .CK(T13664_Q), .D(T9591_Y));
KC_DFFHQ_X1 T13668 ( .Q(T13668_Q), .CK(T13634_Q), .D(T9591_Y));
KC_DFFHQ_X1 T13650 ( .Q(T13650_Q), .CK(T13619_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13649 ( .Q(T13649_Q), .CK(T13619_Q), .D(T15252_Y));
KC_DFFHQ_X1 T13648 ( .Q(T13648_Q), .CK(T13633_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13646 ( .Q(T13646_Q), .CK(T13619_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13636 ( .Q(T13636_Q), .CK(T13620_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13635 ( .Q(T13635_Q), .CK(T13620_Q), .D(T15252_Y));
KC_DFFHQ_X1 T13623 ( .Q(T13623_Q), .CK(T13621_Q), .D(T9591_Y));
KC_DFFHQ_X1 T14920 ( .Q(T14920_Q), .CK(T14036_Q), .D(T9727_Y));
KC_DFFHQ_X1 T14919 ( .Q(T14919_Q), .CK(T14036_Q), .D(T9734_Y));
KC_DFFHQ_X1 T14918 ( .Q(T14918_Q), .CK(T13666_Q), .D(T15252_Y));
KC_DFFHQ_X1 T14916 ( .Q(T14916_Q), .CK(T14036_Q), .D(T9733_Y));
KC_DFFHQ_X1 T14915 ( .Q(T14915_Q), .CK(T14062_Q), .D(T9734_Y));
KC_DFFHQ_X1 T13765 ( .Q(T13765_Q), .CK(T13666_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13764 ( .Q(T13764_Q), .CK(T13645_Q), .D(T15252_Y));
KC_DFFHQ_X1 T13754 ( .Q(T13754_Q), .CK(T13666_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13752 ( .Q(T13752_Q), .CK(T13633_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13751 ( .Q(T13751_Q), .CK(T13666_Q), .D(T9644_Y));
KC_DFFHQ_X1 T14852 ( .Q(T14852_Q), .CK(T14062_Q), .D(T10492_Y));
KC_DFFHQ_X1 T14831 ( .Q(T14831_Q), .CK(T13926_Q), .D(T9844_Y));
KC_DFFHQ_X1 T14827 ( .Q(T14827_Q), .CK(T14061_Q), .D(T9727_Y));
KC_DFFHQ_X1 T14826 ( .Q(T14826_Q), .CK(T14062_Q), .D(T9727_Y));
KC_DFFHQ_X1 T13925 ( .Q(T13925_Q), .CK(T14061_Q), .D(T10492_Y));
KC_DFFHQ_X1 T13909 ( .Q(T13909_Q), .CK(T14061_Q), .D(T9733_Y));
KC_DFFHQ_X1 T13908 ( .Q(T13908_Q), .CK(T14040_Q), .D(T9734_Y));
KC_DFFHQ_X1 T13906 ( .Q(T13906_Q), .CK(T14061_Q), .D(T125_Q));
KC_DFFHQ_X1 T13904 ( .Q(T13904_Q), .CK(T14040_Q), .D(T9733_Y));
KC_DFFHQ_X1 T13903 ( .Q(T13903_Q), .CK(T14061_Q), .D(T9734_Y));
KC_DFFHQ_X1 T13892 ( .Q(T13892_Q), .CK(T14040_Q), .D(T9727_Y));
KC_DFFHQ_X1 T13878 ( .Q(T13878_Q), .CK(T14061_Q), .D(T9735_Y));
KC_DFFHQ_X1 T13876 ( .Q(T13876_Q), .CK(T14040_Q), .D(T10492_Y));
KC_DFFHQ_X1 T13875 ( .Q(T13875_Q), .CK(T14843_Q), .D(T10492_Y));
KC_DFFHQ_X1 T14089 ( .Q(T14089_Q), .CK(T14025_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14087 ( .Q(T14087_Q), .CK(T14084_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14066 ( .Q(T14066_Q), .CK(T14040_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14065 ( .Q(T14065_Q), .CK(T14061_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14064 ( .Q(T14064_Q), .CK(T14062_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14043 ( .Q(T14043_Q), .CK(T14843_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14041 ( .Q(T14041_Q), .CK(T14036_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14029 ( .Q(T14029_Q), .CK(T14028_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14889 ( .Q(T14889_Q), .CK(T14321_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14888 ( .Q(T14888_Q), .CK(T14028_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14874 ( .Q(T14874_Q), .CK(T14866_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14196 ( .Q(T14196_Q), .CK(T14332_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14191 ( .Q(T14191_Q), .CK(T14866_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14190 ( .Q(T14190_Q), .CK(T14028_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14189 ( .Q(T14189_Q), .CK(T14866_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14180 ( .Q(T14180_Q), .CK(T14025_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14171 ( .Q(T14171_Q), .CK(T14332_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14166 ( .Q(T14166_Q), .CK(T14321_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14165 ( .Q(T14165_Q), .CK(T14025_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14163 ( .Q(T14163_Q), .CK(T14084_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14161 ( .Q(T14161_Q), .CK(T14084_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14160 ( .Q(T14160_Q), .CK(T14321_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14149 ( .Q(T14149_Q), .CK(T14332_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14146 ( .Q(T14146_Q), .CK(T14867_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14145 ( .Q(T14145_Q), .CK(T14084_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14144 ( .Q(T14144_Q), .CK(T14025_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14143 ( .Q(T14143_Q), .CK(T14084_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14142 ( .Q(T14142_Q), .CK(T14321_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14358 ( .Q(T14358_Q), .CK(T14353_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14356 ( .Q(T14356_Q), .CK(T14333_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14337 ( .Q(T14337_Q), .CK(T14355_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14336 ( .Q(T14336_Q), .CK(T14321_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14335 ( .Q(T14335_Q), .CK(T14346_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14334 ( .Q(T14334_Q), .CK(T14332_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14324 ( .Q(T14324_Q), .CK(T14333_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14322 ( .Q(T14322_Q), .CK(T14332_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14312 ( .Q(T14312_Q), .CK(T16467_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14310 ( .Q(T14310_Q), .CK(T14321_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14309 ( .Q(T14309_Q), .CK(T14866_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14308 ( .Q(T14308_Q), .CK(T14321_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14307 ( .Q(T14307_Q), .CK(T14332_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14302 ( .Q(T14302_Q), .CK(T14332_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14295 ( .Q(T14295_Q), .CK(T14867_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14293 ( .Q(T14293_Q), .CK(T14867_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14292 ( .Q(T14292_Q), .CK(T14321_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14291 ( .Q(T14291_Q), .CK(T14028_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14289 ( .Q(T14289_Q), .CK(T16467_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14288 ( .Q(T14288_Q), .CK(T14332_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14905 ( .Q(T14905_Q), .CK(T14392_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14903 ( .Q(T14903_Q), .CK(T14392_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14443 ( .Q(T14443_Q), .CK(T14412_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14442 ( .Q(T14442_Q), .CK(T14406_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14441 ( .Q(T14441_Q), .CK(T14412_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14439 ( .Q(T14439_Q), .CK(T14394_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14431 ( .Q(T14431_Q), .CK(T14405_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14430 ( .Q(T14430_Q), .CK(T14394_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14418 ( .Q(T14418_Q), .CK(T14394_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14417 ( .Q(T14417_Q), .CK(T14393_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14415 ( .Q(T14415_Q), .CK(T14393_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14414 ( .Q(T14414_Q), .CK(T14412_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14413 ( .Q(T14413_Q), .CK(T14406_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14395 ( .Q(T14395_Q), .CK(T14392_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14518 ( .Q(T14518_Q), .CK(T14519_Q), .D(T11331_Y));
KC_DFFHQ_X1 T14514 ( .Q(T14514_Q), .CK(T14948_Q), .D(T3808_Y));
KC_DFFHQ_X1 T14513 ( .Q(T14513_Q), .CK(T14944_Q), .D(T16221_Y));
KC_DFFHQ_X1 T14512 ( .Q(T14512_Q), .CK(T14531_Q), .D(T16223_Y));
KC_DFFHQ_X1 T14510 ( .Q(T14510_Q), .CK(T14948_Q), .D(T11324_Y));
KC_DFFHQ_X1 T14509 ( .Q(T14509_Q), .CK(T14531_Q), .D(T16114_Y));
KC_DFFHQ_X1 T14506 ( .Q(T14506_Q), .CK(T14392_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14505 ( .Q(T14505_Q), .CK(T14394_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14489 ( .Q(T14489_Q), .CK(T14944_Q), .D(T16215_Y));
KC_DFFHQ_X1 T14487 ( .Q(T14487_Q), .CK(T14944_Q), .D(T16229_Y));
KC_DFFHQ_X1 T14486 ( .Q(T14486_Q), .CK(T14944_Q), .D(T16218_Y));
KC_DFFHQ_X1 T14485 ( .Q(T14485_Q), .CK(T14944_Q), .D(T16216_Y));
KC_DFFHQ_X1 T14477 ( .Q(T14477_Q), .CK(T3198_Y), .D(T12780_Y));
KC_DFFHQ_X1 T14473 ( .Q(T14473_Q), .CK(T14531_Q), .D(T16212_Y));
KC_DFFHQ_X1 T14471 ( .Q(T14471_Q), .CK(T14531_Q), .D(T16228_Y));
KC_DFFHQ_X1 T14470 ( .Q(T14470_Q), .CK(T14944_Q), .D(T16214_Y));
KC_DFFHQ_X1 T14469 ( .Q(T14469_Q), .CK(T14531_Q), .D(T10238_Y));
KC_DFFHQ_X1 T14468 ( .Q(T14468_Q), .CK(T14531_Q), .D(T16217_Y));
KC_DFFHQ_X1 T14463 ( .Q(T14463_Q), .CK(T14944_Q), .D(T16226_Y));
KC_DFFHQ_X1 T14460 ( .Q(T14460_Q), .CK(T14531_Q), .D(T16224_Y));
KC_DFFHQ_X1 T14945 ( .Q(T14945_Q), .CK(T14944_Q), .D(T8440_Y));
KC_DFFHQ_X1 T13418 ( .Q(T13418_Q), .CK(T13645_Q), .D(T6443_Y));
KC_DFFHQ_X1 T13417 ( .Q(T13417_Q), .CK(T13665_Q), .D(T6443_Y));
KC_DFFHQ_X1 T13402 ( .Q(T13402_Q), .CK(T13665_Q), .D(T15199_Y));
KC_DFFHQ_X1 T13387 ( .Q(T13387_Q), .CK(T13645_Q), .D(T15199_Y));
KC_DFFHQ_X1 T14792 ( .Q(T14792_Q), .CK(T13633_Q), .D(T9602_Y));
KC_DFFHQ_X1 T13546 ( .Q(T13546_Q), .CK(T14775_Q), .D(T6443_Y));
KC_DFFHQ_X1 T13545 ( .Q(T13545_Q), .CK(T13665_Q), .D(T9602_Y));
KC_DFFHQ_X1 T13539 ( .Q(T13539_Q), .CK(T13645_Q), .D(T9602_Y));
KC_DFFHQ_X1 T13521 ( .Q(T13521_Q), .CK(T14775_Q), .D(T9602_Y));
KC_DFFHQ_X1 T13520 ( .Q(T13520_Q), .CK(T13620_Q), .D(T9602_Y));
KC_DFFHQ_X1 T14914 ( .Q(T14914_Q), .CK(T14034_Q), .D(T9733_Y));
KC_DFFHQ_X1 T14913 ( .Q(T14913_Q), .CK(T14842_Q), .D(T9735_Y));
KC_DFFHQ_X1 T14912 ( .Q(T14912_Q), .CK(T14034_Q), .D(T9734_Y));
KC_DFFHQ_X1 T14911 ( .Q(T14911_Q), .CK(T14035_Q), .D(T9727_Y));
KC_DFFHQ_X1 T14910 ( .Q(T14910_Q), .CK(T14035_Q), .D(T9734_Y));
KC_DFFHQ_X1 T13780 ( .Q(T13780_Q), .CK(T14033_Q), .D(T9727_Y));
KC_DFFHQ_X1 T13779 ( .Q(T13779_Q), .CK(T14033_Q), .D(T9735_Y));
KC_DFFHQ_X1 T13778 ( .Q(T13778_Q), .CK(T14033_Q), .D(T9733_Y));
KC_DFFHQ_X1 T13762 ( .Q(T13762_Q), .CK(T14033_Q), .D(T9734_Y));
KC_DFFHQ_X1 T13761 ( .Q(T13761_Q), .CK(T14842_Q), .D(T9727_Y));
KC_DFFHQ_X1 T13760 ( .Q(T13760_Q), .CK(T14842_Q), .D(T9733_Y));
KC_DFFHQ_X1 T13759 ( .Q(T13759_Q), .CK(T13665_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13750 ( .Q(T13750_Q), .CK(T13645_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13749 ( .Q(T13749_Q), .CK(T14842_Q), .D(T9734_Y));
KC_DFFHQ_X1 T13748 ( .Q(T13748_Q), .CK(T14034_Q), .D(T9727_Y));
KC_DFFHQ_X1 T13747 ( .Q(T13747_Q), .CK(T13665_Q), .D(T15252_Y));
KC_DFFHQ_X1 T14849 ( .Q(T14849_Q), .CK(T14033_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14848 ( .Q(T14848_Q), .CK(T14842_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14847 ( .Q(T14847_Q), .CK(T14035_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14846 ( .Q(T14846_Q), .CK(T14062_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14823 ( .Q(T14823_Q), .CK(T14036_Q), .D(T125_Q));
KC_DFFHQ_X1 T14822 ( .Q(T14822_Q), .CK(T14033_Q), .D(T125_Q));
KC_DFFHQ_X1 T14821 ( .Q(T14821_Q), .CK(T14034_Q), .D(T9735_Y));
KC_DFFHQ_X1 T14820 ( .Q(T14820_Q), .CK(T14035_Q), .D(T125_Q));
KC_DFFHQ_X1 T13924 ( .Q(T13924_Q), .CK(T14034_Q), .D(T10491_Y));
KC_DFFHQ_X1 T13902 ( .Q(T13902_Q), .CK(T14062_Q), .D(T9735_Y));
KC_DFFHQ_X1 T13901 ( .Q(T13901_Q), .CK(T14033_Q), .D(T10492_Y));
KC_DFFHQ_X1 T13900 ( .Q(T13900_Q), .CK(T14843_Q), .D(T9735_Y));
KC_DFFHQ_X1 T13899 ( .Q(T13899_Q), .CK(T14035_Q), .D(T9735_Y));
KC_DFFHQ_X1 T13891 ( .Q(T13891_Q), .CK(T14842_Q), .D(T125_Q));
KC_DFFHQ_X1 T13890 ( .Q(T13890_Q), .CK(T14034_Q), .D(T125_Q));
KC_DFFHQ_X1 T13889 ( .Q(T13889_Q), .CK(T14843_Q), .D(T125_Q));
KC_DFFHQ_X1 T13888 ( .Q(T13888_Q), .CK(T14062_Q), .D(T125_Q));
KC_DFFHQ_X1 T13874 ( .Q(T13874_Q), .CK(T14842_Q), .D(T10492_Y));
KC_DFFHQ_X1 T13873 ( .Q(T13873_Q), .CK(T14034_Q), .D(T10492_Y));
KC_DFFHQ_X1 T13872 ( .Q(T13872_Q), .CK(T14036_Q), .D(T9735_Y));
KC_DFFHQ_X1 T14086 ( .Q(T14086_Q), .CK(T14154_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14085 ( .Q(T14085_Q), .CK(T14153_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14063 ( .Q(T14063_Q), .CK(T14033_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14039 ( .Q(T14039_Q), .CK(T14034_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14038 ( .Q(T14038_Q), .CK(T14842_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14037 ( .Q(T14037_Q), .CK(T14036_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14027 ( .Q(T14027_Q), .CK(T14026_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14887 ( .Q(T14887_Q), .CK(T16467_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14886 ( .Q(T14886_Q), .CK(T14026_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14885 ( .Q(T14885_Q), .CK(T14866_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14871 ( .Q(T14871_Q), .CK(T14025_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14870 ( .Q(T14870_Q), .CK(T14026_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14869 ( .Q(T14869_Q), .CK(T16467_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14868 ( .Q(T14868_Q), .CK(T14867_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14188 ( .Q(T14188_Q), .CK(T14026_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14187 ( .Q(T14187_Q), .CK(T14154_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14186 ( .Q(T14186_Q), .CK(T14153_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14178 ( .Q(T14178_Q), .CK(T14867_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14177 ( .Q(T14177_Q), .CK(T14026_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14176 ( .Q(T14176_Q), .CK(T16467_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14175 ( .Q(T14175_Q), .CK(T14084_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14159 ( .Q(T14159_Q), .CK(T14025_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14158 ( .Q(T14158_Q), .CK(T14154_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14157 ( .Q(T14157_Q), .CK(T14025_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14156 ( .Q(T14156_Q), .CK(T14153_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14155 ( .Q(T14155_Q), .CK(T14084_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14141 ( .Q(T14141_Q), .CK(T14154_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14139 ( .Q(T14139_Q), .CK(T14153_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14351 ( .Q(T14351_Q), .CK(T14153_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14350 ( .Q(T14350_Q), .CK(T14347_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14349 ( .Q(T14349_Q), .CK(T14327_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14348 ( .Q(T14348_Q), .CK(T14389_Q), .D(T16255_Y));
KC_DFFHQ_X1 T14330 ( .Q(T14330_Q), .CK(T14153_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14329 ( .Q(T14329_Q), .CK(T14026_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14328 ( .Q(T14328_Q), .CK(T14026_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14320 ( .Q(T14320_Q), .CK(T14026_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14319 ( .Q(T14319_Q), .CK(T14154_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14306 ( .Q(T14306_Q), .CK(T14153_Q), .D(T9933_Y));
KC_DFFHQ_X1 T14305 ( .Q(T14305_Q), .CK(T14154_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14287 ( .Q(T14287_Q), .CK(T16467_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14286 ( .Q(T14286_Q), .CK(T14867_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14285 ( .Q(T14285_Q), .CK(T14028_Q), .D(T9943_Y));
KC_DFFHQ_X1 T14284 ( .Q(T14284_Q), .CK(T14154_Q), .D(T9954_Y));
KC_DFFHQ_X1 T14899 ( .Q(T14899_Q), .CK(T14389_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14898 ( .Q(T14898_Q), .CK(T14347_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14437 ( .Q(T14437_Q), .CK(T14327_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14436 ( .Q(T14436_Q), .CK(T14389_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14435 ( .Q(T14435_Q), .CK(T14327_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14434 ( .Q(T14434_Q), .CK(T14347_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14429 ( .Q(T14429_Q), .CK(T14327_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14428 ( .Q(T14428_Q), .CK(T14389_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14411 ( .Q(T14411_Q), .CK(T14347_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14410 ( .Q(T14410_Q), .CK(T14347_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14409 ( .Q(T14409_Q), .CK(T14389_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14408 ( .Q(T14408_Q), .CK(T14389_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14407 ( .Q(T14407_Q), .CK(T14347_Q), .D(T10186_Y));
KC_DFFHQ_X1 T14391 ( .Q(T14391_Q), .CK(T14327_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14390 ( .Q(T14390_Q), .CK(T14327_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14508 ( .Q(T14508_Q), .CK(T14944_Q), .D(T16206_Y));
KC_DFFHQ_X1 T14507 ( .Q(T14507_Q), .CK(T14944_Q), .D(T16205_Y));
KC_DFFHQ_X1 T14504 ( .Q(T14504_Q), .CK(T14347_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14503 ( .Q(T14503_Q), .CK(T14327_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14502 ( .Q(T14502_Q), .CK(T14389_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14483 ( .Q(T14483_Q), .CK(T14944_Q), .D(T16209_Y));
KC_DFFHQ_X1 T14482 ( .Q(T14482_Q), .CK(T14944_Q), .D(T16208_Y));
KC_DFFHQ_X1 T14467 ( .Q(T14467_Q), .CK(T14531_Q), .D(T16204_Y));
KC_DFFHQ_X1 T14459 ( .Q(T14459_Q), .CK(T14944_Q), .D(T16203_Y));
KC_DFFHQ_X1 T14942 ( .Q(T14942_Q), .CK(T14944_Q), .D(T5148_Y));
KC_DFFHQ_X1 T14523 ( .Q(T14523_Q), .CK(T14542_Q), .D(T4421_Y));
KC_DFFHQ_X1 T14551 ( .Q(T14551_Q), .CK(T14545_Q), .D(T11443_Y));
KC_DFFHQ_X1 T14550 ( .Q(T14550_Q), .CK(T14545_Q), .D(T12337_Y));
KC_DFFHQ_X1 T14549 ( .Q(T14549_Q), .CK(T14545_Q), .D(T11441_Y));
KC_DFFHQ_X1 T14548 ( .Q(T14548_Q), .CK(T14545_Q), .D(T11439_Y));
KC_DFFHQ_X1 T14547 ( .Q(T14547_Q), .CK(T14545_Q), .D(T4504_Y));
KC_DFFHQ_X1 T14584 ( .Q(T14584_Q), .CK(T13496_Q), .D(T15242_Y));
KC_DFFHQ_X1 T14717 ( .Q(T14717_Q), .CK(T13467_Q), .D(T15242_Y));
KC_DFFHQ_X1 T14713 ( .Q(T14713_Q), .CK(T13496_Q), .D(T15243_Y));
KC_DFFHQ_X1 T14675 ( .Q(T14675_Q), .CK(T14638_Q), .D(T10416_Y));
KC_DFFHQ_X1 T14673 ( .Q(T14673_Q), .CK(T14638_Q), .D(T15193_Y));
KC_DFFHQ_X1 T14649 ( .Q(T14649_Q), .CK(T14643_Q), .D(T9788_Y));
KC_DFFHQ_X1 T14731 ( .Q(T14731_Q), .CK(T13608_Q), .D(T15203_Y));
KC_DFFHQ_X1 T14715 ( .Q(T14715_Q), .CK(T14691_Q), .D(T15196_Y));
KC_DFFHQ_X1 T14714 ( .Q(T14714_Q), .CK(T14691_Q), .D(T9608_Y));
KC_DFFHQ_X1 T14711 ( .Q(T14711_Q), .CK(T14690_Q), .D(T15240_Y));
KC_DFFHQ_X1 T14710 ( .Q(T14710_Q), .CK(T14691_Q), .D(T15209_Y));
KC_DFFHQ_X1 T14674 ( .Q(T14674_Q), .CK(T13815_Q), .D(T10416_Y));
KC_DFFHQ_X1 T14650 ( .Q(T14650_Q), .CK(T13858_Q), .D(T9788_Y));
KC_DFFHQ_X1 T14646 ( .Q(T14646_Q), .CK(T14643_Q), .D(T9793_Y));
KC_DFFHQ_X1 T14644 ( .Q(T14644_Q), .CK(T13792_Q), .D(T9788_Y));
KC_DFFHQ_X1 T14729 ( .Q(T14729_Q), .CK(T14688_Q), .D(T15209_Y));
KC_DFFHQ_X1 T14712 ( .Q(T14712_Q), .CK(T14690_Q), .D(T10401_Y));
KC_DFFHQ_X1 T14709 ( .Q(T14709_Q), .CK(T14688_Q), .D(T10401_Y));
KC_DFFHQ_X1 T14707 ( .Q(T14707_Q), .CK(T14690_Q), .D(T15208_Y));
KC_DFFHQ_X1 T14640 ( .Q(T14640_Q), .CK(T14642_Q), .D(T9696_Y));
KC_DFFHQ_X1 T14639 ( .Q(T14639_Q), .CK(T14642_Q), .D(T9793_Y));
KC_DFFHQ_X1 T14624 ( .Q(T14624_Q), .CK(T14250_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14621 ( .Q(T14621_Q), .CK(T14224_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14620 ( .Q(T14620_Q), .CK(T14237_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14597 ( .Q(T14597_Q), .CK(T14212_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14727 ( .Q(T14727_Q), .CK(T1651_Y), .D(T12501_Y));
KC_DFFHQ_X1 T14726 ( .Q(T14726_Q), .CK(T1651_Y), .D(T12506_Y));
KC_DFFHQ_X1 T14720 ( .Q(T14720_Q), .CK(T1651_Y), .D(T12910_Y));
KC_DFFHQ_X1 T14706 ( .Q(T14706_Q), .CK(T13608_Q), .D(T15208_Y));
KC_DFFHQ_X1 T14663 ( .Q(T14663_Q), .CK(T13849_Q), .D(T9618_Y));
KC_DFFHQ_X1 T14662 ( .Q(T14662_Q), .CK(T1650_Y), .D(T12580_Y));
KC_DFFHQ_X1 T14634 ( .Q(T14634_Q), .CK(T14012_Q), .D(T10348_Y));
KC_DFFHQ_X1 T14633 ( .Q(T14633_Q), .CK(T13849_Q), .D(T10350_Y));
KC_DFFHQ_X1 T14616 ( .Q(T14616_Q), .CK(T1549_Y), .D(T12698_Y));
KC_DFFHQ_X1 T14596 ( .Q(T14596_Q), .CK(T14591_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14595 ( .Q(T14595_Q), .CK(T13329_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14592 ( .Q(T14592_Q), .CK(T14374_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14722 ( .Q(T14722_Q), .CK(T13492_Q), .D(T9687_Y));
KC_DFFHQ_X1 T14721 ( .Q(T14721_Q), .CK(T13491_Q), .D(T9606_Y));
KC_DFFHQ_X1 T14705 ( .Q(T14705_Q), .CK(T13445_Q), .D(T10444_Y));
KC_DFFHQ_X1 T14704 ( .Q(T14704_Q), .CK(T13745_Q), .D(T10444_Y));
KC_DFFHQ_X1 T14655 ( .Q(T14655_Q), .CK(T14009_Q), .D(T9609_Y));
KC_DFFHQ_X1 T14627 ( .Q(T14627_Q), .CK(T13951_Q), .D(T8533_Y));
KC_DFFHQ_X1 T14607 ( .Q(T14607_Q), .CK(T4900_Y), .D(T2544_Y));
KC_DFFHQ_X1 T14594 ( .Q(T14594_Q), .CK(T14374_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14593 ( .Q(T14593_Q), .CK(T14591_Q), .D(T15226_Y));
KC_DFFHQ_X1 T6461 ( .Q(T6461_Q), .CK(T13757_Q), .D(T9606_Y));
KC_DFFHQ_X1 T14789 ( .Q(T14789_Q), .CK(T13464_Q), .D(T10445_Y));
KC_DFFHQ_X1 T14773 ( .Q(T14773_Q), .CK(T1638_Y), .D(T11128_Y));
KC_DFFHQ_X1 T14656 ( .Q(T14656_Q), .CK(T14864_Q), .D(T6716_Y));
KC_DFFHQ_X1 T14861 ( .Q(T14861_Q), .CK(T14864_Q), .D(T9760_Y));
KC_DFFHQ_X1 T14860 ( .Q(T14860_Q), .CK(T14864_Q), .D(T9749_Y));
KC_DFFHQ_X1 T14840 ( .Q(T14840_Q), .CK(T1638_Y), .D(T11944_Y));
KC_DFFHQ_X1 T14788 ( .Q(T14788_Q), .CK(T13630_Q), .D(T9601_Y));
KC_DFFHQ_X1 T14787 ( .Q(T14787_Q), .CK(T14682_Q), .D(T9599_Y));
KC_DFFHQ_X1 T14786 ( .Q(T14786_Q), .CK(T13630_Q), .D(T9599_Y));
KC_DFFHQ_X1 T14785 ( .Q(T14785_Q), .CK(T13464_Q), .D(T9601_Y));
KC_DFFHQ_X1 T14768 ( .Q(T14768_Q), .CK(T13445_Q), .D(T9599_Y));
KC_DFFHQ_X1 T14884 ( .Q(T14884_Q), .CK(T5315_Y), .D(T12708_Y));
KC_DFFHQ_X1 T14857 ( .Q(T14857_Q), .CK(T5315_Y), .D(T12601_Y));
KC_DFFHQ_X1 T14839 ( .Q(T14839_Q), .CK(T2495_Y), .D(T11942_Y));
KC_DFFHQ_X1 T14836 ( .Q(T14836_Q), .CK(T2495_Y), .D(T11929_Y));
KC_DFFHQ_X1 T14782 ( .Q(T14782_Q), .CK(T13664_Q), .D(T9589_Y));
KC_DFFHQ_X1 T14765 ( .Q(T14765_Q), .CK(T2495_Y), .D(T12548_Y));
KC_DFFHQ_X1 T14951 ( .Q(T14951_Q), .CK(T14948_Q), .D(T11335_Y));
KC_DFFHQ_X1 T14950 ( .Q(T14950_Q), .CK(T3199_Y), .D(T3184_Y));
KC_DFFHQ_X1 T14883 ( .Q(T14883_Q), .CK(T14354_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14880 ( .Q(T14880_Q), .CK(T14353_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14879 ( .Q(T14879_Q), .CK(T14355_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14856 ( .Q(T14856_Q), .CK(T5315_Y), .D(T12936_Y));
KC_DFFHQ_X1 T14855 ( .Q(T14855_Q), .CK(T14079_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14837 ( .Q(T14837_Q), .CK(T14076_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14833 ( .Q(T14833_Q), .CK(T13926_Q), .D(T9741_Y));
KC_DFFHQ_X1 T14832 ( .Q(T14832_Q), .CK(T13927_Q), .D(T9844_Y));
KC_DFFHQ_X1 T14781 ( .Q(T14781_Q), .CK(T13663_Q), .D(T9593_Y));
KC_DFFHQ_X1 T14780 ( .Q(T14780_Q), .CK(T13644_Q), .D(T9593_Y));
KC_DFFHQ_X1 T14762 ( .Q(T14762_Q), .CK(T14775_Q), .D(T9644_Y));
KC_DFFHQ_X1 T14761 ( .Q(T14761_Q), .CK(T3026_Y), .D(T13205_Y));
KC_DFFHQ_X1 T14947 ( .Q(T14947_Q), .CK(T14948_Q), .D(T11979_Y));
KC_DFFHQ_X1 T14946 ( .Q(T14946_Q), .CK(T14531_Q), .D(T16225_Y));
KC_DFFHQ_X1 T14906 ( .Q(T14906_Q), .CK(T14393_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14902 ( .Q(T14902_Q), .CK(T14393_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14901 ( .Q(T14901_Q), .CK(T14944_Q), .D(T3777_Y));
KC_DFFHQ_X1 T14900 ( .Q(T14900_Q), .CK(T14406_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14878 ( .Q(T14878_Q), .CK(T14028_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14876 ( .Q(T14876_Q), .CK(T14867_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14875 ( .Q(T14875_Q), .CK(T14866_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14850 ( .Q(T14850_Q), .CK(T14036_Q), .D(T10492_Y));
KC_DFFHQ_X1 T14828 ( .Q(T14828_Q), .CK(T14062_Q), .D(T9733_Y));
KC_DFFHQ_X1 T14778 ( .Q(T14778_Q), .CK(T13644_Q), .D(T9591_Y));
KC_DFFHQ_X1 T14757 ( .Q(T14757_Q), .CK(T13633_Q), .D(T15252_Y));
KC_DFFHQ_X1 T14897 ( .Q(T14897_Q), .CK(T14389_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14896 ( .Q(T14896_Q), .CK(T14327_Q), .D(T10187_Y));
KC_DFFHQ_X1 T14895 ( .Q(T14895_Q), .CK(T14347_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14873 ( .Q(T14873_Q), .CK(T14154_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14872 ( .Q(T14872_Q), .CK(T14153_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14844 ( .Q(T14844_Q), .CK(T14843_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14825 ( .Q(T14825_Q), .CK(T14843_Q), .D(T9733_Y));
KC_DFFHQ_X1 T14824 ( .Q(T14824_Q), .CK(T14035_Q), .D(T9733_Y));
KC_DFFHQ_X1 T14777 ( .Q(T14777_Q), .CK(T13619_Q), .D(T9602_Y));
KC_DFFHQ_X1 T14776 ( .Q(T14776_Q), .CK(T13617_Q), .D(T9602_Y));
KC_DFFHQ_X1 T14812 ( .Q(T14812_Q), .CK(T13633_Q), .D(T6443_Y));
KC_DFFHQ_X1 T14587 ( .Q(T14587_Q), .CK(T13345_Q), .D(T15241_Y));
KC_DFFHQ_X1 T13429 ( .Q(T13429_Q), .CK(T13492_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13426 ( .Q(T13426_Q), .CK(T13644_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13421 ( .Q(T13421_Q), .CK(T13633_Q), .D(T15199_Y));
KC_DFFHQ_X1 T13415 ( .Q(T13415_Q), .CK(T13491_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13412 ( .Q(T13412_Q), .CK(T13667_Q), .D(T10454_Y));
KC_DFFHQ_X1 T13408 ( .Q(T13408_Q), .CK(T14791_Q), .D(T10456_Y));
KC_DFFHQ_X1 T13406 ( .Q(T13406_Q), .CK(T13665_Q), .D(T9587_Y));
KC_DFFHQ_X1 T13401 ( .Q(T13401_Q), .CK(T14702_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13395 ( .Q(T13395_Q), .CK(T13644_Q), .D(T10447_Y));
KC_DFFHQ_X1 T13393 ( .Q(T13393_Q), .CK(T14791_Q), .D(T10447_Y));
KC_DFFHQ_X1 T13385 ( .Q(T13385_Q), .CK(T13347_Q), .D(T15203_Y));
KC_DFFHQ_X1 T13373 ( .Q(T13373_Q), .CK(T13445_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13366 ( .Q(T13366_Q), .CK(T13376_Q), .D(T15203_Y));
KC_DFFHQ_X1 T13361 ( .Q(T13361_Q), .CK(T14677_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13358 ( .Q(T13358_Q), .CK(T13445_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13356 ( .Q(T13356_Q), .CK(T14678_Q), .D(T15236_Y));
KC_DFFHQ_X1 T13339 ( .Q(T13339_Q), .CK(T14683_Q), .D(T15250_Y));
KC_DFFHQ_X1 T13338 ( .Q(T13338_Q), .CK(T14678_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13336 ( .Q(T13336_Q), .CK(T14678_Q), .D(T15243_Y));
KC_DFFHQ_X1 T13335 ( .Q(T13335_Q), .CK(T13346_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13333 ( .Q(T13333_Q), .CK(T13346_Q), .D(T15243_Y));
KC_DFFHQ_X1 T14811 ( .Q(T14811_Q), .CK(T14682_Q), .D(T10445_Y));
KC_DFFHQ_X1 T14810 ( .Q(T14810_Q), .CK(T13630_Q), .D(T10445_Y));
KC_DFFHQ_X1 T14804 ( .Q(T14804_Q), .CK(T13464_Q), .D(T9600_Y));
KC_DFFHQ_X1 T14802 ( .Q(T14802_Q), .CK(T13663_Q), .D(T9589_Y));
KC_DFFHQ_X1 T14795 ( .Q(T14795_Q), .CK(T14791_Q), .D(T9591_Y));
KC_DFFHQ_X1 T14697 ( .Q(T14697_Q), .CK(T14689_Q), .D(T15208_Y));
KC_DFFHQ_X1 T14684 ( .Q(T14684_Q), .CK(T14683_Q), .D(T10445_Y));
KC_DFFHQ_X1 T14585 ( .Q(T14585_Q), .CK(T13496_Q), .D(T15210_Y));
KC_DFFHQ_X1 T13552 ( .Q(T13552_Q), .CK(T14791_Q), .D(T9589_Y));
KC_DFFHQ_X1 T13549 ( .Q(T13549_Q), .CK(T13619_Q), .D(T6443_Y));
KC_DFFHQ_X1 T13541 ( .Q(T13541_Q), .CK(T13617_Q), .D(T6443_Y));
KC_DFFHQ_X1 T13538 ( .Q(T13538_Q), .CK(T13630_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13532 ( .Q(T13532_Q), .CK(T13642_Q), .D(T10448_Y));
KC_DFFHQ_X1 T13529 ( .Q(T13529_Q), .CK(T13621_Q), .D(T9588_Y));
KC_DFFHQ_X1 T13527 ( .Q(T13527_Q), .CK(T13644_Q), .D(T9589_Y));
KC_DFFHQ_X1 T13523 ( .Q(T13523_Q), .CK(T13620_Q), .D(T6443_Y));
KC_DFFHQ_X1 T13517 ( .Q(T13517_Q), .CK(T14682_Q), .D(T10455_Y));
KC_DFFHQ_X1 T13510 ( .Q(T13510_Q), .CK(T13682_Q), .D(T10446_Y));
KC_DFFHQ_X1 T13504 ( .Q(T13504_Q), .CK(T13666_Q), .D(T6443_Y));
KC_DFFHQ_X1 T13502 ( .Q(T13502_Q), .CK(T13497_Q), .D(T15203_Y));
KC_DFFHQ_X1 T13482 ( .Q(T13482_Q), .CK(T14689_Q), .D(T10394_Y));
KC_DFFHQ_X1 T13474 ( .Q(T13474_Q), .CK(T13757_Q), .D(T15200_Y));
KC_DFFHQ_X1 T13470 ( .Q(T13470_Q), .CK(T13478_Q), .D(T15236_Y));
KC_DFFHQ_X1 T13459 ( .Q(T13459_Q), .CK(T13467_Q), .D(T15236_Y));
KC_DFFHQ_X1 T13452 ( .Q(T13452_Q), .CK(T13466_Q), .D(T10394_Y));
KC_DFFHQ_X1 T13442 ( .Q(T13442_Q), .CK(T14767_Q), .D(T15249_Y));
KC_DFFHQ_X1 T13441 ( .Q(T13441_Q), .CK(T13467_Q), .D(T15241_Y));
KC_DFFHQ_X1 T13439 ( .Q(T13439_Q), .CK(T13467_Q), .D(T15243_Y));
KC_DFFHQ_X1 T13437 ( .Q(T13437_Q), .CK(T13448_Q), .D(T15243_Y));
KC_DFFHQ_X1 T13434 ( .Q(T13434_Q), .CK(T13345_Q), .D(T15210_Y));
KC_DFFHQ_X1 T14770 ( .Q(T14770_Q), .CK(T13745_Q), .D(T9601_Y));
KC_DFFHQ_X1 T14733 ( .Q(T14733_Q), .CK(T14690_Q), .D(T9608_Y));
KC_DFFHQ_X1 T14718 ( .Q(T14718_Q), .CK(T13682_Q), .D(T9606_Y));
KC_DFFHQ_X1 T13678 ( .Q(T13678_Q), .CK(T13490_Q), .D(T9600_Y));
KC_DFFHQ_X1 T13675 ( .Q(T13675_Q), .CK(T13667_Q), .D(T9593_Y));
KC_DFFHQ_X1 T13670 ( .Q(T13670_Q), .CK(T13617_Q), .D(T15252_Y));
KC_DFFHQ_X1 T13661 ( .Q(T13661_Q), .CK(T13445_Q), .D(T9601_Y));
KC_DFFHQ_X1 T13655 ( .Q(T13655_Q), .CK(T4977_Y), .D(T11925_Y));
KC_DFFHQ_X1 T13652 ( .Q(T13652_Q), .CK(T13617_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13647 ( .Q(T13647_Q), .CK(T13645_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13643 ( .Q(T13643_Q), .CK(T14683_Q), .D(T9601_Y));
KC_DFFHQ_X1 T13638 ( .Q(T13638_Q), .CK(T13620_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13628 ( .Q(T13628_Q), .CK(T13446_Q), .D(T9600_Y));
KC_DFFHQ_X1 T13627 ( .Q(T13627_Q), .CK(T14767_Q), .D(T9600_Y));
KC_DFFHQ_X1 T13625 ( .Q(T13625_Q), .CK(T13664_Q), .D(T9592_Y));
KC_DFFHQ_X1 T13622 ( .Q(T13622_Q), .CK(T13618_Q), .D(T9602_Y));
KC_DFFHQ_X1 T13613 ( .Q(T13613_Q), .CK(T14691_Q), .D(T15203_Y));
KC_DFFHQ_X1 T13609 ( .Q(T13609_Q), .CK(T1651_Y), .D(T12513_Y));
KC_DFFHQ_X1 T13603 ( .Q(T13603_Q), .CK(T1651_Y), .D(T12511_Y));
KC_DFFHQ_X1 T13602 ( .Q(T13602_Q), .CK(T14703_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13595 ( .Q(T13595_Q), .CK(T14703_Q), .D(T9687_Y));
KC_DFFHQ_X1 T13591 ( .Q(T13591_Q), .CK(T14690_Q), .D(T15196_Y));
KC_DFFHQ_X1 T13586 ( .Q(T13586_Q), .CK(T1651_Y), .D(T12499_Y));
KC_DFFHQ_X1 T13579 ( .Q(T13579_Q), .CK(T13682_Q), .D(T9687_Y));
KC_DFFHQ_X1 T13576 ( .Q(T13576_Q), .CK(T13466_Q), .D(T9608_Y));
KC_DFFHQ_X1 T13573 ( .Q(T13573_Q), .CK(T1651_Y), .D(T12505_Y));
KC_DFFHQ_X1 T13571 ( .Q(T13571_Q), .CK(T13340_Q), .D(T9605_Y));
KC_DFFHQ_X1 T13569 ( .Q(T13569_Q), .CK(T13496_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13568 ( .Q(T13568_Q), .CK(T13478_Q), .D(T15239_Y));
KC_DFFHQ_X1 T13566 ( .Q(T13566_Q), .CK(T13478_Q), .D(T15238_Y));
KC_DFFHQ_X1 T13564 ( .Q(T13564_Q), .CK(T13495_Q), .D(T15242_Y));
KC_DFFHQ_X1 T14940 ( .Q(T14940_Q), .CK(T1638_Y), .D(T11957_Y));
KC_DFFHQ_X1 T14930 ( .Q(T14930_Q), .CK(T2495_Y), .D(T12999_Y));
KC_DFFHQ_X1 T14927 ( .Q(T14927_Q), .CK(T13618_Q), .D(T15252_Y));
KC_DFFHQ_X1 T14923 ( .Q(T14923_Q), .CK(T13926_Q), .D(T9742_Y));
KC_DFFHQ_X1 T14921 ( .Q(T14921_Q), .CK(T14843_Q), .D(T9727_Y));
KC_DFFHQ_X1 T14917 ( .Q(T14917_Q), .CK(T14843_Q), .D(T9734_Y));
KC_DFFHQ_X1 T14754 ( .Q(T14754_Q), .CK(T14665_Q), .D(T15206_Y));
KC_DFFHQ_X1 T14752 ( .Q(T14752_Q), .CK(T14745_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13777 ( .Q(T13777_Q), .CK(T1638_Y), .D(T11129_Y));
KC_DFFHQ_X1 T13771 ( .Q(T13771_Q), .CK(T4977_Y), .D(T11111_Y));
KC_DFFHQ_X1 T13768 ( .Q(T13768_Q), .CK(T13618_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13766 ( .Q(T13766_Q), .CK(T13618_Q), .D(T9644_Y));
KC_DFFHQ_X1 T13763 ( .Q(T13763_Q), .CK(T13665_Q), .D(T9648_Y));
KC_DFFHQ_X1 T13756 ( .Q(T13756_Q), .CK(T13618_Q), .D(T8522_Y));
KC_DFFHQ_X1 T13753 ( .Q(T13753_Q), .CK(T13633_Q), .D(T9644_Y));
KC_DFFHQ_X1 T13742 ( .Q(T13742_Q), .CK(T14688_Q), .D(T15203_Y));
KC_DFFHQ_X1 T13738 ( .Q(T13738_Q), .CK(T14665_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13715 ( .Q(T13715_Q), .CK(T13939_Q), .D(T9618_Y));
KC_DFFHQ_X1 T13712 ( .Q(T13712_Q), .CK(T13938_Q), .D(T9618_Y));
KC_DFFHQ_X1 T13703 ( .Q(T13703_Q), .CK(T14665_Q), .D(T10416_Y));
KC_DFFHQ_X1 T13700 ( .Q(T13700_Q), .CK(T13719_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13698 ( .Q(T13698_Q), .CK(T14666_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13688 ( .Q(T13688_Q), .CK(T13939_Q), .D(T10351_Y));
KC_DFFHQ_X1 T14862 ( .Q(T14862_Q), .CK(T13952_Q), .D(T9758_Y));
KC_DFFHQ_X1 T14851 ( .Q(T14851_Q), .CK(T14040_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14830 ( .Q(T14830_Q), .CK(T14067_Q), .D(T9741_Y));
KC_DFFHQ_X1 T14668 ( .Q(T14668_Q), .CK(T14664_Q), .D(T10417_Y));
KC_DFFHQ_X1 T14657 ( .Q(T14657_Q), .CK(T13849_Q), .D(T9617_Y));
KC_DFFHQ_X1 T14648 ( .Q(T14648_Q), .CK(T14637_Q), .D(T9793_Y));
KC_DFFHQ_X1 T14632 ( .Q(T14632_Q), .CK(T13804_Q), .D(T10350_Y));
KC_DFFHQ_X1 T14628 ( .Q(T14628_Q), .CK(T13952_Q), .D(T9757_Y));
KC_DFFHQ_X1 T13930 ( .Q(T13930_Q), .CK(T14864_Q), .D(T9759_Y));
KC_DFFHQ_X1 T13923 ( .Q(T13923_Q), .CK(T13937_Q), .D(T8533_Y));
KC_DFFHQ_X1 T13915 ( .Q(T13915_Q), .CK(T14865_Q), .D(T9749_Y));
KC_DFFHQ_X1 T13914 ( .Q(T13914_Q), .CK(T13937_Q), .D(T9749_Y));
KC_DFFHQ_X1 T13907 ( .Q(T13907_Q), .CK(T14040_Q), .D(T125_Q));
KC_DFFHQ_X1 T13905 ( .Q(T13905_Q), .CK(T14040_Q), .D(T9735_Y));
KC_DFFHQ_X1 T13898 ( .Q(T13898_Q), .CK(T13937_Q), .D(T6716_Y));
KC_DFFHQ_X1 T13886 ( .Q(T13886_Q), .CK(T13937_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13883 ( .Q(T13883_Q), .CK(T13950_Q), .D(T9759_Y));
KC_DFFHQ_X1 T13877 ( .Q(T13877_Q), .CK(T14035_Q), .D(T10492_Y));
KC_DFFHQ_X1 T13870 ( .Q(T13870_Q), .CK(T14637_Q), .D(T9803_Y));
KC_DFFHQ_X1 T13866 ( .Q(T13866_Q), .CK(T14637_Q), .D(T9789_Y));
KC_DFFHQ_X1 T13864 ( .Q(T13864_Q), .CK(T13858_Q), .D(T9793_Y));
KC_DFFHQ_X1 T13862 ( .Q(T13862_Q), .CK(T13793_Q), .D(T9793_Y));
KC_DFFHQ_X1 T13844 ( .Q(T13844_Q), .CK(T14625_Q), .D(T9757_Y));
KC_DFFHQ_X1 T13838 ( .Q(T13838_Q), .CK(T13815_Q), .D(T10417_Y));
KC_DFFHQ_X1 T13831 ( .Q(T13831_Q), .CK(T14745_Q), .D(T9699_Y));
KC_DFFHQ_X1 T13824 ( .Q(T13824_Q), .CK(T14659_Q), .D(T9698_Y));
KC_DFFHQ_X1 T13822 ( .Q(T13822_Q), .CK(T13792_Q), .D(T9793_Y));
KC_DFFHQ_X1 T13807 ( .Q(T13807_Q), .CK(T13849_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13806 ( .Q(T13806_Q), .CK(T13957_Q), .D(T10349_Y));
KC_DFFHQ_X1 T13801 ( .Q(T13801_Q), .CK(T13953_Q), .D(T6716_Y));
KC_DFFHQ_X1 T13798 ( .Q(T13798_Q), .CK(T13953_Q), .D(T8533_Y));
KC_DFFHQ_X1 T13794 ( .Q(T13794_Q), .CK(T13856_Q), .D(T9793_Y));
KC_DFFHQ_X1 T13788 ( .Q(T13788_Q), .CK(T14012_Q), .D(T10349_Y));
KC_DFFHQ_X1 T14092 ( .Q(T14092_Q), .CK(T14346_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14088 ( .Q(T14088_Q), .CK(T16467_Q), .D(T9826_Y));
KC_DFFHQ_X1 T14071 ( .Q(T14071_Q), .CK(T14008_Q), .D(T9760_Y));
KC_DFFHQ_X1 T14059 ( .Q(T14059_Q), .CK(T13951_Q), .D(T9760_Y));
KC_DFFHQ_X1 T14051 ( .Q(T14051_Q), .CK(T5315_Y), .D(T12650_Y));
KC_DFFHQ_X1 T14048 ( .Q(T14048_Q), .CK(T14078_Q), .D(T9740_Y));
KC_DFFHQ_X1 T14042 ( .Q(T14042_Q), .CK(T14035_Q), .D(T9852_Y));
KC_DFFHQ_X1 T14019 ( .Q(T14019_Q), .CK(T13792_Q), .D(T9812_Y));
KC_DFFHQ_X1 T14007 ( .Q(T14007_Q), .CK(T14637_Q), .D(T9788_Y));
KC_DFFHQ_X1 T14004 ( .Q(T14004_Q), .CK(T14637_Q), .D(T9811_Y));
KC_DFFHQ_X1 T14002 ( .Q(T14002_Q), .CK(T14643_Q), .D(T9812_Y));
KC_DFFHQ_X1 T13992 ( .Q(T13992_Q), .CK(T14009_Q), .D(T10350_Y));
KC_DFFHQ_X1 T13989 ( .Q(T13989_Q), .CK(T14008_Q), .D(T9757_Y));
KC_DFFHQ_X1 T13984 ( .Q(T13984_Q), .CK(T13953_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13982 ( .Q(T13982_Q), .CK(T14637_Q), .D(T9812_Y));
KC_DFFHQ_X1 T13972 ( .Q(T13972_Q), .CK(T14008_Q), .D(T9808_Y));
KC_DFFHQ_X1 T13970 ( .Q(T13970_Q), .CK(T13793_Q), .D(T9812_Y));
KC_DFFHQ_X1 T13965 ( .Q(T13965_Q), .CK(T13856_Q), .D(T9812_Y));
KC_DFFHQ_X1 T13956 ( .Q(T13956_Q), .CK(T13957_Q), .D(T10409_Y));
KC_DFFHQ_X1 T13949 ( .Q(T13949_Q), .CK(T13791_Q), .D(T9812_Y));
KC_DFFHQ_X1 T15072 ( .Q(T15072_Q), .CK(T3122_Y), .D(T12715_Y));
KC_DFFHQ_X1 T15068 ( .Q(T15068_Q), .CK(T14212_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14892 ( .Q(T14892_Q), .CK(T3122_Y), .D(T12718_Y));
KC_DFFHQ_X1 T14891 ( .Q(T14891_Q), .CK(T14346_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14881 ( .Q(T14881_Q), .CK(T5315_Y), .D(T13210_Y));
KC_DFFHQ_X1 T14622 ( .Q(T14622_Q), .CK(T14276_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14608 ( .Q(T14608_Q), .CK(T4900_Y), .D(T12695_Y));
KC_DFFHQ_X1 T14606 ( .Q(T14606_Q), .CK(T14212_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14604 ( .Q(T14604_Q), .CK(T14276_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14599 ( .Q(T14599_Q), .CK(T14253_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14195 ( .Q(T14195_Q), .CK(T14333_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14182 ( .Q(T14182_Q), .CK(T14333_Q), .D(T10508_Y));
KC_DFFHQ_X1 T14179 ( .Q(T14179_Q), .CK(T14866_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14170 ( .Q(T14170_Q), .CK(T14333_Q), .D(T9879_Y));
KC_DFFHQ_X1 T14167 ( .Q(T14167_Q), .CK(T14346_Q), .D(T9939_Y));
KC_DFFHQ_X1 T14164 ( .Q(T14164_Q), .CK(T14084_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14162 ( .Q(T14162_Q), .CK(T14025_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14152 ( .Q(T14152_Q), .CK(T3122_Y), .D(T13027_Y));
KC_DFFHQ_X1 T14140 ( .Q(T14140_Q), .CK(T16467_Q), .D(T9875_Y));
KC_DFFHQ_X1 T14136 ( .Q(T14136_Q), .CK(T14255_Q), .D(T10323_Y));
KC_DFFHQ_X1 T14134 ( .Q(T14134_Q), .CK(T14252_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14123 ( .Q(T14123_Q), .CK(T14255_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14121 ( .Q(T14121_Q), .CK(T14209_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14119 ( .Q(T14119_Q), .CK(T14252_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14114 ( .Q(T14114_Q), .CK(T14210_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14107 ( .Q(T14107_Q), .CK(T14250_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14101 ( .Q(T14101_Q), .CK(T14251_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14366 ( .Q(T14366_Q), .CK(T2047_Y), .D(T13047_Y));
KC_DFFHQ_X1 T14363 ( .Q(T14363_Q), .CK(T2047_Y), .D(T12747_Y));
KC_DFFHQ_X1 T14361 ( .Q(T14361_Q), .CK(T14354_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14345 ( .Q(T14345_Q), .CK(T2047_Y), .D(T13046_Y));
KC_DFFHQ_X1 T14342 ( .Q(T14342_Q), .CK(T2047_Y), .D(T12744_Y));
KC_DFFHQ_X1 T14340 ( .Q(T14340_Q), .CK(T14346_Q), .D(T16260_Y));
KC_DFFHQ_X1 T14338 ( .Q(T14338_Q), .CK(T14331_Q), .D(T10181_Y));
KC_DFFHQ_X1 T14325 ( .Q(T14325_Q), .CK(T14346_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14314 ( .Q(T14314_Q), .CK(T14333_Q), .D(T10087_Y));
KC_DFFHQ_X1 T14311 ( .Q(T14311_Q), .CK(T14867_Q), .D(T9953_Y));
KC_DFFHQ_X1 T14303 ( .Q(T14303_Q), .CK(T3122_Y), .D(T12732_Y));
KC_DFFHQ_X1 T14301 ( .Q(T14301_Q), .CK(T14333_Q), .D(T9964_Y));
KC_DFFHQ_X1 T14297 ( .Q(T14297_Q), .CK(T14333_Q), .D(T10055_Y));
KC_DFFHQ_X1 T14294 ( .Q(T14294_Q), .CK(T14028_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14290 ( .Q(T14290_Q), .CK(T14866_Q), .D(T9962_Y));
KC_DFFHQ_X1 T14283 ( .Q(T14283_Q), .CK(T14209_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14280 ( .Q(T14280_Q), .CK(T14212_Q), .D(T9910_Y));
KC_DFFHQ_X1 T14274 ( .Q(T14274_Q), .CK(T14255_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14266 ( .Q(T14266_Q), .CK(T14236_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14264 ( .Q(T14264_Q), .CK(T14236_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14263 ( .Q(T14263_Q), .CK(T14276_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14260 ( .Q(T14260_Q), .CK(T14212_Q), .D(T9912_Y));
KC_DFFHQ_X1 T14254 ( .Q(T14254_Q), .CK(T14237_Q), .D(T9911_Y));
KC_DFFHQ_X1 T14249 ( .Q(T14249_Q), .CK(T14236_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14244 ( .Q(T14244_Q), .CK(T14270_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14242 ( .Q(T14242_Q), .CK(T14236_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14241 ( .Q(T14241_Q), .CK(T14252_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14232 ( .Q(T14232_Q), .CK(T14225_Q), .D(T15227_Y));
KC_DFFHQ_X1 T14231 ( .Q(T14231_Q), .CK(T14255_Q), .D(T9888_Y));
KC_DFFHQ_X1 T14219 ( .Q(T14219_Q), .CK(T14251_Q), .D(T9907_Y));
KC_DFFHQ_X1 T14218 ( .Q(T14218_Q), .CK(T14236_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14215 ( .Q(T14215_Q), .CK(T14276_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14908 ( .Q(T14908_Q), .CK(T14405_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14904 ( .Q(T14904_Q), .CK(T14393_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14448 ( .Q(T14448_Q), .CK(T14406_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14445 ( .Q(T14445_Q), .CK(T14394_Q), .D(T5949_Y));
KC_DFFHQ_X1 T14440 ( .Q(T14440_Q), .CK(T14405_Q), .D(T10193_Y));
KC_DFFHQ_X1 T14438 ( .Q(T14438_Q), .CK(T14405_Q), .D(T5970_Y));
KC_DFFHQ_X1 T14422 ( .Q(T14422_Q), .CK(T14412_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14416 ( .Q(T14416_Q), .CK(T14405_Q), .D(T10182_Y));
KC_DFFHQ_X1 T14398 ( .Q(T14398_Q), .CK(T14406_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14397 ( .Q(T14397_Q), .CK(T14392_Q), .D(T5948_Y));
KC_DFFHQ_X1 T14388 ( .Q(T14388_Q), .CK(T14211_Q), .D(T10325_Y));
KC_DFFHQ_X1 T14522 ( .Q(T14522_Q), .CK(T3199_Y), .D(T12119_Y));
KC_DFFHQ_X1 T14517 ( .Q(T14517_Q), .CK(T14519_Q), .D(T11332_Y));
KC_DFFHQ_X1 T14511 ( .Q(T14511_Q), .CK(T14531_Q), .D(T16227_Y));
KC_DFFHQ_X1 T14493 ( .Q(T14493_Q), .CK(T3199_Y), .D(T12781_Y));
KC_DFFHQ_X1 T14492 ( .Q(T14492_Q), .CK(T3198_Y), .D(T12782_Y));
KC_DFFHQ_X1 T14488 ( .Q(T14488_Q), .CK(T14531_Q), .D(T16220_Y));
KC_DFFHQ_X1 T14484 ( .Q(T14484_Q), .CK(T14531_Q), .D(T3778_Y));
KC_DFFHQ_X1 T14480 ( .Q(T14480_Q), .CK(T3199_Y), .D(T12117_Y));
KC_DFFHQ_X1 T14475 ( .Q(T14475_Q), .CK(T3198_Y), .D(T12777_Y));
KC_DFFHQ_X1 T14472 ( .Q(T14472_Q), .CK(T14531_Q), .D(T16219_Y));
KC_DFFHQ_X1 T14466 ( .Q(T14466_Q), .CK(T14531_Q), .D(T16207_Y));
KC_DFFHQ_X1 T14465 ( .Q(T14465_Q), .CK(T3199_Y), .D(T12118_Y));
KC_DFFHQ_X1 T14461 ( .Q(T14461_Q), .CK(T14531_Q), .D(T16213_Y));
KC_DFFHQ_X1 T14455 ( .Q(T14455_Q), .CK(T13329_Q), .D(T9906_Y));
KC_DFFHQ_X1 T14454 ( .Q(T14454_Q), .CK(T13329_Q), .D(T15226_Y));
KC_DFFHQ_X1 T14453 ( .Q(T14453_Q), .CK(T13329_Q), .D(T9903_Y));
KC_DFFHQ_X1 T14536 ( .Q(T14536_Q), .CK(T14532_Q), .D(T2685_Y));
KC_DFFHQ_X1 T14526 ( .Q(T14526_Q), .CK(T14532_Q), .D(T2690_Y));
KC_DFFHQ_X1 T14546 ( .Q(T14546_Q), .CK(T14539_Q), .D(T12168_Y));
KC_DFFHQ_X1 T14544 ( .Q(T14544_Q), .CK(T14539_Q), .D(T11411_Y));
KC_DFFHQ_X1 T14540 ( .Q(T14540_Q), .CK(T14539_Q), .D(T11395_Y));
KC_DFFHQ_X1 T14952 ( .Q(T14952_Q), .CK(T14519_Q), .D(T11986_Y));
KC_DFFHQ_X1 T14943 ( .Q(T14943_Q), .CK(T14531_Q), .D(T16222_Y));
KC_DFFHQ_X1 T14894 ( .Q(T14894_Q), .CK(T14944_Q), .D(T3776_Y));
KC_DFFHQ_X1 T14877 ( .Q(T14877_Q), .CK(T14028_Q), .D(T9876_Y));
KC_DFFHQ_X1 T14853 ( .Q(T14853_Q), .CK(T14031_Q), .D(T9740_Y));
KC_DFFHQ_X1 T14845 ( .Q(T14845_Q), .CK(T14061_Q), .D(T10491_Y));
KC_DFFHQ_X1 T14834 ( .Q(T14834_Q), .CK(T14067_Q), .D(T9844_Y));
KC_DFFHQ_X1 T14784 ( .Q(T14784_Q), .CK(T13464_Q), .D(T9599_Y));
KC_DFFHQ_X1 T14783 ( .Q(T14783_Q), .CK(T13621_Q), .D(T9589_Y));
KC_DFFHQ_X1 T14779 ( .Q(T14779_Q), .CK(T13666_Q), .D(T9602_Y));
KC_DFFHQ_X1 T14769 ( .Q(T14769_Q), .CK(T1638_Y), .D(T11134_Y));
KC_DFFHQ_X1 T14766 ( .Q(T14766_Q), .CK(T3026_Y), .D(T12923_Y));
KC_DFFHQ_X1 T14763 ( .Q(T14763_Q), .CK(T14775_Q), .D(T8522_Y));
KC_DFFHQ_X1 T14756 ( .Q(T14756_Q), .CK(T13665_Q), .D(T9644_Y));
KC_DFFHQ_X1 T14730 ( .Q(T14730_Q), .CK(T14688_Q), .D(T9608_Y));
KC_DFFHQ_X1 T14725 ( .Q(T14725_Q), .CK(T1651_Y), .D(T12500_Y));
KC_DFFHQ_X1 T14716 ( .Q(T14716_Q), .CK(T13496_Q), .D(T15241_Y));
KC_DFFHQ_X1 T14708 ( .Q(T14708_Q), .CK(T14688_Q), .D(T15208_Y));
KC_DFFHQ_X1 T14645 ( .Q(T14645_Q), .CK(T14642_Q), .D(T9812_Y));
KC_DFFHQ_X1 T14626 ( .Q(T14626_Q), .CK(T13951_Q), .D(T9757_Y));
KC_DFFHQ_X1 T14623 ( .Q(T14623_Q), .CK(T14276_Q), .D(T10324_Y));
KC_DFFHQ_X1 T14615 ( .Q(T14615_Q), .CK(T1549_Y), .D(T12896_Y));
KC_DFFHQ_X1 T14612 ( .Q(T14612_Q), .CK(T4900_Y), .D(T12691_Y));
KC_DFFHQ_X1 T14598 ( .Q(T14598_Q), .CK(T14211_Q), .D(T9913_Y));
KC_DFFHQ_X1 T14590 ( .Q(T14590_Q), .CK(T13329_Q), .D(T15225_Y));
KC_DFFHQ_X1 T14583 ( .Q(T14583_Q), .CK(T13467_Q), .D(T15210_Y));
KC_OAI22_X1 T13284 ( .A1(T12443_Y), .B0(T921_Y), .B1(T229_Y),     .A0(T8784_Y), .Y(T13284_Y));
KC_OAI22_X1 T13283 ( .A1(T9388_Y), .B0(T924_Y), .B1(T7670_Y),     .A0(T7569_Y), .Y(T13283_Y));
KC_OAI22_X1 T13282 ( .A1(T7576_Y), .B0(T15655_Y), .B1(T8780_Y),     .A0(T9379_Y), .Y(T13282_Y));
KC_OAI22_X1 T13246 ( .A1(T12450_Y), .B0(T8907_Y), .B1(T936_Y),     .A0(T968_Y), .Y(T13246_Y));
KC_OAI22_X1 T13240 ( .A1(T7828_Y), .B0(T917_Y), .B1(T7823_Y),     .A0(T7688_Y), .Y(T13240_Y));
KC_OAI22_X1 T13256 ( .A1(T7917_Y), .B0(T1206_Y), .B1(T7918_Y),     .A0(T7902_Y), .Y(T13256_Y));
KC_OAI22_X1 T13254 ( .A1(T8103_Y), .B0(T1273_Y), .B1(T8139_Y),     .A0(T16391_Y), .Y(T13254_Y));
KC_OAI22_X1 T13253 ( .A1(T7909_Y), .B0(T1321_Y), .B1(T8872_Y),     .A0(T8916_Y), .Y(T13253_Y));
KC_OAI22_X1 T13238 ( .A1(T7658_Y), .B0(T8754_Y), .B1(T740_Y),     .A0(T742_Y), .Y(T13238_Y));
KC_OAI22_X1 T13281 ( .A1(T7816_Y), .B0(T7827_Y), .B1(T12607_Y),     .A0(T7564_Y), .Y(T13281_Y));
KC_OAI22_X1 T13255 ( .A1(T8101_Y), .B0(T8078_Y), .B1(T12886_Y),     .A0(T7905_Y), .Y(T13255_Y));
KC_OAI22_X1 T13265 ( .A1(T614_Y), .B0(T168_Y), .B1(T15538_Y),     .A0(T561_Q), .Y(T13265_Y));
KC_OAI22_X1 T13217 ( .A1(T15331_Y), .B0(T5194_Q), .B1(T108_Y),     .A0(T621_Q), .Y(T13217_Y));
KC_OAI22_X1 T13270 ( .A1(T15355_Y), .B0(T450_Q), .B1(T6313_Y),     .A0(T812_Q), .Y(T13270_Y));
KC_OAI22_X1 T13220 ( .A1(T15171_Y), .B0(T5223_Q), .B1(T249_Y),     .A0(T649_Q), .Y(T13220_Y));
KC_OAI22_X1 T13219 ( .A1(T6289_Y), .B0(T5227_Q), .B1(T304_Y),     .A0(T817_Q), .Y(T13219_Y));
KC_OAI22_X1 T13218 ( .A1(T15349_Y), .B0(T446_Q), .B1(T250_Y),     .A0(T5229_Q), .Y(T13218_Y));
KC_OAI22_X1 T13269 ( .A1(T6288_Y), .B0(T445_Q), .B1(T6264_Y),     .A0(T847_Q), .Y(T13269_Y));
KC_OAI22_X1 T13226 ( .A1(T333_Y), .B0(T4845_Q), .B1(T6332_Y),     .A0(T653_Q), .Y(T13226_Y));
KC_OAI22_X1 T13221 ( .A1(T345_Y), .B0(T5240_Q), .B1(T6266_Y),     .A0(T843_Q), .Y(T13221_Y));
KC_OAI22_X1 T13232 ( .A1(T12395_Y), .B0(T6485_Y), .B1(T557_Y),     .A0(T12395_Y), .Y(T13232_Y));
KC_OAI22_X1 T13249 ( .A1(T15842_Y), .B0(T8895_Y), .B1(T7892_Y),     .A0(T8899_Y), .Y(T13249_Y));
KC_OAI22_X1 T13248 ( .A1(T15842_Y), .B0(T8894_Y), .B1(T7892_Y),     .A0(T8898_Y), .Y(T13248_Y));
KC_OAI22_X1 T13247 ( .A1(T15842_Y), .B0(T13260_Y), .B1(T7892_Y),     .A0(T9445_Y), .Y(T13247_Y));
KC_OAI22_X1 T13245 ( .A1(T15842_Y), .B0(T8939_Y), .B1(T7892_Y),     .A0(T8942_Y), .Y(T13245_Y));
KC_OAI22_X1 T13244 ( .A1(T15842_Y), .B0(T9411_Y), .B1(T7892_Y),     .A0(T9415_Y), .Y(T13244_Y));
KC_OAI22_X1 T13243 ( .A1(T15842_Y), .B0(T8803_Y), .B1(T7892_Y),     .A0(T9407_Y), .Y(T13243_Y));
KC_OAI22_X1 T13242 ( .A1(T15842_Y), .B0(T9001_Y), .B1(T7892_Y),     .A0(T9010_Y), .Y(T13242_Y));
KC_OAI22_X1 T13250 ( .A1(T1327_Y), .B0(T1255_Y), .B1(T16387_Y),     .A0(T8034_Y), .Y(T13250_Y));
KC_OAI22_X1 T13287 ( .A1(T6625_Y), .B0(T15740_Y), .B1(T10918_Y),     .A0(T9331_Y), .Y(T13287_Y));
KC_OAI22_X1 T13286 ( .A1(T6638_Y), .B0(T896_Y), .B1(T10918_Y),     .A0(T7410_Y), .Y(T13286_Y));
KC_OAI22_X1 T13285 ( .A1(T6630_Y), .B0(T9318_Y), .B1(T10918_Y),     .A0(T7413_Y), .Y(T13285_Y));
KC_OAI22_X1 T13274 ( .A1(T15659_Y), .B0(T124_Q), .B1(T10918_Y),     .A0(T7590_Y), .Y(T13274_Y));
KC_OAI22_X1 T13272 ( .A1(T6700_Y), .B0(T9316_Y), .B1(T10918_Y),     .A0(T7412_Y), .Y(T13272_Y));
KC_OAI22_X1 T13233 ( .A1(T9306_Y), .B0(T7410_Y), .B1(T15406_Y),     .A0(T8655_Y), .Y(T13233_Y));
KC_OAI22_X1 T13239 ( .A1(T12422_Y), .B0(T15654_Y), .B1(T783_Y),     .A0(T7839_Y), .Y(T13239_Y));
KC_OAI22_X1 T13237 ( .A1(T7617_Y), .B0(T7618_Y), .B1(T659_Y),     .A0(T7611_Y), .Y(T13237_Y));
KC_OAI22_X1 T13276 ( .A1(T16381_Y), .B0(T7868_Y), .B1(T7869_Y),     .A0(T16380_Y), .Y(T13276_Y));
KC_OAI22_X1 T13257 ( .A1(T8112_Y), .B0(T9000_Y), .B1(T8995_Y),     .A0(T961_Y), .Y(T13257_Y));
KC_OAI22_X1 T13201 ( .A1(T7977_Y), .B0(T1008_Y), .B1(T10047_Y),     .A0(T10316_Y), .Y(T13201_Y));
KC_OAI22_X1 T13200 ( .A1(T10043_Y), .B0(T7998_Y), .B1(T10316_Y),     .A0(T987_Y), .Y(T13200_Y));
KC_OAI22_X1 T13023 ( .A1(T7999_Y), .B0(T16394_Y), .B1(T10317_Y),     .A0(T10316_Y), .Y(T13023_Y));
KC_OAI22_X1 T13022 ( .A1(T7997_Y), .B0(T1009_Y), .B1(T10026_Y),     .A0(T10316_Y), .Y(T13022_Y));
KC_OAI22_X1 T13038 ( .A1(T10044_Y), .B0(T10317_Y), .B1(T1457_Y),     .A0(T7999_Y), .Y(T13038_Y));
KC_OAI22_X1 T13037 ( .A1(T10044_Y), .B0(T10026_Y), .B1(T15497_Y),     .A0(T7997_Y), .Y(T13037_Y));
KC_OAI22_X1 T13036 ( .A1(T10044_Y), .B0(T10043_Y), .B1(T16308_Y),     .A0(T7998_Y), .Y(T13036_Y));
KC_OAI22_X1 T13035 ( .A1(T10044_Y), .B0(T10047_Y), .B1(T16414_Y),     .A0(T7977_Y), .Y(T13035_Y));
KC_OAI22_X1 T13050 ( .A1(T16040_Y), .B0(T5879_Y), .B1(T10173_Y),     .A0(T15014_Y), .Y(T13050_Y));
KC_OAI22_X1 T13202 ( .A1(T7799_Y), .B0(T8025_Y), .B1(T1089_Y),     .A0(T16377_Y), .Y(T13202_Y));
KC_OAI22_X1 T13025 ( .A1(T10328_Y), .B0(T1060_Y), .B1(T8025_Y),     .A0(T16377_Y), .Y(T13025_Y));
KC_OAI22_X1 T13049 ( .A1(T12752_Y), .B0(T1362_Y), .B1(T10144_Y),     .A0(T4902_Y), .Y(T13049_Y));
KC_OAI22_X1 T13026 ( .A1(T15152_Y), .B0(T2620_Y), .B1(T15470_Y),     .A0(T16437_Y), .Y(T13026_Y));
KC_OAI22_X1 T13189 ( .A1(T6200_Y), .B0(T6520_Y), .B1(T2339_Y),     .A0(T11752_Y), .Y(T13189_Y));
KC_OAI22_X1 T13183 ( .A1(T6198_Y), .B0(T6519_Y), .B1(T2339_Y),     .A0(T11757_Y), .Y(T13183_Y));
KC_OAI22_X1 T12983 ( .A1(T291_Y), .B0(T6518_Y), .B1(T15332_Y),     .A0(T11044_Y), .Y(T12983_Y));
KC_OAI22_X1 T13196 ( .A1(T6543_Y), .B0(T6519_Y), .B1(T15332_Y),     .A0(T11047_Y), .Y(T13196_Y));
KC_OAI22_X1 T13195 ( .A1(T6498_Y), .B0(T6522_Y), .B1(T15332_Y),     .A0(T11045_Y), .Y(T13195_Y));
KC_OAI22_X1 T13030 ( .A1(T15478_Y), .B0(T1991_Y), .B1(T1124_Y),     .A0(T5881_Y), .Y(T13030_Y));
KC_OAI22_X1 T13040 ( .A1(T2604_Y), .B0(T2628_Q), .B1(T2034_Y),     .A0(T5363_Q), .Y(T13040_Y));
KC_OAI22_X1 T13303 ( .A1(T15906_Y), .B0(T6737_Y), .B1(T5444_Y),     .A0(T4931_Y), .Y(T13303_Y));
KC_OAI22_X1 T13114 ( .A1(T15943_Y), .B0(T2239_Y), .B1(T8238_Y),     .A0(T2751_Y), .Y(T13114_Y));
KC_OAI22_X1 T13107 ( .A1(T15943_Y), .B0(T6026_Y), .B1(T8238_Y),     .A0(T2127_Y), .Y(T13107_Y));
KC_OAI22_X1 T13101 ( .A1(T15943_Y), .B0(T5902_Y), .B1(T8238_Y),     .A0(T15854_Y), .Y(T13101_Y));
KC_OAI22_X1 T13100 ( .A1(T15916_Y), .B0(T5878_Y), .B1(T8238_Y),     .A0(T15855_Y), .Y(T13100_Y));
KC_OAI22_X1 T13099 ( .A1(T15943_Y), .B0(T5902_Y), .B1(T8238_Y),     .A0(T15853_Y), .Y(T13099_Y));
KC_OAI22_X1 T13098 ( .A1(T15943_Y), .B0(T5878_Y), .B1(T8238_Y),     .A0(T15856_Y), .Y(T13098_Y));
KC_OAI22_X1 T13117 ( .A1(T8238_Y), .B0(T2848_Y), .B1(T10739_Y),     .A0(T2237_Q), .Y(T13117_Y));
KC_OAI22_X1 T13144 ( .A1(T16489_Y), .B0(T2802_Y), .B1(T5991_Y),     .A0(T12808_Y), .Y(T13144_Y));
KC_OAI22_X1 T13267 ( .A1(T6184_Y), .B0(T15590_Y), .B1(T11665_Y),     .A0(T1788_Y), .Y(T13267_Y));
KC_OAI22_X1 T13156 ( .A1(T12228_Y), .B0(T6000_Y), .B1(T1786_Y),     .A0(T2854_Y), .Y(T13156_Y));
KC_OAI22_X1 T13149 ( .A1(T11032_Y), .B0(T2802_Y), .B1(T2239_Y),     .A0(T15712_Y), .Y(T13149_Y));
KC_OAI22_X1 T13148 ( .A1(T5002_Y), .B0(T2802_Y), .B1(T6004_Y),     .A0(T16130_Y), .Y(T13148_Y));
KC_OAI22_X1 T13322 ( .A1(T11032_Y), .B0(T6101_Y), .B1(T5002_Y),     .A0(T15633_Y), .Y(T13322_Y));
KC_OAI22_X1 T13310 ( .A1(T6184_Y), .B0(T5902_Y), .B1(T11665_Y),     .A0(T2246_Y), .Y(T13310_Y));
KC_OAI22_X1 T13163 ( .A1(T6184_Y), .B0(T5983_Y), .B1(T11665_Y),     .A0(T2250_Y), .Y(T13163_Y));
KC_OAI22_X1 T13159 ( .A1(T6184_Y), .B0(T6040_Y), .B1(T11665_Y),     .A0(T2280_Y), .Y(T13159_Y));
KC_OAI22_X1 T13158 ( .A1(T15618_Y), .B0(T6055_Y), .B1(T11665_Y),     .A0(T2280_Y), .Y(T13158_Y));
KC_OAI22_X1 T13157 ( .A1(T6184_Y), .B0(T6026_Y), .B1(T11665_Y),     .A0(T2245_Y), .Y(T13157_Y));
KC_OAI22_X1 T13178 ( .A1(T6180_Y), .B0(T2247_Y), .B1(T12064_Y),     .A0(T6225_Y), .Y(T13178_Y));
KC_OAI22_X1 T13194 ( .A1(T6541_Y), .B0(T6520_Y), .B1(T15332_Y),     .A0(T11825_Y), .Y(T13194_Y));
KC_OAI22_X1 T13003 ( .A1(T9667_Y), .B0(T6592_Y), .B1(T6456_Y),     .A0(T6760_Y), .Y(T13003_Y));
KC_OAI22_X1 T13001 ( .A1(T9652_Y), .B0(T6592_Y), .B1(T478_Y),     .A0(T6760_Y), .Y(T13001_Y));
KC_OAI22_X1 T13210 ( .A1(T9836_Y), .B0(T2620_Y), .B1(T1109_Y),     .A0(T875_Y), .Y(T13210_Y));
KC_OAI22_X1 T13209 ( .A1(T9938_Y), .B0(T2620_Y), .B1(T15473_Y),     .A0(T875_Y), .Y(T13209_Y));
KC_OAI22_X1 T13032 ( .A1(T1986_Y), .B0(T1994_Y), .B1(T9971_Y),     .A0(T2005_Q), .Y(T13032_Y));
KC_OAI22_X1 T13027 ( .A1(T10118_Y), .B0(T2620_Y), .B1(T1097_Y),     .A0(T875_Y), .Y(T13027_Y));
KC_OAI22_X1 T13047 ( .A1(T15090_Y), .B0(T2620_Y), .B1(T4852_Y),     .A0(T875_Y), .Y(T13047_Y));
KC_OAI22_X1 T13046 ( .A1(T15088_Y), .B0(T2620_Y), .B1(T1524_Y),     .A0(T875_Y), .Y(T13046_Y));
KC_OAI22_X1 T13039 ( .A1(T16368_Y), .B0(T2611_Y), .B1(T2615_Y),     .A0(T10059_Y), .Y(T13039_Y));
KC_OAI22_X1 T13073 ( .A1(T12790_Y), .B0(T5766_Y), .B1(T11009_Y),     .A0(T5783_Y), .Y(T13073_Y));
KC_OAI22_X1 T13106 ( .A1(T8238_Y), .B0(T15574_Y), .B1(T3401_Y),     .A0(T3355_Y), .Y(T13106_Y));
KC_OAI22_X1 T13123 ( .A1(T15974_Y), .B0(T6235_Y), .B1(T15943_Y),     .A0(T2839_Y), .Y(T13123_Y));
KC_OAI22_X1 T13143 ( .A1(T15974_Y), .B0(T2803_Y), .B1(T4991_Y),     .A0(T16039_Y), .Y(T13143_Y));
KC_OAI22_X1 T13164 ( .A1(T6087_Y), .B0(T16167_Y), .B1(T6039_Y),     .A0(T2618_Q), .Y(T13164_Y));
KC_OAI22_X1 T13175 ( .A1(T3429_Y), .B0(T5523_Y), .B1(T16105_Y),     .A0(T10622_Y), .Y(T13175_Y));
KC_OAI22_X1 T13193 ( .A1(T3489_Y), .B0(T6531_Y), .B1(T2937_Y),     .A0(T2929_Y), .Y(T13193_Y));
KC_OAI22_X1 T13000 ( .A1(T9663_Y), .B0(T6592_Y), .B1(T423_Y),     .A0(T6760_Y), .Y(T13000_Y));
KC_OAI22_X1 T12998 ( .A1(T8523_Y), .B0(T6592_Y), .B1(T15397_Y),     .A0(T6760_Y), .Y(T12998_Y));
KC_OAI22_X1 T13062 ( .A1(T5730_Y), .B0(T5730_Y), .B1(T16181_Y),     .A0(T5735_Y), .Y(T13062_Y));
KC_OAI22_X1 T13072 ( .A1(T3845_Y), .B0(T5773_Y), .B1(T5427_Y),     .A0(T15863_Y), .Y(T13072_Y));
KC_OAI22_X1 T12981 ( .A1(T5062_Y), .B0(T5062_Y), .B1(T5062_Y),     .A0(T3307_Y), .Y(T12981_Y));
KC_OAI22_X1 T13319 ( .A1(T5051_Y), .B0(T6081_Y), .B1(T10979_Y),     .A0(T6044_Y), .Y(T13319_Y));
KC_OAI22_X1 T13162 ( .A1(T6064_Y), .B0(T2824_Y), .B1(T11029_Y),     .A0(T15802_Q), .Y(T13162_Y));
KC_OAI22_X1 T13161 ( .A1(T15615_Y), .B0(T3468_Y), .B1(T12829_Y),     .A0(T6156_Y), .Y(T13161_Y));
KC_OAI22_X1 T13160 ( .A1(T6081_Y), .B0(T6069_Y), .B1(T10968_Y),     .A0(T3516_Y), .Y(T13160_Y));
KC_OAI22_X1 T13177 ( .A1(T3390_Y), .B0(T4070_Y), .B1(T4018_Y),     .A0(T4024_Y), .Y(T13177_Y));
KC_OAI22_X1 T13173 ( .A1(T3427_Y), .B0(T10619_Y), .B1(T6181_Y),     .A0(T12283_Y), .Y(T13173_Y));
KC_OAI22_X1 T13172 ( .A1(T6087_Y), .B0(T12271_Y), .B1(T12322_Y),     .A0(T12254_Y), .Y(T13172_Y));
KC_OAI22_X1 T13327 ( .A1(T16135_Y), .B0(T3514_Y), .B1(T2880_Y),     .A0(T5109_Y), .Y(T13327_Y));
KC_OAI22_X1 T13190 ( .A1(T10609_Y), .B0(T2865_Y), .B1(T12256_Y),     .A0(T16148_Y), .Y(T13190_Y));
KC_OAI22_X1 T13188 ( .A1(T4127_Y), .B0(T3489_Y), .B1(T5520_Y),     .A0(T3528_Q), .Y(T13188_Y));
KC_OAI22_X1 T13187 ( .A1(T3427_Y), .B0(T3489_Y), .B1(T2893_Y),     .A0(T6236_Y), .Y(T13187_Y));
KC_OAI22_X1 T13186 ( .A1(T3481_Y), .B0(T10985_Y), .B1(T6209_Y),     .A0(T12108_Y), .Y(T13186_Y));
KC_OAI22_X1 T13182 ( .A1(T5046_Y), .B0(T12304_Y), .B1(T6188_Y),     .A0(T12299_Y), .Y(T13182_Y));
KC_OAI22_X1 T13308 ( .A1(T3840_Y), .B0(T5101_Y), .B1(T3841_Y),     .A0(T12342_Y), .Y(T13308_Y));
KC_OAI22_X1 T13078 ( .A1(T3794_Y), .B0(T5767_Y), .B1(T5800_Y),     .A0(T11410_Y), .Y(T13078_Y));
KC_OAI22_X1 T13077 ( .A1(T5770_Y), .B0(T3795_Y), .B1(T15867_Y),     .A0(T5101_Y), .Y(T13077_Y));
KC_OAI22_X1 T13066 ( .A1(T5816_Y), .B0(T5806_Y), .B1(T15867_Y),     .A0(T5101_Y), .Y(T13066_Y));
KC_OAI22_X1 T13093 ( .A1(T3834_Y), .B0(T8188_Y), .B1(T3842_Y),     .A0(T11409_Y), .Y(T13093_Y));
KC_OAI22_X1 T13092 ( .A1(T11405_Y), .B0(T15908_Y), .B1(T3829_Y),     .A0(T8190_Y), .Y(T13092_Y));
KC_OAI22_X1 T13087 ( .A1(T3840_Y), .B0(T5101_Y), .B1(T5800_Y),     .A0(T144_Q), .Y(T13087_Y));
KC_OAI22_X1 T13086 ( .A1(T3849_Y), .B0(T15873_Y), .B1(T5803_Y),     .A0(T4450_Y), .Y(T13086_Y));
KC_OAI22_X1 T13081 ( .A1(T3828_Y), .B0(T16154_Y), .B1(T15897_Y),     .A0(T14550_Q), .Y(T13081_Y));
KC_OAI22_X1 T13124 ( .A1(T4510_Y), .B0(T5120_Y), .B1(T11511_Y),     .A0(T11507_Y), .Y(T13124_Y));
KC_OAI22_X1 T13176 ( .A1(T6176_Y), .B0(T6155_Y), .B1(T11708_Y),     .A0(T2806_Y), .Y(T13176_Y));
KC_OAI22_X1 T13174 ( .A1(T6532_Y), .B0(T6157_Y), .B1(T6155_Y),     .A0(T2838_Y), .Y(T13174_Y));
KC_OAI22_X1 T13171 ( .A1(T6137_Y), .B0(T4095_Y), .B1(T12289_Y),     .A0(T10602_Y), .Y(T13171_Y));
KC_OAI22_X1 T13169 ( .A1(T4077_Y), .B0(T16124_Y), .B1(T8382_Y),     .A0(T8380_Y), .Y(T13169_Y));
KC_OAI22_X1 T13168 ( .A1(T3443_Y), .B0(T6517_Y), .B1(T4085_Y),     .A0(T6157_Y), .Y(T13168_Y));
KC_OAI22_X1 T13166 ( .A1(T3368_Y), .B0(T6527_Y), .B1(T4085_Y),     .A0(T10567_Y), .Y(T13166_Y));
KC_OAI22_X1 T13180 ( .A1(T6188_Y), .B0(T6079_Y), .B1(T5051_Y),     .A0(T6824_Y), .Y(T13180_Y));
KC_OAI22_X1 T13179 ( .A1(T3427_Y), .B0(T2865_Y), .B1(T12304_Y),     .A0(T6824_Y), .Y(T13179_Y));
KC_OAI22_X1 T13305 ( .A1(T4389_Y), .B0(T3826_Y), .B1(T4448_Y),     .A0(T16154_Y), .Y(T13305_Y));
KC_OAI22_X1 T13076 ( .A1(T3842_Y), .B0(T11313_Y), .B1(T4486_Y),     .A0(T14942_Q), .Y(T13076_Y));
KC_OAI22_X1 T13071 ( .A1(T5800_Y), .B0(T5767_Y), .B1(T5778_Y),     .A0(T16153_Y), .Y(T13071_Y));
KC_OAI22_X1 T13090 ( .A1(T4394_Y), .B0(T14551_Q), .B1(T5802_Y),     .A0(T14546_Q), .Y(T13090_Y));
KC_OAI22_X1 T13085 ( .A1(T4426_Y), .B0(T4462_Y), .B1(T4459_Y),     .A0(T4459_Y), .Y(T13085_Y));
KC_OAI22_X1 T13084 ( .A1(T4383_Y), .B0(T15869_Y), .B1(T3833_Y),     .A0(T4486_Y), .Y(T13084_Y));
KC_OAI22_X1 T13083 ( .A1(T4446_Y), .B0(T3833_Y), .B1(T4382_Y),     .A0(T3824_Y), .Y(T13083_Y));
KC_OAI22_X1 T13118 ( .A1(T12355_Y), .B0(T4532_Y), .B1(T15994_Y),     .A0(T16466_Q), .Y(T13118_Y));
KC_OAI22_X1 T13115 ( .A1(T6780_Y), .B0(T4474_Y), .B1(T15969_Y),     .A0(T11574_Y), .Y(T13115_Y));
KC_OAI22_X1 T13309 ( .A1(T11995_Y), .B0(T4623_Y), .B1(T12345_Y),     .A0(T16112_Y), .Y(T13309_Y));
KC_OAI22_X1 T13184 ( .A1(T6202_Y), .B0(T6103_Y), .B1(T4739_Y),     .A0(T12302_Y), .Y(T13184_Y));
KC_OAI22_X1 T13185 ( .A1(T4736_Y), .B0(T15630_Y), .B1(T12308_Y),     .A0(T6103_Y), .Y(T13185_Y));
KC_OAI22_X1 T13280 ( .A1(T636_Y), .B0(T7867_Y), .B1(T7866_Y),     .A0(T9363_Y), .Y(T13280_Y));
KC_OAI22_X1 T13279 ( .A1(T718_Y), .B0(T763_Y), .B1(T7869_Y),     .A0(T16379_Y), .Y(T13279_Y));
KC_OAI22_X1 T13278 ( .A1(T15433_Y), .B0(T763_Y), .B1(T7866_Y),     .A0(T12883_Y), .Y(T13278_Y));
KC_OAI22_X1 T13277 ( .A1(T854_Y), .B0(T15654_Y), .B1(T7869_Y),     .A0(T7800_Y), .Y(T13277_Y));
KC_OAI22_X1 T13275 ( .A1(T6629_Y), .B0(T6819_Y), .B1(T10918_Y),     .A0(T7591_Y), .Y(T13275_Y));
KC_OAI22_X1 T13273 ( .A1(T6699_Y), .B0(T6835_Y), .B1(T10918_Y),     .A0(T7414_Y), .Y(T13273_Y));
KC_OAI22_X1 T13203 ( .A1(T10331_Y), .B0(T8025_Y), .B1(T15471_Y),     .A0(T16377_Y), .Y(T13203_Y));
KC_OAI22_X1 T13314 ( .A1(T8238_Y), .B0(T2848_Y), .B1(T10659_Y),     .A0(T2236_Q), .Y(T13314_Y));
KC_OAI22_X1 T13311 ( .A1(T6184_Y), .B0(T2239_Y), .B1(T11665_Y),     .A0(T16042_Y), .Y(T13311_Y));
KC_OAI22_X1 T13289 ( .A1(T2037_Y), .B0(T16366_Y), .B1(T2036_Y),     .A0(T15502_Y), .Y(T13289_Y));
KC_OAI22_X1 T13320 ( .A1(T6181_Y), .B0(T16167_Y), .B1(T6155_Y),     .A0(T12104_Y), .Y(T13320_Y));
KC_OAI22_X1 T13321 ( .A1(T6176_Y), .B0(T2865_Y), .B1(T8508_Y),     .A0(T15802_Q), .Y(T13321_Y));
KC_OAI22_X1 T13318 ( .A1(T5054_Y), .B0(T6392_Y), .B1(T5522_Y),     .A0(T15233_Y), .Y(T13318_Y));
KC_OAI22_X1 T13205 ( .A1(T9666_Y), .B0(T6592_Y), .B1(T15383_Y),     .A0(T6760_Y), .Y(T13205_Y));
KC_OAI22_X1 T13326 ( .A1(T4091_Y), .B0(T6587_Y), .B1(T10580_Y),     .A0(T10564_Y), .Y(T13326_Y));
KC_OAI22_X1 T13325 ( .A1(T10580_Y), .B0(T6176_Y), .B1(T4085_Y),     .A0(T6155_Y), .Y(T13325_Y));
KC_OAI22_X1 T13307 ( .A1(T15867_Y), .B0(T5101_Y), .B1(T3794_Y),     .A0(T5800_Y), .Y(T13307_Y));
KC_OAI22_X1 T13306 ( .A1(T5842_Y), .B0(T8452_Y), .B1(T3856_Y),     .A0(T16153_Y), .Y(T13306_Y));
KC_OAI22_X1 T13296 ( .A1(T11967_Y), .B0(T3825_Y), .B1(T3857_Y),     .A0(T5789_Y), .Y(T13296_Y));
KC_OAI22_X1 T15875 ( .A1(T15869_Y), .B0(T3836_Y), .B1(T15557_Y),     .A0(T5815_Y), .Y(T15875_Y));
KC_OAI22_X1 T13304 ( .A1(T4448_Y), .B0(T3794_Y), .B1(T4382_Y),     .A0(T11348_Y), .Y(T13304_Y));
KC_OAI22_X1 T13295 ( .A1(T11966_Y), .B0(T16153_Y), .B1(T4445_Y),     .A0(T14548_Q), .Y(T13295_Y));
KC_OAI22_X1 T13002 ( .A1(T9638_Y), .B0(T6592_Y), .B1(T431_Y),     .A0(T6760_Y), .Y(T13002_Y));
KC_OAI22_X1 T12999 ( .A1(T8525_Y), .B0(T6592_Y), .B1(T424_Y),     .A0(T6760_Y), .Y(T12999_Y));
KC_OAI22_X1 T13091 ( .A1(T5783_Y), .B0(T5824_Y), .B1(T5840_Y),     .A0(T144_Q), .Y(T13091_Y));
KC_OAI22_X1 T13089 ( .A1(T5827_Y), .B0(T4445_Y), .B1(T4440_Y),     .A0(T144_Q), .Y(T13089_Y));
KC_OAI22_X1 T13109 ( .A1(T3401_Y), .B0(T5908_Y), .B1(T2168_Y),     .A0(T5896_Y), .Y(T13109_Y));
KC_OAI22_X1 T13122 ( .A1(T15943_Y), .B0(T10932_Y), .B1(T2168_Y),     .A0(T6081_Y), .Y(T13122_Y));
KC_OAI22_X1 T13116 ( .A1(T5925_Y), .B0(T5878_Y), .B1(T8238_Y),     .A0(T8241_Y), .Y(T13116_Y));
KC_OAI22_X1 T13134 ( .A1(T15592_Y), .B0(T11571_Y), .B1(T5956_Y),     .A0(T11451_Y), .Y(T13134_Y));
KC_OAI22_X1 T13191 ( .A1(T2888_Y), .B0(T12038_Y), .B1(T6583_Y),     .A0(T6560_Y), .Y(T13191_Y));
KC_OAI22_X1 T13313 ( .A1(T8235_Y), .B0(T5119_Y), .B1(T3945_Y),     .A0(T11570_Y), .Y(T13313_Y));
KC_DFFSNHQ_X1 T13216 ( .Q(T13216_Q), .D(T102_Y), .CK(T138_Y),     .SN(T7073_Y));
KC_DFFSNHQ_X1 T13229 ( .Q(T13229_Q), .D(T8628_Y), .CK(T138_Y),     .SN(T7074_Y));
KC_DFFSNHQ_X1 T13241 ( .Q(T13241_Q), .D(T16314_Y), .CK(T4828_Y),     .SN(T14976_Y));
KC_DFFSNHQ_X1 T13263 ( .Q(T13263_Q), .D(T4850_Y), .CK(T4851_Y),     .SN(T993_Y));
KC_DFFSNHQ_X1 T13033 ( .Q(T13033_Q), .D(T16159_Y), .CK(T1140_Y),     .SN(T10697_Y));
KC_DFFSNHQ_X1 T13059 ( .Q(T13059_Q), .D(T5381_Y), .CK(T1604_Y),     .SN(T13053_SN));
KC_DFFSNHQ_X1 T13058 ( .Q(T13058_Q), .D(T10206_Y), .CK(T10226_Y),     .SN(T13053_SN));
KC_DFFSNHQ_X1 T13053 ( .Q(T13053_Q), .D(T1302_Y), .CK(T1604_Y),     .SN(T13053_SN));
KC_DFFSNHQ_X1 T16231 ( .Q(T16231_Q), .D(T1678_Q), .CK(T16407_Y),     .SN(T2000_Y));
KC_DFFSNHQ_X1 T13019 ( .Q(T13019_Q), .D(T5313_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13010 ( .Q(T13010_Q), .D(T13018_Q), .CK(T16407_Y),     .SN(T2000_Y));
KC_DFFSNHQ_X1 T13008 ( .Q(T13008_Q), .D(T16231_Q), .CK(T16407_Y),     .SN(T2000_Y));
KC_DFFSNHQ_X1 T13031 ( .Q(T13031_Q), .D(T15071_Y), .CK(T15190_Y),     .SN(T14999_Y));
KC_DFFSNHQ_X1 T13020 ( .Q(T13020_Q), .D(T1970_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13017 ( .Q(T13017_Q), .D(T13014_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13016 ( .Q(T13016_Q), .D(T13013_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13015 ( .Q(T13015_Q), .D(T13016_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13014 ( .Q(T13014_Q), .D(T1978_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13013 ( .Q(T13013_Q), .D(T13017_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13007 ( .Q(T13007_Q), .D(T1981_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13006 ( .Q(T13006_Q), .D(T13020_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13042 ( .Q(T13042_Q), .D(T13048_Q), .CK(T5725_Y),     .SN(T15003_Y));
KC_DFFSNHQ_X1 T13293 ( .Q(T13293_Q), .D(T13052_Q), .CK(T2050_Y),     .SN(T2062_Y));
KC_DFFSNHQ_X1 T13051 ( .Q(T13051_Q), .D(T13293_Q), .CK(T2050_Y),     .SN(T2062_Y));
KC_DFFSNHQ_X1 T13065 ( .Q(T13065_Q), .D(T2120_Y), .CK(T14554_Q),     .SN(T15034_Y));
KC_DFFSNHQ_X1 T13108 ( .Q(T13108_Q), .D(T13107_Y), .CK(T14960_Q),     .SN(T15015_Y));
KC_DFFSNHQ_X1 T13132 ( .Q(T13132_Q), .D(T2170_Y), .CK(T14570_Q),     .SN(T15015_Y));
KC_DFFSNHQ_X1 T13129 ( .Q(T13129_Q), .D(T12813_Y), .CK(T14564_Q),     .SN(T15015_Y));
KC_DFFSNHQ_X1 T13127 ( .Q(T13127_Q), .D(T12809_Y), .CK(T14564_Q),     .SN(T15015_Y));
KC_DFFSNHQ_X1 T13298 ( .Q(T13298_Q), .D(T5017_Y), .CK(T3264_Y),     .SN(T15034_Y));
KC_DFFSNHQ_X1 T13112 ( .Q(T13112_Q), .D(T2743_Y), .CK(T14557_Q),     .SN(T15013_Y));
KC_DFFSNHQ_X1 T13111 ( .Q(T13111_Q), .D(T2745_Y), .CK(T14557_Q),     .SN(T15013_Y));
KC_DFFSNHQ_X1 T13128 ( .Q(T13128_Q), .D(T13116_Y), .CK(T14557_Q),     .SN(T15015_Y));
KC_DFFSNHQ_X1 T13141 ( .Q(T13141_Q), .D(T11593_Y), .CK(T2790_Y),     .SN(T14566_Q));
KC_DFFSNHQ_X1 T13140 ( .Q(T13140_Q), .D(T13141_Q), .CK(T2790_Y),     .SN(T14566_Q));
KC_DFFSNHQ_X1 T13133 ( .Q(T13133_Q), .D(T5998_Y), .CK(T14564_Q),     .SN(T2169_Y));
KC_DFFSNHQ_X1 T13079 ( .Q(T13079_Q), .D(T3212_Y), .CK(T14542_Q),     .SN(T3221_Y));
KC_DFFSNHQ_X1 T13067 ( .Q(T13067_Q), .D(T3208_Y), .CK(T3209_Y),     .SN(T3221_Y));
KC_DFFSNHQ_X1 T13297 ( .Q(T13297_Q), .D(T5450_Y), .CK(T3264_Y),     .SN(T15034_Y));
KC_DFFSNHQ_X1 T13110 ( .Q(T13110_Q), .D(T3261_Y), .CK(T3264_Y),     .SN(T15034_Y));
KC_DFFSNHQ_X1 T13096 ( .Q(T13096_Q), .D(T3275_Y), .CK(T3264_Y),     .SN(T2709_Y));
KC_DFFSNHQ_X1 T13126 ( .Q(T13126_Q), .D(T11515_Y), .CK(T2790_Y),     .SN(T2761_Y));
KC_DFFSNHQ_X1 T13130 ( .Q(T13130_Q), .D(T4473_Y), .CK(T3879_Y),     .SN(T3888_Y));
KC_DFFSNHQ_X1 T13312 ( .Q(T13312_Q), .D(T5472_Y), .CK(T3993_Y),     .SN(T5023_Y));
KC_DFFSNHQ_X1 T13155 ( .Q(T13155_Q), .D(T3987_Y), .CK(T3993_Y),     .SN(T15035_Y));
KC_DFFSNHQ_X1 T13154 ( .Q(T13154_Q), .D(T3985_Y), .CK(T3993_Y),     .SN(T15035_Y));
KC_DFFSNHQ_X1 T13151 ( .Q(T13151_Q), .D(T3983_Y), .CK(T3993_Y),     .SN(T15035_Y));
KC_DFFSNHQ_X1 T13150 ( .Q(T13150_Q), .D(T3986_Y), .CK(T3993_Y),     .SN(T15035_Y));
KC_DFFSNHQ_X1 T13145 ( .Q(T13145_Q), .D(T12236_Y), .CK(T4045_Y),     .SN(T15035_Y));
KC_DFFSNHQ_X1 T13167 ( .Q(T13167_Q), .D(T9100_Y), .CK(T2736_Y),     .SN(T15022_Y));
KC_DFFSNHQ_X1 T13165 ( .Q(T13165_Q), .D(T6421_Y), .CK(T2736_Y),     .SN(T15022_Y));
KC_DFFSNHQ_X1 T13323 ( .Q(T13323_Q), .D(T15758_Y), .CK(T4728_Y),     .SN(T15022_Y));
KC_DFFSNHQ_X1 T13198 ( .Q(T13198_Q), .D(T13058_Q), .CK(T10226_Y),     .SN(T13053_SN));
KC_DFFSNHQ_X1 T13292 ( .Q(T13292_Q), .D(T12111_Y), .CK(T2078_Y),     .SN(T2063_Y));
KC_DFFSNHQ_X1 T13324 ( .Q(T13324_Q), .D(T15759_Y), .CK(T4728_Y),     .SN(T15022_Y));
KC_DFFSNHQ_X1 T13018 ( .Q(T13018_Q), .D(T1682_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13012 ( .Q(T13012_Q), .D(T1982_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13009 ( .Q(T13009_Q), .D(T13019_Q), .CK(T16407_Y),     .SN(T14988_Y));
KC_DFFSNHQ_X1 T13029 ( .Q(T13029_Q), .D(T1680_Y), .CK(T15190_Y),     .SN(T2000_Y));
KC_DFFSNHQ_X1 T13028 ( .Q(T13028_Q), .D(T2026_Y), .CK(T2667_Y),     .SN(T2582_Y));
KC_DFFSNHQ_X1 T13048 ( .Q(T13048_Q), .D(T2045_Y), .CK(T5725_Y),     .SN(T15003_Y));
KC_DFFSNHQ_X1 T13291 ( .Q(T13291_Q), .D(T13051_Q), .CK(T2050_Y),     .SN(T2062_Y));
KC_DFFSNHQ_X1 T13052 ( .Q(T13052_Q), .D(T13063_Q), .CK(T2050_Y),     .SN(T2062_Y));
KC_DFFSNHQ_X1 T13063 ( .Q(T13063_Q), .D(T12148_Y), .CK(T2050_Y),     .SN(T2062_Y));
KC_DFFSNHQ_X1 T13056 ( .Q(T13056_Q), .D(T1291_Y), .CK(T1604_Y),     .SN(T13053_SN));
KC_DFFSNHQ_X1 T13070 ( .Q(T13070_Q), .D(T15700_Y), .CK(T3879_Y),     .SN(T2688_Y));
KC_DFFSNHQ_X1 T13316 ( .Q(T13316_Q), .D(T3301_Y), .CK(T3264_Y),     .SN(T15034_Y));
KC_DFFSNHQ_X1 T13104 ( .Q(T13104_Q), .D(T3271_Y), .CK(T3264_Y),     .SN(T15034_Y));
KC_DFFSNHQ_X1 T13103 ( .Q(T13103_Q), .D(T3302_Y), .CK(T3264_Y),     .SN(T15034_Y));
KC_DFFSNHQ_X1 T13119 ( .Q(T13119_Q), .D(T3313_Y), .CK(T3264_Y),     .SN(T5023_Y));
KC_DFFSNHQ_X1 T13136 ( .Q(T13136_Q), .D(T12827_Y), .CK(T14564_Q),     .SN(T2169_Y));
KC_DFFSNHQ_X1 T13135 ( .Q(T13135_Q), .D(T14566_Q), .CK(T2790_Y),     .SN(T1748_Y));
KC_DFFSNHQ_X1 T12980 ( .Q(T12980_Q), .D(T5468_Y), .CK(T3993_Y),     .SN(T5023_Y));
KC_DFFSNHQ_X1 T13170 ( .Q(T13170_Q), .D(T2869_Y), .CK(T14557_Q),     .SN(T15021_Y));
KC_DFFSNHQ_X1 T13299 ( .Q(T13299_Q), .D(T2720_Y), .CK(T3264_Y),     .SN(T15034_Y));
KC_OAI13_X1 T12472 ( .B0(T8560_Y), .A(T8561_Y), .B2(T5202_Q),     .Y(T12472_Y), .B1(T106_Q));
KC_OAI13_X1 T12471 ( .B0(T5614_Y), .A(T15318_Y), .B2(T1201_Y),     .Y(T12471_Y), .B1(T16310_Y));
KC_OAI13_X1 T12470 ( .B0(T5612_Y), .A(T878_Y), .B2(T5598_Y),     .Y(T12470_Y), .B1(T8540_Y));
KC_OAI13_X1 T12475 ( .B0(T6912_Y), .A(T878_Y), .B2(T6913_Y),     .Y(T12475_Y), .B1(T6935_Y));
KC_OAI13_X1 T12614 ( .B0(T7677_Y), .A(T646_Y), .B2(T7698_Y),     .Y(T12614_Y), .B1(T7584_Y));
KC_OAI13_X1 T12608 ( .B0(T9396_Y), .A(T878_Y), .B2(T16317_Y),     .Y(T12608_Y), .B1(T7584_Y));
KC_OAI13_X1 T12527 ( .B0(T15025_Y), .A(T13260_Y), .B2(T4810_Q),     .Y(T12527_Y), .B1(T180_Q));
KC_OAI13_X1 T12606 ( .B0(T7570_Y), .A(T7579_Y), .B2(T9384_Y),     .Y(T12606_Y), .B1(T7832_Y));
KC_OAI13_X1 T12722 ( .B0(T7857_Y), .A(T8102_Y), .B2(T8949_Y),     .Y(T12722_Y), .B1(T8081_Y));
KC_OAI13_X1 T12477 ( .B0(T8852_Y), .A(T8573_Y), .B2(T6931_Y),     .Y(T12477_Y), .B1(T311_Y));
KC_OAI13_X1 T12496 ( .B0(T8894_Y), .A(T8624_Y), .B2(T7069_Y),     .Y(T12496_Y), .B1(T6348_Y));
KC_OAI13_X1 T12890 ( .B0(T8895_Y), .A(T9514_Y), .B2(T9515_Y),     .Y(T12890_Y), .B1(T6613_Y));
KC_OAI13_X1 T12882 ( .B0(T9411_Y), .A(T9348_Y), .B2(T9346_Y),     .Y(T12882_Y), .B1(T6671_Y));
KC_OAI13_X1 T12576 ( .B0(T8664_Y), .A(T8803_Y), .B2(T189_Q),     .Y(T12576_Y), .B1(T183_Q));
KC_OAI13_X1 T12615 ( .B0(T916_Y), .A(T8750_Y), .B2(T5350_Q),     .Y(T12615_Y), .B1(T5357_Q));
KC_OAI13_X1 T12611 ( .B0(T9001_Y), .A(T8712_Y), .B2(T7605_Y),     .Y(T12611_Y), .B1(T6662_Y));
KC_OAI13_X1 T12605 ( .B0(T528_Q), .A(T8894_Y), .B2(T550_Q),     .Y(T12605_Y), .B1(T544_Q));
KC_OAI13_X1 T12885 ( .B0(T8036_Y), .A(T960_Y), .B2(T8903_Y),     .Y(T12885_Y), .B1(T8072_Y));
KC_OAI13_X1 T12889 ( .B0(T9160_Y), .A(T4811_Y), .B2(T9472_Q),     .Y(T12889_Y), .B1(T16183_Y));
KC_OAI13_X1 T12478 ( .B0(T245_Y), .A(T6954_Y), .B2(T8593_Y),     .Y(T12478_Y), .B1(T820_Q));
KC_OAI13_X1 T12476 ( .B0(T301_Y), .A(T6916_Y), .B2(T8570_Y),     .Y(T12476_Y), .B1(T823_Q));
KC_OAI13_X1 T12474 ( .B0(T244_Y), .A(T6901_Y), .B2(T8565_Y),     .Y(T12474_Y), .B1(T815_Q));
KC_OAI13_X1 T12880 ( .B0(T315_Y), .A(T6299_Y), .B2(T9264_Y),     .Y(T12880_Y), .B1(T848_Q));
KC_OAI13_X1 T12495 ( .B0(T334_Y), .A(T6329_Y), .B2(T8617_Y),     .Y(T12495_Y), .B1(T838_Q));
KC_OAI13_X1 T12494 ( .B0(T9409_Y), .A(T8621_Y), .B2(T9277_Y),     .Y(T12494_Y), .B1(T333_Y));
KC_OAI13_X1 T12492 ( .B0(T8802_Y), .A(T8620_Y), .B2(T6922_Y),     .Y(T12492_Y), .B1(T339_Y));
KC_OAI13_X1 T12491 ( .B0(T9408_Y), .A(T8622_Y), .B2(T9281_Y),     .Y(T12491_Y), .B1(T6332_Y));
KC_OAI13_X1 T12575 ( .B0(T14981_Y), .A(T9412_Y), .B2(T690_Q),     .Y(T12575_Y), .B1(T688_Q));
KC_OAI13_X1 T12609 ( .B0(T8854_Y), .A(T8721_Y), .B2(T7598_Y),     .Y(T12609_Y), .B1(T737_Y));
KC_OAI13_X1 T12604 ( .B0(T932_Y), .A(T8693_Y), .B2(T729_Q),     .Y(T12604_Y), .B1(T724_Q));
KC_OAI13_X1 T12720 ( .B0(T8061_Y), .A(T1196_Y), .B2(T8943_Y),     .Y(T12720_Y), .B1(T13250_Y));
KC_OAI13_X1 T12749 ( .B0(T9094_Y), .A(T1004_Q), .B2(T770_Q),     .Y(T12749_Y), .B1(T780_Q));
KC_OAI13_X1 T12497 ( .B0(T317_Y), .A(T7080_Y), .B2(T8612_Y),     .Y(T12497_Y), .B1(T834_Q));
KC_OAI13_X1 T12525 ( .B0(T9410_Y), .A(T8641_Y), .B2(T7300_Y),     .Y(T12525_Y), .B1(T15647_Y));
KC_OAI13_X1 T12610 ( .B0(T886_Y), .A(T7591_Y), .B2(T7610_Y),     .Y(T12610_Y), .B1(T7616_Y));
KC_OAI13_X1 T12884 ( .B0(T9401_Y), .A(T1196_Y), .B2(T989_Y),     .Y(T12884_Y), .B1(T7880_Y));
KC_OAI13_X1 T12883 ( .B0(T763_Y), .A(T8792_Y), .B2(T16159_Y),     .Y(T12883_Y), .B1(T4872_Y));
KC_OAI13_X1 T12678 ( .B0(T15654_Y), .A(T8792_Y), .B2(T16159_Y),     .Y(T12678_Y), .B1(T4872_Y));
KC_OAI13_X1 T12677 ( .B0(T7868_Y), .A(T8792_Y), .B2(T16159_Y),     .Y(T12677_Y), .B1(T4872_Y));
KC_OAI13_X1 T12612 ( .B0(T7613_Y), .A(T12613_Y), .B2(T7633_Y),     .Y(T12612_Y), .B1(T7634_Y));
KC_OAI13_X1 T12603 ( .B0(T7556_Y), .A(T7951_Y), .B2(T1084_Q),     .Y(T12603_Y), .B1(T5343_Q));
KC_OAI13_X1 T12690 ( .B0(T1208_Q), .A(T9916_Y), .B2(T9918_Y),     .Y(T12690_Y), .B1(T9919_Y));
KC_OAI13_X1 T12724 ( .B0(T4848_Y), .A(T16383_Y), .B2(T16275_Y),     .Y(T12724_Y), .B1(T13033_Q));
KC_OAI13_X1 T12752 ( .B0(T13125_Y), .A(T10144_Y), .B2(T1362_Y),     .Y(T12752_Y), .B1(T10934_Y));
KC_OAI13_X1 T12771 ( .B0(T1168_Y), .A(T12208_Y), .B2(T5412_Y),     .Y(T12771_Y), .B1(T5411_Y));
KC_OAI13_X1 T12513 ( .B0(T6481_Y), .A(T7139_Y), .B2(T372_Y),     .Y(T12513_Y), .B1(T13575_Q));
KC_OAI13_X1 T12509 ( .B0(T6481_Y), .A(T7192_Y), .B2(T367_Y),     .Y(T12509_Y), .B1(T13586_Q));
KC_OAI13_X1 T12498 ( .B0(T6481_Y), .A(T7141_Y), .B2(T355_Y),     .Y(T12498_Y), .B1(T13597_Q));
KC_OAI13_X1 T12582 ( .B0(T15393_Y), .A(T1453_Y), .B2(T1476_Y),     .Y(T12582_Y), .B1(T7489_Y));
KC_OAI13_X1 T12577 ( .B0(T15393_Y), .A(T1453_Y), .B2(T1476_Y),     .Y(T12577_Y), .B1(T7541_Y));
KC_OAI13_X1 T12977 ( .B0(T15393_Y), .A(T1493_Y), .B2(T1476_Y),     .Y(T12977_Y), .B1(T10015_Y));
KC_OAI13_X1 T12726 ( .B0(T10015_Y), .A(T1493_Y), .B2(T7703_Y),     .Y(T12726_Y), .B1(T1476_Y));
KC_OAI13_X1 T12908 ( .B0(T15393_Y), .A(T1418_Y), .B2(T4884_Y),     .Y(T12908_Y), .B1(T6993_Y));
KC_OAI13_X1 T12490 ( .B0(T15393_Y), .A(T1418_Y), .B2(T4884_Y),     .Y(T12490_Y), .B1(T9542_Y));
KC_OAI13_X1 T12489 ( .B0(T15393_Y), .A(T1418_Y), .B2(T4884_Y),     .Y(T12489_Y), .B1(T6983_Y));
KC_OAI13_X1 T12488 ( .B0(T15670_Y), .A(T1419_Y), .B2(T4884_Y),     .Y(T12488_Y), .B1(T6992_Y));
KC_OAI13_X1 T12486 ( .B0(T15670_Y), .A(T1419_Y), .B2(T4884_Y),     .Y(T12486_Y), .B1(T10389_Y));
KC_OAI13_X1 T12485 ( .B0(T15393_Y), .A(T1418_Y), .B2(T4884_Y),     .Y(T12485_Y), .B1(T9543_Y));
KC_OAI13_X1 T12483 ( .B0(T6993_Y), .A(T1418_Y), .B2(T16448_Y),     .Y(T12483_Y), .B1(T4884_Y));
KC_OAI13_X1 T12482 ( .B0(T9542_Y), .A(T1418_Y), .B2(T16448_Y),     .Y(T12482_Y), .B1(T4884_Y));
KC_OAI13_X1 T12481 ( .B0(T6983_Y), .A(T1418_Y), .B2(T16448_Y),     .Y(T12481_Y), .B1(T4884_Y));
KC_OAI13_X1 T12480 ( .B0(T9543_Y), .A(T1418_Y), .B2(T16448_Y),     .Y(T12480_Y), .B1(T4884_Y));
KC_OAI13_X1 T12479 ( .B0(T6992_Y), .A(T1419_Y), .B2(T16448_Y),     .Y(T12479_Y), .B1(T4884_Y));
KC_OAI13_X1 T12512 ( .B0(T6481_Y), .A(T7215_Y), .B2(T15379_Y),     .Y(T12512_Y), .B1(T13609_Q));
KC_OAI13_X1 T12511 ( .B0(T6481_Y), .A(T7127_Y), .B2(T369_Y),     .Y(T12511_Y), .B1(T14728_Q));
KC_OAI13_X1 T12510 ( .B0(T6481_Y), .A(T7131_Y), .B2(T370_Y),     .Y(T12510_Y), .B1(T13573_Q));
KC_OAI13_X1 T12508 ( .B0(T6481_Y), .A(T7190_Y), .B2(T351_Y),     .Y(T12508_Y), .B1(T13607_Q));
KC_OAI13_X1 T12507 ( .B0(T6481_Y), .A(T7132_Y), .B2(T15375_Y),     .Y(T12507_Y), .B1(T13584_Q));
KC_OAI13_X1 T12506 ( .B0(T6481_Y), .A(T7130_Y), .B2(T354_Y),     .Y(T12506_Y), .B1(T13606_Q));
KC_OAI13_X1 T12505 ( .B0(T6481_Y), .A(T7187_Y), .B2(T353_Y),     .Y(T12505_Y), .B1(T13603_Q));
KC_OAI13_X1 T12504 ( .B0(T6481_Y), .A(T7189_Y), .B2(T366_Y),     .Y(T12504_Y), .B1(T13585_Q));
KC_OAI13_X1 T12501 ( .B0(T6481_Y), .A(T7179_Y), .B2(T358_Y),     .Y(T12501_Y), .B1(T14726_Q));
KC_OAI13_X1 T12500 ( .B0(T6481_Y), .A(T7178_Y), .B2(T364_Y),     .Y(T12500_Y), .B1(T14727_Q));
KC_OAI13_X1 T12499 ( .B0(T6481_Y), .A(T7140_Y), .B2(T365_Y),     .Y(T12499_Y), .B1(T14725_Q));
KC_OAI13_X1 T12921 ( .B0(T1483_Y), .A(T5668_Y), .B2(T15676_Y),     .Y(T12921_Y), .B1(T13691_Q));
KC_OAI13_X1 T12920 ( .B0(T9721_Y), .A(T1453_Y), .B2(T7703_Y),     .Y(T12920_Y), .B1(T1476_Y));
KC_OAI13_X1 T12919 ( .B0(T1483_Y), .A(T5667_Y), .B2(T6749_Y),     .Y(T12919_Y), .B1(T14662_Q));
KC_OAI13_X1 T12542 ( .B0(T1483_Y), .A(T7336_Y), .B2(T402_Y),     .Y(T12542_Y), .B1(T13717_Q));
KC_OAI13_X1 T12541 ( .B0(T1483_Y), .A(T5666_Y), .B2(T15395_Y),     .Y(T12541_Y), .B1(T13716_Q));
KC_OAI13_X1 T12536 ( .B0(T1483_Y), .A(T7335_Y), .B2(T401_Y),     .Y(T12536_Y), .B1(T13692_Q));
KC_OAI13_X1 T12906 ( .B0(T7952_Y), .A(T10809_Y), .B2(T15667_Y),     .Y(T12906_Y), .B1(T14661_Q));
KC_OAI13_X1 T12586 ( .B0(T15393_Y), .A(T1453_Y), .B2(T1476_Y),     .Y(T12586_Y), .B1(T9720_Y));
KC_OAI13_X1 T12585 ( .B0(T7541_Y), .A(T1453_Y), .B2(T7703_Y),     .Y(T12585_Y), .B1(T1476_Y));
KC_OAI13_X1 T12584 ( .B0(T9720_Y), .A(T1453_Y), .B2(T7703_Y),     .Y(T12584_Y), .B1(T1476_Y));
KC_OAI13_X1 T12581 ( .B0(T7489_Y), .A(T1453_Y), .B2(T7703_Y),     .Y(T12581_Y), .B1(T1476_Y));
KC_OAI13_X1 T12580 ( .B0(T1483_Y), .A(T7508_Y), .B2(T587_Y),     .Y(T12580_Y), .B1(T13812_Q));
KC_OAI13_X1 T12579 ( .B0(T15393_Y), .A(T1453_Y), .B2(T1476_Y),     .Y(T12579_Y), .B1(T9721_Y));
KC_OAI13_X1 T12578 ( .B0(T1483_Y), .A(T7488_Y), .B2(T589_Y),     .Y(T12578_Y), .B1(T13978_Q));
KC_OAI13_X1 T12638 ( .B0(T1483_Y), .A(T7790_Y), .B2(T15439_Y),     .Y(T12638_Y), .B1(T13960_Q));
KC_OAI13_X1 T12637 ( .B0(T1483_Y), .A(T7699_Y), .B2(T15436_Y),     .Y(T12637_Y), .B1(T13942_Q));
KC_OAI13_X1 T12636 ( .B0(T1483_Y), .A(T7784_Y), .B2(T853_Y),     .Y(T12636_Y), .B1(T13943_Q));
KC_OAI13_X1 T12635 ( .B0(T9810_Y), .A(T1492_Y), .B2(T7703_Y),     .Y(T12635_Y), .B1(T7707_Y));
KC_OAI13_X1 T12634 ( .B0(T1483_Y), .A(T7785_Y), .B2(T851_Y),     .Y(T12634_Y), .B1(T14013_Q));
KC_OAI13_X1 T12623 ( .B0(T1483_Y), .A(T7783_Y), .B2(T821_Y),     .Y(T12623_Y), .B1(T13958_Q));
KC_OAI13_X1 T12622 ( .B0(T1483_Y), .A(T7706_Y), .B2(T827_Y),     .Y(T12622_Y), .B1(T13959_Q));
KC_OAI13_X1 T12621 ( .B0(T15393_Y), .A(T1492_Y), .B2(T7707_Y),     .Y(T12621_Y), .B1(T9810_Y));
KC_OAI13_X1 T12896 ( .B0(T15470_Y), .A(T10762_Y), .B2(T1483_Y),     .Y(T12896_Y), .B1(T14613_Q));
KC_OAI13_X1 T12893 ( .B0(T7952_Y), .A(T16441_Y), .B2(T1080_Y),     .Y(T12893_Y), .B1(T14612_Q));
KC_OAI13_X1 T12702 ( .B0(T1483_Y), .A(T7967_Y), .B2(T1081_Y),     .Y(T12702_Y), .B1(T14614_Q));
KC_OAI13_X1 T12701 ( .B0(T1483_Y), .A(T7958_Y), .B2(T1033_Y),     .Y(T12701_Y), .B1(T14128_Q));
KC_OAI13_X1 T12700 ( .B0(T1483_Y), .A(T7957_Y), .B2(T1027_Y),     .Y(T12700_Y), .B1(T14127_Q));
KC_OAI13_X1 T12699 ( .B0(T1483_Y), .A(T8014_Y), .B2(T1083_Y),     .Y(T12699_Y), .B1(T14616_Q));
KC_OAI13_X1 T12698 ( .B0(T1483_Y), .A(T8015_Y), .B2(T1082_Y),     .Y(T12698_Y), .B1(T14615_Q));
KC_OAI13_X1 T12695 ( .B0(T7952_Y), .A(T8012_Y), .B2(T1038_Y),     .Y(T12695_Y), .B1(T14129_Q));
KC_OAI13_X1 T12694 ( .B0(T7952_Y), .A(T7959_Y), .B2(T1035_Y),     .Y(T12694_Y), .B1(T14126_Q));
KC_OAI13_X1 T12693 ( .B0(T7952_Y), .A(T8005_Y), .B2(T15468_Y),     .Y(T12693_Y), .B1(T14608_Q));
KC_OAI13_X1 T12978 ( .B0(T15393_Y), .A(T1493_Y), .B2(T1476_Y),     .Y(T12978_Y), .B1(T10018_Y));
KC_OAI13_X1 T12730 ( .B0(T10017_Y), .A(T1493_Y), .B2(T7703_Y),     .Y(T12730_Y), .B1(T1476_Y));
KC_OAI13_X1 T12729 ( .B0(T15393_Y), .A(T1493_Y), .B2(T1476_Y),     .Y(T12729_Y), .B1(T10014_Y));
KC_OAI13_X1 T12728 ( .B0(T10014_Y), .A(T1493_Y), .B2(T7703_Y),     .Y(T12728_Y), .B1(T1476_Y));
KC_OAI13_X1 T12727 ( .B0(T15393_Y), .A(T1493_Y), .B2(T1476_Y),     .Y(T12727_Y), .B1(T10017_Y));
KC_OAI13_X1 T12484 ( .B0(T15670_Y), .A(T1419_Y), .B2(T4884_Y),     .Y(T12484_Y), .B1(T9540_Y));
KC_OAI13_X1 T12544 ( .B0(T6481_Y), .A(T7348_Y), .B2(T15396_Y),     .Y(T12544_Y), .B1(T14720_Q));
KC_OAI13_X1 T12633 ( .B0(T15393_Y), .A(T1492_Y), .B2(T7707_Y),     .Y(T12633_Y), .B1(T9787_Y));
KC_OAI13_X1 T12632 ( .B0(T15393_Y), .A(T1492_Y), .B2(T7707_Y),     .Y(T12632_Y), .B1(T7781_Y));
KC_OAI13_X1 T12631 ( .B0(T7704_Y), .A(T1492_Y), .B2(T7703_Y),     .Y(T12631_Y), .B1(T7707_Y));
KC_OAI13_X1 T12630 ( .B0(T15393_Y), .A(T1492_Y), .B2(T7707_Y),     .Y(T12630_Y), .B1(T7704_Y));
KC_OAI13_X1 T12628 ( .B0(T7781_Y), .A(T1492_Y), .B2(T7703_Y),     .Y(T12628_Y), .B1(T7707_Y));
KC_OAI13_X1 T12616 ( .B0(T9787_Y), .A(T1492_Y), .B2(T7703_Y),     .Y(T12616_Y), .B1(T7707_Y));
KC_OAI13_X1 T12697 ( .B0(T7952_Y), .A(T8006_Y), .B2(T16398_Y),     .Y(T12697_Y), .B1(T14609_Q));
KC_OAI13_X1 T12696 ( .B0(T7952_Y), .A(T8007_Y), .B2(T1026_Y),     .Y(T12696_Y), .B1(T14124_Q));
KC_OAI13_X1 T12692 ( .B0(T7952_Y), .A(T8008_Y), .B2(T16396_Y),     .Y(T12692_Y), .B1(T14125_Q));
KC_OAI13_X1 T12750 ( .B0(T1366_Y), .A(T1365_Y), .B2(T15529_Y),     .Y(T12750_Y), .B1(T1362_Y));
KC_OAI13_X1 T12828 ( .B0(T15973_Y), .A(T11595_Y), .B2(T10225_Y),     .Y(T12828_Y), .B1(T15974_Y));
KC_OAI13_X1 T12941 ( .B0(T635_Y), .A(T15154_Y), .B2(T4973_Y),     .Y(T12941_Y), .B1(T635_Y));
KC_OAI13_X1 T12719 ( .B0(T9973_Y), .A(T9971_Y), .B2(T16369_Y),     .Y(T12719_Y), .B1(T868_Y));
KC_OAI13_X1 T12713 ( .B0(T1990_Y), .A(T11257_Y), .B2(T2016_Q),     .Y(T12713_Y), .B1(T1106_Y));
KC_OAI13_X1 T12709 ( .B0(T9951_Y), .A(T11258_Y), .B2(T2028_Q),     .Y(T12709_Y), .B1(T868_Y));
KC_OAI13_X1 T12738 ( .B0(T1509_Y), .A(T5395_Y), .B2(T16305_Y),     .Y(T12738_Y), .B1(T12096_Y));
KC_OAI13_X1 T12737 ( .B0(T2053_Q), .A(T2043_Y), .B2(T1495_Y),     .Y(T12737_Y), .B1(T2042_Y));
KC_OAI13_X1 T12736 ( .B0(T2957_Y), .A(T15506_Y), .B2(T1527_Y),     .Y(T12736_Y), .B1(T9974_Y));
KC_OAI13_X1 T12734 ( .B0(T10065_Y), .A(T2057_Y), .B2(T16365_Y),     .Y(T12734_Y), .B1(T15503_Y));
KC_OAI13_X1 T12770 ( .B0(T10183_Y), .A(T10185_Y), .B2(T10183_Y),     .Y(T12770_Y), .B1(T10183_Y));
KC_OAI13_X1 T12812 ( .B0(T15943_Y), .A(T12198_Y), .B2(T16302_Y),     .Y(T12812_Y), .B1(T8250_Y));
KC_OAI13_X1 T12824 ( .B0(T6026_Y), .A(T2201_Y), .B2(T16096_Y),     .Y(T12824_Y), .B1(T2217_Y));
KC_OAI13_X1 T12823 ( .B0(T5982_Y), .A(T11585_Y), .B2(T16070_Y),     .Y(T12823_Y), .B1(T2217_Y));
KC_OAI13_X1 T12822 ( .B0(T5902_Y), .A(T6301_Y), .B2(T16074_Y),     .Y(T12822_Y), .B1(T2217_Y));
KC_OAI13_X1 T12821 ( .B0(T5878_Y), .A(T2198_Y), .B2(T16072_Y),     .Y(T12821_Y), .B1(T2217_Y));
KC_OAI13_X1 T12820 ( .B0(T15590_Y), .A(T2203_Y), .B2(T16075_Y),     .Y(T12820_Y), .B1(T2217_Y));
KC_OAI13_X1 T12819 ( .B0(T5983_Y), .A(T2210_Y), .B2(T16097_Y),     .Y(T12819_Y), .B1(T2217_Y));
KC_OAI13_X1 T12818 ( .B0(T6004_Y), .A(T2202_Y), .B2(T16071_Y),     .Y(T12818_Y), .B1(T2217_Y));
KC_OAI13_X1 T12835 ( .B0(T4957_Y), .A(T15164_Y), .B2(T6342_Y),     .Y(T12835_Y), .B1(T6013_Y));
KC_OAI13_X1 T12869 ( .B0(T2358_Y), .A(T2352_Y), .B2(T15638_Y),     .Y(T12869_Y), .B1(T2317_Y));
KC_OAI13_X1 T12879 ( .B0(T4978_Y), .A(T4980_Y), .B2(T4963_Y),     .Y(T12879_Y), .B1(T2369_Y));
KC_OAI13_X1 T12521 ( .B0(T6481_Y), .A(T2428_Y), .B2(T15384_Y),     .Y(T12521_Y), .B1(T14765_Q));
KC_OAI13_X1 T12520 ( .B0(T6481_Y), .A(T2429_Y), .B2(T375_Y),     .Y(T12520_Y), .B1(T13656_Q));
KC_OAI13_X1 T12548 ( .B0(T6456_Y), .A(T4990_Y), .B2(T6481_Y),     .Y(T12548_Y), .B1(T13782_Q));
KC_OAI13_X1 T12933 ( .B0(T632_Y), .A(T11932_Y), .B2(T14836_Q),     .Y(T12933_Y), .B1(T2447_Y));
KC_OAI13_X1 T12601 ( .B0(T7952_Y), .A(T3056_Y), .B2(T15424_Y),     .Y(T12601_Y), .B1(T14856_Q));
KC_OAI13_X1 T12591 ( .B0(T7952_Y), .A(T2479_Y), .B2(T6762_Y),     .Y(T12591_Y), .B1(T13835_Q));
KC_OAI13_X1 T12587 ( .B0(T7952_Y), .A(T5272_Y), .B2(T609_Y),     .Y(T12587_Y), .B1(T14857_Q));
KC_OAI13_X1 T12670 ( .B0(T7952_Y), .A(T5850_Y), .B2(T871_Y),     .Y(T12670_Y), .B1(T14859_Q));
KC_OAI13_X1 T12942 ( .B0(T16245_Y), .A(T2554_Y), .B2(T1482_Y),     .Y(T12942_Y), .B1(T14892_Q));
KC_OAI13_X1 T12715 ( .B0(T15473_Y), .A(T2563_Y), .B2(T16245_Y),     .Y(T12715_Y), .B1(T14882_Q));
KC_OAI13_X1 T12714 ( .B0(T1109_Y), .A(T5329_Y), .B2(T16245_Y),     .Y(T12714_Y), .B1(T14881_Q));
KC_OAI13_X1 T12708 ( .B0(T1097_Y), .A(T2569_Y), .B2(T7952_Y),     .Y(T12708_Y), .B1(T14152_Q));
KC_OAI13_X1 T12747 ( .B0(T4852_Y), .A(T16256_Y), .B2(T16245_Y),     .Y(T12747_Y), .B1(T14366_Q));
KC_OAI13_X1 T12744 ( .B0(T1524_Y), .A(T2595_Y), .B2(T16245_Y),     .Y(T12744_Y), .B1(T14345_Q));
KC_OAI13_X1 T12740 ( .B0(T1509_Y), .A(T2607_Y), .B2(T10058_Y),     .Y(T12740_Y), .B1(T1527_Y));
KC_OAI13_X1 T12735 ( .B0(T5920_Y), .A(T2057_Y), .B2(T15501_Y),     .Y(T12735_Y), .B1(T15503_Y));
KC_OAI13_X1 T12768 ( .B0(T16245_Y), .A(T2634_Y), .B2(T4871_Y),     .Y(T12768_Y), .B1(T14425_Q));
KC_OAI13_X1 T12763 ( .B0(T16245_Y), .A(T2636_Y), .B2(T4864_Y),     .Y(T12763_Y), .B1(T14403_Q));
KC_OAI13_X1 T12762 ( .B0(T16245_Y), .A(T2638_Y), .B2(T4867_Y),     .Y(T12762_Y), .B1(T14363_Q));
KC_OAI13_X1 T12758 ( .B0(T16245_Y), .A(T2635_Y), .B2(T4886_Y),     .Y(T12758_Y), .B1(T14427_Q));
KC_OAI13_X1 T12757 ( .B0(T16245_Y), .A(T2637_Y), .B2(T4883_Y),     .Y(T12757_Y), .B1(T14426_Q));
KC_OAI13_X1 T12967 ( .B0(T12847_Y), .A(T12049_Y), .B2(T2822_Y),     .Y(T12967_Y), .B1(T2818_Y));
KC_OAI13_X1 T12848 ( .B0(T11686_Y), .A(T6561_Y), .B2(T10595_Y),     .Y(T12848_Y), .B1(T6115_Y));
KC_OAI13_X1 T12847 ( .B0(T6576_Y), .A(T10611_Y), .B2(T8261_Y),     .Y(T12847_Y), .B1(T16132_Y));
KC_OAI13_X1 T12974 ( .B0(T2921_Y), .A(T11742_Y), .B2(T6513_Y),     .Y(T12974_Y), .B1(T6239_Y));
KC_OAI13_X1 T12872 ( .B0(T2883_Y), .A(T6561_Y), .B2(T11723_Y),     .Y(T12872_Y), .B1(T12873_Y));
KC_OAI13_X1 T12867 ( .B0(T2896_Y), .A(T12106_Y), .B2(T12101_Y),     .Y(T12867_Y), .B1(T12103_Y));
KC_OAI13_X1 T12862 ( .B0(T2914_Y), .A(T6196_Y), .B2(T2899_Y),     .Y(T12862_Y), .B1(T2900_Y));
KC_OAI13_X1 T12861 ( .B0(T2904_Y), .A(T6196_Y), .B2(T6513_Y),     .Y(T12861_Y), .B1(T2902_Y));
KC_OAI13_X1 T12468 ( .B0(T11740_Y), .A(T6196_Y), .B2(T2357_Y),     .Y(T12468_Y), .B1(T2914_Y));
KC_OAI13_X1 T12877 ( .B0(T2938_Y), .A(T10999_Y), .B2(T4055_Y),     .Y(T12877_Y), .B1(T11000_Y));
KC_OAI13_X1 T12876 ( .B0(T2961_Y), .A(T12297_Y), .B2(T2959_Y),     .Y(T12876_Y), .B1(T5540_Y));
KC_OAI13_X1 T12923 ( .B0(T2447_Y), .A(T2999_Y), .B2(T15679_Y),     .Y(T12923_Y), .B1(T13639_Q));
KC_OAI13_X1 T12519 ( .B0(T15383_Y), .A(T2996_Y), .B2(T2447_Y),     .Y(T12519_Y), .B1(T14761_Q));
KC_OAI13_X1 T12518 ( .B0(T2447_Y), .A(T2997_Y), .B2(T374_Y),     .Y(T12518_Y), .B1(T13653_Q));
KC_OAI13_X1 T12945 ( .B0(T424_Y), .A(T3016_Y), .B2(T2447_Y),     .Y(T12945_Y), .B1(T14930_Q));
KC_OAI13_X1 T12547 ( .B0(T15397_Y), .A(T3019_Y), .B2(T2447_Y),     .Y(T12547_Y), .B1(T13755_Q));
KC_OAI13_X1 T12668 ( .B0(T3076_Y), .A(T3678_Y), .B2(T3073_Y),     .Y(T12668_Y), .B1(T3679_Y));
KC_OAI13_X1 T12667 ( .B0(T3068_Y), .A(T3678_Y), .B2(T3073_Y),     .Y(T12667_Y), .B1(T3679_Y));
KC_OAI13_X1 T12666 ( .B0(T3076_Y), .A(T3678_Y), .B2(T3679_Y),     .Y(T12666_Y), .B1(T15441_Y));
KC_OAI13_X1 T12657 ( .B0(T7952_Y), .A(T2510_Y), .B2(T874_Y),     .Y(T12657_Y), .B1(T14083_Q));
KC_OAI13_X1 T12650 ( .B0(T7952_Y), .A(T5550_Y), .B2(T870_Y),     .Y(T12650_Y), .B1(T14069_Q));
KC_OAI13_X1 T12646 ( .B0(T15441_Y), .A(T3678_Y), .B2(T3679_Y),     .Y(T12646_Y), .B1(T3068_Y));
KC_OAI13_X1 T12645 ( .B0(T3068_Y), .A(T3678_Y), .B2(T880_Y),     .Y(T12645_Y), .B1(T15441_Y));
KC_OAI13_X1 T12644 ( .B0(T880_Y), .A(T3678_Y), .B2(T15441_Y),     .Y(T12644_Y), .B1(T3076_Y));
KC_OAI13_X1 T12717 ( .B0(T16245_Y), .A(T5326_Y), .B2(T1138_Y),     .Y(T12717_Y), .B1(T14198_Q));
KC_OAI13_X1 T12716 ( .B0(T16245_Y), .A(T5863_Y), .B2(T1136_Y),     .Y(T12716_Y), .B1(T14172_Q));
KC_OAI13_X1 T12951 ( .B0(T15826_Y), .A(T5765_Y), .B2(T15819_Y),     .Y(T12951_Y), .B1(T8188_Y));
KC_OAI13_X1 T12790 ( .B0(T3203_Y), .A(T16160_Y), .B2(T11983_Y),     .Y(T12790_Y), .B1(T11336_Y));
KC_OAI13_X1 T12789 ( .B0(T11354_Y), .A(T16160_Y), .B2(T12132_Y),     .Y(T12789_Y), .B1(T3799_Y));
KC_OAI13_X1 T12960 ( .B0(T16000_Y), .A(T15162_Y), .B2(T3332_Y),     .Y(T12960_Y), .B1(T16000_Y));
KC_OAI13_X1 T12826 ( .B0(T15981_Y), .A(T3322_Y), .B2(T15579_Y),     .Y(T12826_Y), .B1(T5483_Y));
KC_OAI13_X1 T12817 ( .B0(T3316_Y), .A(T6278_Y), .B2(T15591_Y),     .Y(T12817_Y), .B1(T3363_Y));
KC_OAI13_X1 T12829 ( .B0(T12357_Y), .A(T5996_Y), .B2(T15005_Y),     .Y(T12829_Y), .B1(T15882_Y));
KC_OAI13_X1 T12852 ( .B0(T3459_Y), .A(T6141_Y), .B2(T2839_Y),     .Y(T12852_Y), .B1(T10588_Y));
KC_OAI13_X1 T12846 ( .B0(T3443_Y), .A(T12972_Y), .B2(T4089_Y),     .Y(T12846_Y), .B1(T6119_Y));
KC_OAI13_X1 T12845 ( .B0(T3445_Y), .A(T15622_Y), .B2(T3458_Y),     .Y(T12845_Y), .B1(T6080_Y));
KC_OAI13_X1 T12464 ( .B0(T4073_Y), .A(T5045_Y), .B2(T6119_Y),     .Y(T12464_Y), .B1(T3515_Y));
KC_OAI13_X1 T12866 ( .B0(T13182_Y), .A(T6561_Y), .B2(T6820_Y),     .Y(T12866_Y), .B1(T3485_Y));
KC_OAI13_X1 T12865 ( .B0(T3487_Y), .A(T6561_Y), .B2(T3497_Y),     .Y(T12865_Y), .B1(T2925_Y));
KC_OAI13_X1 T12875 ( .B0(T6510_Y), .A(T6561_Y), .B2(T3521_Q),     .Y(T12875_Y), .B1(T10570_Y));
KC_OAI13_X1 T12955 ( .B0(T3787_Y), .A(T11394_Y), .B2(T11977_Y),     .Y(T12955_Y), .B1(T15868_Y));
KC_OAI13_X1 T12792 ( .B0(T3794_Y), .A(T3796_Y), .B2(T413_Y),     .Y(T12792_Y), .B1(T5780_Y));
KC_OAI13_X1 T12788 ( .B0(T5801_Y), .A(T4465_Q), .B2(T5771_Y),     .Y(T12788_Y), .B1(T11365_Y));
KC_OAI13_X1 T12797 ( .B0(T11380_Y), .A(T11393_Y), .B2(T5830_Y),     .Y(T12797_Y), .B1(T11375_Y));
KC_OAI13_X1 T12807 ( .B0(T5874_Y), .A(T3872_Y), .B2(T5870_Y),     .Y(T12807_Y), .B1(T15571_Y));
KC_OAI13_X1 T12806 ( .B0(T4491_Q), .A(T3900_Q), .B2(T3885_Q),     .Y(T12806_Y), .B1(T4493_Q));
KC_OAI13_X1 T12804 ( .B0(T15919_Y), .A(T3866_Y), .B2(T15917_Y),     .Y(T12804_Y), .B1(T15918_Y));
KC_OAI13_X1 T12814 ( .B0(T3914_Y), .A(T5100_Y), .B2(T15578_Y),     .Y(T12814_Y), .B1(T5120_Y));
KC_OAI13_X1 T12965 ( .B0(T4058_Y), .A(T4068_Y), .B2(T11636_Y),     .Y(T12965_Y), .B1(T6078_Y));
KC_OAI13_X1 T12842 ( .B0(T8167_Y), .A(T4025_Y), .B2(T6084_Y),     .Y(T12842_Y), .B1(T3417_Y));
KC_OAI13_X1 T12841 ( .B0(T8167_Y), .A(T4025_Y), .B2(T6084_Y),     .Y(T12841_Y), .B1(T3417_Y));
KC_OAI13_X1 T12857 ( .B0(T4064_Y), .A(T8503_Y), .B2(T11714_Y),     .Y(T12857_Y), .B1(T6437_Y));
KC_OAI13_X1 T12856 ( .B0(T12253_Y), .A(T16140_Y), .B2(T5522_Y),     .Y(T12856_Y), .B1(T4017_Y));
KC_OAI13_X1 T12851 ( .B0(T3445_Y), .A(T11711_Y), .B2(T11710_Y),     .Y(T12851_Y), .B1(T3443_Y));
KC_OAI13_X1 T12968 ( .B0(T16141_Y), .A(T10993_Y), .B2(T6111_Y),     .Y(T12968_Y), .B1(T6155_Y));
KC_OAI13_X1 T12975 ( .B0(T4204_Y), .A(T3025_Y), .B2(T3073_Y),     .Y(T12975_Y), .B1(T16449_Y));
KC_OAI13_X1 T12524 ( .B0(T15441_Y), .A(T3025_Y), .B2(T16449_Y),     .Y(T12524_Y), .B1(T10433_Y));
KC_OAI13_X1 T12523 ( .B0(T15441_Y), .A(T3585_Y), .B2(T16449_Y),     .Y(T12523_Y), .B1(T10432_Y));
KC_OAI13_X1 T12522 ( .B0(T15441_Y), .A(T3585_Y), .B2(T16449_Y),     .Y(T12522_Y), .B1(T4203_Y));
KC_OAI13_X1 T12517 ( .B0(T10433_Y), .A(T3025_Y), .B2(T3073_Y),     .Y(T12517_Y), .B1(T16449_Y));
KC_OAI13_X1 T12516 ( .B0(T15441_Y), .A(T3585_Y), .B2(T16449_Y),     .Y(T12516_Y), .B1(T4204_Y));
KC_OAI13_X1 T12515 ( .B0(T4203_Y), .A(T3025_Y), .B2(T3073_Y),     .Y(T12515_Y), .B1(T16449_Y));
KC_OAI13_X1 T12514 ( .B0(T10432_Y), .A(T3025_Y), .B2(T3073_Y),     .Y(T12514_Y), .B1(T16449_Y));
KC_OAI13_X1 T12664 ( .B0(T4267_Y), .A(T4283_Y), .B2(T3073_Y),     .Y(T12664_Y), .B1(T3679_Y));
KC_OAI13_X1 T12663 ( .B0(T15441_Y), .A(T4283_Y), .B2(T3679_Y),     .Y(T12663_Y), .B1(T4267_Y));
KC_OAI13_X1 T12661 ( .B0(T15441_Y), .A(T4283_Y), .B2(T3679_Y),     .Y(T12661_Y), .B1(T9860_Y));
KC_OAI13_X1 T12660 ( .B0(T9859_Y), .A(T4283_Y), .B2(T3073_Y),     .Y(T12660_Y), .B1(T3679_Y));
KC_OAI13_X1 T12656 ( .B0(T15441_Y), .A(T4283_Y), .B2(T3679_Y),     .Y(T12656_Y), .B1(T4266_Y));
KC_OAI13_X1 T12655 ( .B0(T4266_Y), .A(T4283_Y), .B2(T3073_Y),     .Y(T12655_Y), .B1(T3679_Y));
KC_OAI13_X1 T12643 ( .B0(T9860_Y), .A(T4283_Y), .B2(T3073_Y),     .Y(T12643_Y), .B1(T3679_Y));
KC_OAI13_X1 T12746 ( .B0(T4318_Y), .A(T3735_Y), .B2(T3073_Y),     .Y(T12746_Y), .B1(T7707_Y));
KC_OAI13_X1 T12745 ( .B0(T15441_Y), .A(T3735_Y), .B2(T7707_Y),     .Y(T12745_Y), .B1(T4318_Y));
KC_OAI13_X1 T12742 ( .B0(T10095_Y), .A(T3735_Y), .B2(T3073_Y),     .Y(T12742_Y), .B1(T7707_Y));
KC_OAI13_X1 T12741 ( .B0(T15441_Y), .A(T3735_Y), .B2(T7707_Y),     .Y(T12741_Y), .B1(T10095_Y));
KC_OAI13_X1 T12756 ( .B0(T16248_Y), .A(T3735_Y), .B2(T3073_Y),     .Y(T12756_Y), .B1(T7707_Y));
KC_OAI13_X1 T12755 ( .B0(T10096_Y), .A(T3735_Y), .B2(T3073_Y),     .Y(T12755_Y), .B1(T7707_Y));
KC_OAI13_X1 T12754 ( .B0(T15441_Y), .A(T3735_Y), .B2(T7707_Y),     .Y(T12754_Y), .B1(T16248_Y));
KC_OAI13_X1 T12753 ( .B0(T15441_Y), .A(T3735_Y), .B2(T7707_Y),     .Y(T12753_Y), .B1(T10096_Y));
KC_OAI13_X1 T12953 ( .B0(T8184_Y), .A(T144_Q), .B2(T4487_Q),     .Y(T12953_Y), .B1(T5767_Y));
KC_OAI13_X1 T12950 ( .B0(T4402_Y), .A(T15555_Y), .B2(T3792_Y),     .Y(T12950_Y), .B1(T16157_Y));
KC_OAI13_X1 T12791 ( .B0(T13076_Y), .A(T15838_Y), .B2(T16154_Y),     .Y(T12791_Y), .B1(T11322_Y));
KC_OAI13_X1 T12801 ( .B0(T4464_Y), .A(T4440_Y), .B2(T4487_Q),     .Y(T12801_Y), .B1(T4431_Y));
KC_OAI13_X1 T12796 ( .B0(T5760_Y), .A(T4445_Y), .B2(T145_Q),     .Y(T12796_Y), .B1(T5838_Y));
KC_OAI13_X1 T12795 ( .B0(T12796_Y), .A(T11393_Y), .B2(T15845_Y),     .Y(T12795_Y), .B1(T11421_Y));
KC_OAI13_X1 T12805 ( .B0(T15967_Y), .A(T15933_Y), .B2(T11451_Y),     .Y(T12805_Y), .B1(T5867_Y));
KC_OAI13_X1 T12803 ( .B0(T4505_Y), .A(T3896_Y), .B2(T5448_Y),     .Y(T12803_Y), .B1(T4505_Y));
KC_OAI13_X1 T12811 ( .B0(T10931_Y), .A(T4513_Y), .B2(T5459_Y),     .Y(T12811_Y), .B1(T12196_Y));
KC_OAI13_X1 T12810 ( .B0(T11521_Y), .A(T5156_Y), .B2(T11521_Y),     .Y(T12810_Y), .B1(T11521_Y));
KC_OAI13_X1 T12959 ( .B0(T4544_Y), .A(T5125_Y), .B2(T4562_Y),     .Y(T12959_Y), .B1(T5157_Y));
KC_OAI13_X1 T12825 ( .B0(T4548_Y), .A(T12233_Y), .B2(T11536_Y),     .Y(T12825_Y), .B1(T5986_Y));
KC_OAI13_X1 T12834 ( .B0(T8331_Y), .A(T6012_Y), .B2(T8331_Y),     .Y(T12834_Y), .B1(T5067_Y));
KC_OAI13_X1 T12833 ( .B0(T4580_Y), .A(T4595_Y), .B2(T5159_Q),     .Y(T12833_Y), .B1(T6022_Y));
KC_OAI13_X1 T12840 ( .B0(T4652_Y), .A(T4684_Y), .B2(T6030_Y),     .Y(T12840_Y), .B1(T8344_Y));
KC_OAI13_X1 T12839 ( .B0(T4657_Y), .A(T4678_Y), .B2(T8344_Y),     .Y(T12839_Y), .B1(T6042_Y));
KC_OAI13_X1 T12838 ( .B0(T6360_Y), .A(T2521_Y), .B2(T4689_Y),     .Y(T12838_Y), .B1(T15135_Y));
KC_OAI13_X1 T12837 ( .B0(T4646_Y), .A(T4681_Y), .B2(T6030_Y),     .Y(T12837_Y), .B1(T8457_Y));
KC_OAI13_X1 T12836 ( .B0(T16047_Y), .A(T4676_Y), .B2(T8457_Y),     .Y(T12836_Y), .B1(T6042_Y));
KC_OAI13_X1 T12855 ( .B0(T10981_Y), .A(T6448_Y), .B2(T16146_Y),     .Y(T12855_Y), .B1(T6169_Y));
KC_OAI13_X1 T12868 ( .B0(T4704_Y), .A(T6589_Y), .B2(T4758_Q),     .Y(T12868_Y), .B1(T4759_Q));
KC_OAI13_X1 T12881 ( .B0(T110_Y), .A(T6860_Y), .B2(T9292_Y),     .Y(T12881_Y), .B1(T826_Q));
KC_OAI13_X1 T12891 ( .B0(T10142_Y), .A(T972_Y), .B2(T1394_Y),     .Y(T12891_Y), .B1(T9987_Y));
KC_OAI13_X1 T12887 ( .B0(T10142_Y), .A(T972_Y), .B2(T10303_Y),     .Y(T12887_Y), .B1(T1394_Y));
KC_OAI13_X1 T12895 ( .B0(T7952_Y), .A(T10761_Y), .B2(T16399_Y),     .Y(T12895_Y), .B1(T14610_Q));
KC_OAI13_X1 T12892 ( .B0(T7952_Y), .A(T10759_Y), .B2(T15435_Y),     .Y(T12892_Y), .B1(T14607_Q));
KC_OAI13_X1 T12973 ( .B0(T2920_Y), .A(T10555_Y), .B2(T10551_Y),     .Y(T12973_Y), .B1(T2897_Y));
KC_OAI13_X1 T12970 ( .B0(T12971_Y), .A(T6561_Y), .B2(T13172_Y),     .Y(T12970_Y), .B1(T3484_Y));
KC_OAI13_X1 T12969 ( .B0(T2884_Y), .A(T6561_Y), .B2(T8376_Y),     .Y(T12969_Y), .B1(T12056_Y));
KC_OAI13_X1 T12963 ( .B0(T3307_Y), .A(T12981_Y), .B2(T3297_Y),     .Y(T12963_Y), .B1(T3299_Y));
KC_OAI13_X1 T12966 ( .B0(T4019_Y), .A(T16140_Y), .B2(T15709_Y),     .Y(T12966_Y), .B1(T4020_Y));
KC_OAI13_X1 T12957 ( .B0(T16029_Y), .A(T12239_Y), .B2(T11724_Y),     .Y(T12957_Y), .B1(T15610_Y));
KC_OAI13_X1 T12954 ( .B0(T6740_Y), .A(T10902_Y), .B2(T4457_Y),     .Y(T12954_Y), .B1(T5767_Y));
KC_OAI13_X1 T12907 ( .B0(T9540_Y), .A(T1419_Y), .B2(T16448_Y),     .Y(T12907_Y), .B1(T4884_Y));
KC_OAI13_X1 T12487 ( .B0(T9541_Y), .A(T1419_Y), .B2(T16448_Y),     .Y(T12487_Y), .B1(T4884_Y));
KC_OAI13_X1 T12909 ( .B0(T6481_Y), .A(T7188_Y), .B2(T15671_Y),     .Y(T12909_Y), .B1(T13657_Q));
KC_OAI13_X1 T12493 ( .B0(T8893_Y), .A(T8619_Y), .B2(T7052_Y),     .Y(T12493_Y), .B1(T334_Y));
KC_OAI13_X1 T12936 ( .B0(T7952_Y), .A(T3030_Y), .B2(T15902_Y),     .Y(T12936_Y), .B1(T14051_Q));
KC_OAI13_X1 T12574 ( .B0(T5252_Q), .A(T9324_Y), .B2(T9322_Y),     .Y(T12574_Y), .B1(T905_Y));
KC_OAI13_X1 T12675 ( .B0(T16245_Y), .A(T2499_Y), .B2(T884_Y),     .Y(T12675_Y), .B1(T14151_Q));
KC_OAI13_X1 T12671 ( .B0(T7952_Y), .A(T2506_Y), .B2(T866_Y),     .Y(T12671_Y), .B1(T14081_Q));
KC_OAI13_X1 T12669 ( .B0(T3068_Y), .A(T3678_Y), .B2(T3073_Y),     .Y(T12669_Y), .B1(T880_Y));
KC_OAI13_X1 T12665 ( .B0(T3076_Y), .A(T3678_Y), .B2(T3073_Y),     .Y(T12665_Y), .B1(T880_Y));
KC_OAI13_X1 T12662 ( .B0(T15441_Y), .A(T4283_Y), .B2(T3679_Y),     .Y(T12662_Y), .B1(T9859_Y));
KC_OAI13_X1 T12618 ( .B0(T1483_Y), .A(T7792_Y), .B2(T852_Y),     .Y(T12618_Y), .B1(T13946_Q));
KC_OAI13_X1 T12718 ( .B0(T16245_Y), .A(T2552_Y), .B2(T1108_Y),     .Y(T12718_Y), .B1(T15072_Q));
KC_OAI13_X1 T12691 ( .B0(T7952_Y), .A(T8009_Y), .B2(T1079_Y),     .Y(T12691_Y), .B1(T14611_Q));
KC_OAI13_X1 T12725 ( .B0(T10018_Y), .A(T1493_Y), .B2(T7703_Y),     .Y(T12725_Y), .B1(T1476_Y));
KC_OAI13_X1 T12761 ( .B0(T2065_Y), .A(T5979_Y), .B2(T4868_Y),     .Y(T12761_Y), .B1(T16266_Y));
KC_OAI13_X1 T12751 ( .B0(T13121_Y), .A(T1366_Y), .B2(T10156_Y),     .Y(T12751_Y), .B1(T10936_Y));
KC_OAI13_X1 T12858 ( .B0(T12854_Y), .A(T2879_Y), .B2(T10595_Y),     .Y(T12858_Y), .B1(T13175_Y));
KC_OAI13_X1 T12870 ( .B0(T10996_Y), .A(T16140_Y), .B2(T3394_Y),     .Y(T12870_Y), .B1(T5046_Y));
KC_OAI13_X1 T12910 ( .B0(T6481_Y), .A(T10878_Y), .B2(T6468_Y),     .Y(T12910_Y), .B1(T13583_Q));
KC_AO22BB_X1 T12607 ( .D(T794_Y), .A(T382_Y), .C(T8136_Y), .B(T8679_Y),     .Y(T12607_Y));
KC_AO22BB_X1 T12526 ( .D(T6485_Y), .A(T675_Y), .C(T557_Y), .B(T6485_Y),     .Y(T12526_Y));
KC_AO22BB_X1 T12721 ( .D(T8946_Y), .A(T8064_Y), .C(T1197_Y),     .B(T8037_Y), .Y(T12721_Y));
KC_AO22BB_X1 T12613 ( .D(T1127_Q), .A(T7636_Y), .C(T498_Y),     .B(T12603_Y), .Y(T12613_Y));
KC_AO22BB_X1 T12706 ( .D(T1089_Y), .A(T1092_Q), .C(T1100_Q),     .B(T15466_Y), .Y(T12706_Y));
KC_AO22BB_X1 T12642 ( .D(T7799_Y), .A(T9926_Y), .C(T15472_Y),     .B(T1185_Q), .Y(T12642_Y));
KC_AO22BB_X1 T12641 ( .D(T7799_Y), .A(T10326_Y), .C(T15663_Y),     .B(T1183_Q), .Y(T12641_Y));
KC_AO22BB_X1 T12620 ( .D(T10331_Y), .A(T9926_Y), .C(T15472_Y),     .B(T1186_Q), .Y(T12620_Y));
KC_AO22BB_X1 T12619 ( .D(T10331_Y), .A(T10326_Y), .C(T15663_Y),     .B(T1184_Q), .Y(T12619_Y));
KC_AO22BB_X1 T12901 ( .D(T10329_Y), .A(T10326_Y), .C(T15663_Y),     .B(T4869_Q), .Y(T12901_Y));
KC_AO22BB_X1 T12900 ( .D(T10329_Y), .A(T10327_Y), .C(T16400_Y),     .B(T1190_Q), .Y(T12900_Y));
KC_AO22BB_X1 T12705 ( .D(T7799_Y), .A(T10327_Y), .C(T16400_Y),     .B(T1189_Q), .Y(T12705_Y));
KC_AO22BB_X1 T12704 ( .D(T10329_Y), .A(T9926_Y), .C(T15472_Y),     .B(T1203_Q), .Y(T12704_Y));
KC_AO22BB_X1 T12703 ( .D(T10328_Y), .A(T9926_Y), .C(T15472_Y),     .B(T1215_Q), .Y(T12703_Y));
KC_AO22BB_X1 T12915 ( .D(T2492_Y), .A(T2474_Y), .C(T11016_Y),     .B(T5236_Y), .Y(T12915_Y));
KC_AO22BB_X1 T12914 ( .D(T2492_Y), .A(T2474_Y), .C(T10907_Y),     .B(T1326_Y), .Y(T12914_Y));
KC_AO22BB_X1 T12503 ( .D(T2492_Y), .A(T2474_Y), .C(T10906_Y),     .B(T1333_Y), .Y(T12503_Y));
KC_AO22BB_X1 T12502 ( .D(T2492_Y), .A(T2474_Y), .C(T10883_Y),     .B(T1331_Y), .Y(T12502_Y));
KC_AO22BB_X1 T12640 ( .D(T10261_Y), .A(T1571_Y), .C(T10916_Y),     .B(T1470_Y), .Y(T12640_Y));
KC_AO22BB_X1 T12639 ( .D(T10261_Y), .A(T1571_Y), .C(T15032_Y),     .B(T1351_Y), .Y(T12639_Y));
KC_AO22BB_X1 T12626 ( .D(T10261_Y), .A(T1571_Y), .C(T14987_Y),     .B(T1475_Y), .Y(T12626_Y));
KC_AO22BB_X1 T12624 ( .D(T10261_Y), .A(T1571_Y), .C(T11011_Y),     .B(T5295_Y), .Y(T12624_Y));
KC_AO22BB_X1 T12897 ( .D(T10254_Y), .A(T1571_Y), .C(T15032_Y),     .B(T1478_Y), .Y(T12897_Y));
KC_AO22BB_X1 T12686 ( .D(T10254_Y), .A(T1571_Y), .C(T10916_Y),     .B(T1486_Y), .Y(T12686_Y));
KC_AO22BB_X1 T12680 ( .D(T10254_Y), .A(T1571_Y), .C(T14989_Y),     .B(T1355_Y), .Y(T12680_Y));
KC_AO22BB_X1 T12917 ( .D(T2492_Y), .A(T2474_Y), .C(T10912_Y),     .B(T1411_Y), .Y(T12917_Y));
KC_AO22BB_X1 T12916 ( .D(T2492_Y), .A(T2474_Y), .C(T14989_Y),     .B(T1414_Y), .Y(T12916_Y));
KC_AO22BB_X1 T12922 ( .D(T10261_Y), .A(T2474_Y), .C(T10884_Y),     .B(T1447_Y), .Y(T12922_Y));
KC_AO22BB_X1 T12546 ( .D(T2492_Y), .A(T2474_Y), .C(T15032_Y),     .B(T1413_Y), .Y(T12546_Y));
KC_AO22BB_X1 T12543 ( .D(T10261_Y), .A(T2474_Y), .C(T10907_Y),     .B(T1441_Y), .Y(T12543_Y));
KC_AO22BB_X1 T12539 ( .D(T2492_Y), .A(T2474_Y), .C(T11011_Y),     .B(T1432_Y), .Y(T12539_Y));
KC_AO22BB_X1 T12538 ( .D(T10261_Y), .A(T2474_Y), .C(T10905_Y),     .B(T1443_Y), .Y(T12538_Y));
KC_AO22BB_X1 T12537 ( .D(T10261_Y), .A(T2474_Y), .C(T10883_Y),     .B(T1444_Y), .Y(T12537_Y));
KC_AO22BB_X1 T12535 ( .D(T2492_Y), .A(T2474_Y), .C(T14990_Y),     .B(T1434_Y), .Y(T12535_Y));
KC_AO22BB_X1 T12531 ( .D(T2492_Y), .A(T2474_Y), .C(T10917_Y),     .B(T1433_Y), .Y(T12531_Y));
KC_AO22BB_X1 T12530 ( .D(T2492_Y), .A(T2474_Y), .C(T11010_Y),     .B(T1436_Y), .Y(T12530_Y));
KC_AO22BB_X1 T12629 ( .D(T10261_Y), .A(T1571_Y), .C(T10906_Y),     .B(T1461_Y), .Y(T12629_Y));
KC_AO22BB_X1 T12689 ( .D(T10254_Y), .A(T1571_Y), .C(T10906_Y),     .B(T1489_Y), .Y(T12689_Y));
KC_AO22BB_X1 T12688 ( .D(T10254_Y), .A(T1571_Y), .C(T11010_Y),     .B(T1490_Y), .Y(T12688_Y));
KC_AO22BB_X1 T12684 ( .D(T10254_Y), .A(T1571_Y), .C(T10884_Y),     .B(T1488_Y), .Y(T12684_Y));
KC_AO22BB_X1 T12683 ( .D(T10254_Y), .A(T1571_Y), .C(T10907_Y),     .B(T5338_Y), .Y(T12683_Y));
KC_AO22BB_X1 T12679 ( .D(T10254_Y), .A(T1571_Y), .C(T10883_Y),     .B(T1580_Y), .Y(T12679_Y));
KC_AO22BB_X1 T12617 ( .D(T10254_Y), .A(T2475_Y), .C(T10912_Y),     .B(T4899_Y), .Y(T12617_Y));
KC_AO22BB_X1 T12685 ( .D(T10254_Y), .A(T1571_Y), .C(T10918_Y),     .B(T1583_Y), .Y(T12685_Y));
KC_AO22BB_X1 T12682 ( .D(T10254_Y), .A(T10195_Y), .C(T11016_Y),     .B(T1582_Y), .Y(T12682_Y));
KC_AO22BB_X1 T12681 ( .D(T10254_Y), .A(T10195_Y), .C(T10905_Y),     .B(T1581_Y), .Y(T12681_Y));
KC_AO22BB_X1 T12918 ( .D(T14989_Y), .A(T2491_Y), .C(T4985_Y),     .B(T10406_Y), .Y(T12918_Y));
KC_AO22BB_X1 T12572 ( .D(T2477_Y), .A(T2450_Y), .C(T14990_Y),     .B(T9686_Y), .Y(T12572_Y));
KC_AO22BB_X1 T12555 ( .D(T10916_Y), .A(T2491_Y), .C(T4985_Y),     .B(T8535_Y), .Y(T12555_Y));
KC_AO22BB_X1 T12540 ( .D(T14987_Y), .A(T2491_Y), .C(T4985_Y),     .B(T10408_Y), .Y(T12540_Y));
KC_AO22BB_X1 T12534 ( .D(T11011_Y), .A(T2491_Y), .C(T4985_Y),     .B(T10407_Y), .Y(T12534_Y));
KC_AO22BB_X1 T12533 ( .D(T14987_Y), .A(T2491_Y), .C(T2477_Y),     .B(T9657_Y), .Y(T12533_Y));
KC_AO22BB_X1 T12532 ( .D(T15032_Y), .A(T2491_Y), .C(T4985_Y),     .B(T8534_Y), .Y(T12532_Y));
KC_AO22BB_X1 T12528 ( .D(T14989_Y), .A(T2491_Y), .C(T2477_Y),     .B(T9604_Y), .Y(T12528_Y));
KC_AO22BB_X1 T12583 ( .D(T10261_Y), .A(T2491_Y), .C(T14989_Y),     .B(T15419_Y), .Y(T12583_Y));
KC_AO22BB_X1 T12815 ( .D(T5928_Y), .A(T11502_Y), .C(T1850_Y),     .B(T1285_Y), .Y(T12815_Y));
KC_AO22BB_X1 T12929 ( .D(T2477_Y), .A(T2450_Y), .C(T10912_Y),     .B(T9679_Y), .Y(T12929_Y));
KC_AO22BB_X1 T12949 ( .D(T10917_Y), .A(T2491_Y), .C(T4985_Y),     .B(T9646_Y), .Y(T12949_Y));
KC_AO22BB_X1 T12948 ( .D(T11010_Y), .A(T2491_Y), .C(T4985_Y),     .B(T8532_Y), .Y(T12948_Y));
KC_AO22BB_X1 T12947 ( .D(T10907_Y), .A(T2491_Y), .C(T4985_Y),     .B(T8527_Y), .Y(T12947_Y));
KC_AO22BB_X1 T12946 ( .D(T10906_Y), .A(T2491_Y), .C(T4985_Y),     .B(T8531_Y), .Y(T12946_Y));
KC_AO22BB_X1 T12573 ( .D(T2477_Y), .A(T2450_Y), .C(T10905_Y),     .B(T9678_Y), .Y(T12573_Y));
KC_AO22BB_X1 T12570 ( .D(T2477_Y), .A(T2450_Y), .C(T11011_Y),     .B(T9681_Y), .Y(T12570_Y));
KC_AO22BB_X1 T12569 ( .D(T2477_Y), .A(T2450_Y), .C(T11016_Y),     .B(T9677_Y), .Y(T12569_Y));
KC_AO22BB_X1 T12554 ( .D(T10905_Y), .A(T2491_Y), .C(T4985_Y),     .B(T8530_Y), .Y(T12554_Y));
KC_AO22BB_X1 T12551 ( .D(T2477_Y), .A(T2450_Y), .C(T10918_Y),     .B(T9680_Y), .Y(T12551_Y));
KC_AO22BB_X1 T12935 ( .D(T10912_Y), .A(T2491_Y), .C(T4985_Y),     .B(T10477_Y), .Y(T12935_Y));
KC_AO22BB_X1 T12594 ( .D(T10918_Y), .A(T2491_Y), .C(T4985_Y),     .B(T10478_Y), .Y(T12594_Y));
KC_AO22BB_X1 T12593 ( .D(T11016_Y), .A(T2450_Y), .C(T4985_Y),     .B(T10474_Y), .Y(T12593_Y));
KC_AO22BB_X1 T12794 ( .D(T2109_Y), .A(T2105_Y), .C(T11489_Y),     .B(T2148_Y), .Y(T12794_Y));
KC_AO22BB_X1 T12813 ( .D(T8238_Y), .A(T1761_Q), .C(T2239_Y),     .B(T16156_Y), .Y(T12813_Y));
KC_AO22BB_X1 T12809 ( .D(T8238_Y), .A(T2385_Q), .C(T6026_Y),     .B(T16156_Y), .Y(T12809_Y));
KC_AO22BB_X1 T12832 ( .D(T2240_Y), .A(T6070_Y), .C(T6000_Y),     .B(T2206_Y), .Y(T12832_Y));
KC_AO22BB_X1 T12863 ( .D(T2334_Y), .A(T8172_Y), .C(T2332_Y),     .B(T2360_Q), .Y(T12863_Y));
KC_AO22BB_X1 T12469 ( .D(T2334_Y), .A(T8172_Y), .C(T5520_Y),     .B(T2361_Q), .Y(T12469_Y));
KC_AO22BB_X1 T12878 ( .D(T6604_Y), .A(T15645_Y), .C(T8171_Y),     .B(T2375_Y), .Y(T12878_Y));
KC_AO22BB_X1 T12928 ( .D(T2477_Y), .A(T2450_Y), .C(T10884_Y),     .B(T10438_Y), .Y(T12928_Y));
KC_AO22BB_X1 T12927 ( .D(T2465_Y), .A(T2450_Y), .C(T10917_Y),     .B(T2440_Y), .Y(T12927_Y));
KC_AO22BB_X1 T12571 ( .D(T2477_Y), .A(T2450_Y), .C(T10906_Y),     .B(T9640_Y), .Y(T12571_Y));
KC_AO22BB_X1 T12568 ( .D(T2465_Y), .A(T2450_Y), .C(T11016_Y),     .B(T9670_Y), .Y(T12568_Y));
KC_AO22BB_X1 T12563 ( .D(T2465_Y), .A(T2450_Y), .C(T10905_Y),     .B(T2453_Y), .Y(T12563_Y));
KC_AO22BB_X1 T12562 ( .D(T2477_Y), .A(T2450_Y), .C(T11010_Y),     .B(T9656_Y), .Y(T12562_Y));
KC_AO22BB_X1 T12561 ( .D(T2477_Y), .A(T2450_Y), .C(T10916_Y),     .B(T9671_Y), .Y(T12561_Y));
KC_AO22BB_X1 T12560 ( .D(T2465_Y), .A(T2475_Y), .C(T10907_Y),     .B(T9653_Y), .Y(T12560_Y));
KC_AO22BB_X1 T12553 ( .D(T2477_Y), .A(T2450_Y), .C(T10917_Y),     .B(T9645_Y), .Y(T12553_Y));
KC_AO22BB_X1 T12550 ( .D(T2465_Y), .A(T2475_Y), .C(T10884_Y),     .B(T2434_Y), .Y(T12550_Y));
KC_AO22BB_X1 T12549 ( .D(T2465_Y), .A(T2475_Y), .C(T10918_Y),     .B(T2435_Y), .Y(T12549_Y));
KC_AO22BB_X1 T12937 ( .D(T10883_Y), .A(T2475_Y), .C(T4985_Y),     .B(T9754_Y), .Y(T12937_Y));
KC_AO22BB_X1 T12602 ( .D(T2508_Y), .A(T2590_Y), .C(T10918_Y),     .B(T634_Y), .Y(T12602_Y));
KC_AO22BB_X1 T12600 ( .D(T10261_Y), .A(T2491_Y), .C(T10917_Y),     .B(T633_Y), .Y(T12600_Y));
KC_AO22BB_X1 T12599 ( .D(T10261_Y), .A(T2491_Y), .C(T10912_Y),     .B(T610_Y), .Y(T12599_Y));
KC_AO22BB_X1 T12598 ( .D(T16265_Y), .A(T2475_Y), .C(T14990_Y),     .B(T9772_Y), .Y(T12598_Y));
KC_AO22BB_X1 T12597 ( .D(T10884_Y), .A(T2491_Y), .C(T4985_Y),     .B(T9753_Y), .Y(T12597_Y));
KC_AO22BB_X1 T12596 ( .D(T10261_Y), .A(T2491_Y), .C(T11016_Y),     .B(T611_Y), .Y(T12596_Y));
KC_AO22BB_X1 T12592 ( .D(T14990_Y), .A(T2491_Y), .C(T4985_Y),     .B(T10475_Y), .Y(T12592_Y));
KC_AO22BB_X1 T12590 ( .D(T2480_Y), .A(T610_Y), .C(T9746_Y),     .B(T9748_Y), .Y(T12590_Y));
KC_AO22BB_X1 T12589 ( .D(T2508_Y), .A(T2475_Y), .C(T11016_Y),     .B(T2493_Y), .Y(T12589_Y));
KC_AO22BB_X1 T12588 ( .D(T2508_Y), .A(T2475_Y), .C(T10884_Y),     .B(T2536_Y), .Y(T12588_Y));
KC_AO22BB_X1 T12676 ( .D(T875_Y), .A(T14994_Y), .C(T15050_Y),     .B(T3108_Y), .Y(T12676_Y));
KC_AO22BB_X1 T12672 ( .D(T875_Y), .A(T14994_Y), .C(T9838_Y),     .B(T3110_Y), .Y(T12672_Y));
KC_AO22BB_X1 T12658 ( .D(T2508_Y), .A(T2475_Y), .C(T10917_Y),     .B(T4904_Y), .Y(T12658_Y));
KC_AO22BB_X1 T12654 ( .D(T2508_Y), .A(T2590_Y), .C(T10883_Y),     .B(T2537_Y), .Y(T12654_Y));
KC_AO22BB_X1 T12653 ( .D(T2508_Y), .A(T2590_Y), .C(T10905_Y),     .B(T2533_Y), .Y(T12653_Y));
KC_AO22BB_X1 T12651 ( .D(T2508_Y), .A(T2590_Y), .C(T10907_Y),     .B(T5317_Y), .Y(T12651_Y));
KC_AO22BB_X1 T12649 ( .D(T2523_Y), .A(T15507_Y), .C(T2543_Y),     .B(T16113_Y), .Y(T12649_Y));
KC_AO22BB_X1 T12748 ( .D(T16244_Y), .A(T2566_Y), .C(T11016_Y),     .B(T2619_Y), .Y(T12748_Y));
KC_AO22BB_X1 T12733 ( .D(T2629_Y), .A(T2631_Q), .C(T10057_Y),     .B(T2583_Q), .Y(T12733_Y));
KC_AO22BB_X1 T12732 ( .D(T15155_Y), .A(T14994_Y), .C(T875_Y),     .B(T3720_Y), .Y(T12732_Y));
KC_AO22BB_X1 T12769 ( .D(T16244_Y), .A(T2566_Y), .C(T10884_Y),     .B(T2646_Y), .Y(T12769_Y));
KC_AO22BB_X1 T12765 ( .D(T16244_Y), .A(T2566_Y), .C(T10883_Y),     .B(T2645_Y), .Y(T12765_Y));
KC_AO22BB_X1 T12764 ( .D(T16244_Y), .A(T2566_Y), .C(T10912_Y),     .B(T2647_Y), .Y(T12764_Y));
KC_AO22BB_X1 T12760 ( .D(T16244_Y), .A(T2566_Y), .C(T10905_Y),     .B(T2650_Y), .Y(T12760_Y));
KC_AO22BB_X1 T12759 ( .D(T16244_Y), .A(T2566_Y), .C(T10918_Y),     .B(T2644_Y), .Y(T12759_Y));
KC_AO22BB_X1 T12784 ( .D(T5741_Y), .A(T10249_Y), .C(T5747_Y),     .B(T14490_Q), .Y(T12784_Y));
KC_AO22BB_X1 T12802 ( .D(T3860_Y), .A(T5791_Y), .C(T10245_Y),     .B(T9162_Y), .Y(T12802_Y));
KC_AO22BB_X1 T12831 ( .D(T15881_Y), .A(T12263_Y), .C(T12001_Y),     .B(T8481_Y), .Y(T12831_Y));
KC_AO22BB_X1 T12853 ( .D(T3482_Y), .A(T15234_Y), .C(T3426_Y),     .B(T16167_Y), .Y(T12853_Y));
KC_AO22BB_X1 T12849 ( .D(T3436_Y), .A(T12065_Y), .C(T3526_Y),     .B(T2867_Y), .Y(T12849_Y));
KC_AO22BB_X1 T12874 ( .D(T6101_Y), .A(T8352_Q), .C(T6583_Y),     .B(T10995_Y), .Y(T12874_Y));
KC_AO22BB_X1 T12873 ( .D(T2888_Y), .A(T3517_Y), .C(T10999_Y),     .B(T11698_Y), .Y(T12873_Y));
KC_AO22BB_X1 T12566 ( .D(T2465_Y), .A(T2475_Y), .C(T10906_Y),     .B(T5081_Y), .Y(T12566_Y));
KC_AO22BB_X1 T12565 ( .D(T2465_Y), .A(T2475_Y), .C(T11011_Y),     .B(T9668_Y), .Y(T12565_Y));
KC_AO22BB_X1 T12558 ( .D(T2465_Y), .A(T2475_Y), .C(T11010_Y),     .B(T3023_Y), .Y(T12558_Y));
KC_AO22BB_X1 T12557 ( .D(T2465_Y), .A(T2475_Y), .C(T10916_Y),     .B(T9654_Y), .Y(T12557_Y));
KC_AO22BB_X1 T12934 ( .D(T2465_Y), .A(T2475_Y), .C(T14990_Y),     .B(T10472_Y), .Y(T12934_Y));
KC_AO22BB_X1 T12930 ( .D(T2465_Y), .A(T2475_Y), .C(T14989_Y),     .B(T8526_Y), .Y(T12930_Y));
KC_AO22BB_X1 T12976 ( .D(T2508_Y), .A(T2590_Y), .C(T14989_Y),     .B(T3074_Y), .Y(T12976_Y));
KC_AO22BB_X1 T12674 ( .D(T16244_Y), .A(T2590_Y), .C(T14989_Y),     .B(T5079_Y), .Y(T12674_Y));
KC_AO22BB_X1 T12673 ( .D(T16244_Y), .A(T2590_Y), .C(T14987_Y),     .B(T9839_Y), .Y(T12673_Y));
KC_AO22BB_X1 T12652 ( .D(T16265_Y), .A(T2590_Y), .C(T14989_Y),     .B(T5316_Y), .Y(T12652_Y));
KC_AO22BB_X1 T12648 ( .D(T2508_Y), .A(T2590_Y), .C(T10906_Y),     .B(T3077_Y), .Y(T12648_Y));
KC_AO22BB_X1 T12647 ( .D(T2508_Y), .A(T2590_Y), .C(T14987_Y),     .B(T9878_Y), .Y(T12647_Y));
KC_AO22BB_X1 T12940 ( .D(T2508_Y), .A(T2590_Y), .C(T15032_Y),     .B(T3123_Y), .Y(T12940_Y));
KC_AO22BB_X1 T12939 ( .D(T2508_Y), .A(T2590_Y), .C(T14990_Y),     .B(T3116_Y), .Y(T12939_Y));
KC_AO22BB_X1 T12938 ( .D(T16244_Y), .A(T2590_Y), .C(T14990_Y),     .B(T10507_Y), .Y(T12938_Y));
KC_AO22BB_X1 T12712 ( .D(T2508_Y), .A(T2566_Y), .C(T11010_Y),     .B(T3120_Y), .Y(T12712_Y));
KC_AO22BB_X1 T12711 ( .D(T2508_Y), .A(T2566_Y), .C(T10916_Y),     .B(T3121_Y), .Y(T12711_Y));
KC_AO22BB_X1 T12710 ( .D(T2508_Y), .A(T2566_Y), .C(T11011_Y),     .B(T3119_Y), .Y(T12710_Y));
KC_AO22BB_X1 T12707 ( .D(T16244_Y), .A(T2590_Y), .C(T15032_Y),     .B(T3118_Y), .Y(T12707_Y));
KC_AO22BB_X1 T12743 ( .D(T16244_Y), .A(T2566_Y), .C(T10907_Y),     .B(T3148_Y), .Y(T12743_Y));
KC_AO22BB_X1 T12739 ( .D(T16244_Y), .A(T2566_Y), .C(T11011_Y),     .B(T3147_Y), .Y(T12739_Y));
KC_AO22BB_X1 T12731 ( .D(T16244_Y), .A(T2566_Y), .C(T10916_Y),     .B(T3157_Y), .Y(T12731_Y));
KC_AO22BB_X1 T12767 ( .D(T16244_Y), .A(T2566_Y), .C(T11010_Y),     .B(T2649_Y), .Y(T12767_Y));
KC_AO22BB_X1 T12783 ( .D(T15548_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14492_Q), .Y(T12783_Y));
KC_AO22BB_X1 T12781 ( .D(T5740_Y), .A(T10249_Y), .C(T5747_Y),     .B(T14496_Q), .Y(T12781_Y));
KC_AO22BB_X1 T12780 ( .D(T5734_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14476_Q), .Y(T12780_Y));
KC_AO22BB_X1 T12779 ( .D(T15688_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14491_Q), .Y(T12779_Y));
KC_AO22BB_X1 T12778 ( .D(T5738_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14493_Q), .Y(T12778_Y));
KC_AO22BB_X1 T12777 ( .D(T5729_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14464_Q), .Y(T12777_Y));
KC_AO22BB_X1 T12776 ( .D(T15550_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14475_Q), .Y(T12776_Y));
KC_AO22BB_X1 T12775 ( .D(T5736_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14474_Q), .Y(T12775_Y));
KC_AO22BB_X1 T12774 ( .D(T5706_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14478_Q), .Y(T12774_Y));
KC_AO22BB_X1 T12773 ( .D(T5704_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14462_Q), .Y(T12773_Y));
KC_AO22BB_X1 T12772 ( .D(T15546_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14522_Q), .Y(T12772_Y));
KC_AO22BB_X1 T12854 ( .D(T3445_Y), .A(T15621_Y), .C(T3429_Y),     .B(T8510_Y), .Y(T12854_Y));
KC_AO22BB_X1 T12465 ( .D(T6080_Y), .A(T10583_Y), .C(T3458_Y),     .B(T10585_Y), .Y(T12465_Y));
KC_AO22BB_X1 T12971 ( .D(T8407_Y), .A(T12317_Y), .C(T2888_Y),     .B(T11682_Y), .Y(T12971_Y));
KC_AO22BB_X1 T12956 ( .D(T3789_Y), .A(T11379_Y), .C(T3840_Y),     .B(T11977_Y), .Y(T12956_Y));
KC_AO22BB_X1 T12793 ( .D(T3841_Y), .A(T5830_Y), .C(T5780_Y),     .B(T11317_Y), .Y(T12793_Y));
KC_AO22BB_X1 T12816 ( .D(T3880_Y), .A(T15580_Y), .C(T11519_Y),     .B(T3882_Y), .Y(T12816_Y));
KC_AO22BB_X1 T12473 ( .D(T9563_Y), .A(T4191_Y), .C(T6438_Y),     .B(T9563_Y), .Y(T12473_Y));
KC_AO22BB_X1 T12787 ( .D(T4399_Y), .A(T11393_Y), .C(T14942_Q),     .B(T4396_Y), .Y(T12787_Y));
KC_AO22BB_X1 T12786 ( .D(T5746_Y), .A(T5746_Y), .C(T6031_S),     .B(T15554_Y), .Y(T12786_Y));
KC_AO22BB_X1 T12799 ( .D(T4388_Y), .A(T5838_Y), .C(T5822_Y),     .B(T4446_Y), .Y(T12799_Y));
KC_AO22BB_X1 T12850 ( .D(T8398_Y), .A(T4717_Q), .C(T15757_Y),     .B(T10600_Y), .Y(T12850_Y));
KC_AO22BB_X1 T12844 ( .D(T6420_S), .A(T12298_Y), .C(T12298_Y),     .B(T4737_Y), .Y(T12844_Y));
KC_AO22BB_X1 T12859 ( .D(T6187_Y), .A(T4741_Y), .C(T8406_Y),     .B(T12844_Y), .Y(T12859_Y));
KC_AO22BB_X1 T12905 ( .D(T10331_Y), .A(T10327_Y), .C(T16400_Y),     .B(T1187_Q), .Y(T12905_Y));
KC_AO22BB_X1 T12904 ( .D(T15471_Y), .A(T4861_Q), .C(T1100_Q),     .B(T15466_Y), .Y(T12904_Y));
KC_AO22BB_X1 T12903 ( .D(T10328_Y), .A(T10326_Y), .C(T15663_Y),     .B(T1188_Q), .Y(T12903_Y));
KC_AO22BB_X1 T12902 ( .D(T10328_Y), .A(T10327_Y), .C(T16400_Y),     .B(T1202_Q), .Y(T12902_Y));
KC_AO22BB_X1 T12913 ( .D(T2492_Y), .A(T2474_Y), .C(T14987_Y),     .B(T1435_Y), .Y(T12913_Y));
KC_AO22BB_X1 T12912 ( .D(T2492_Y), .A(T2474_Y), .C(T10884_Y),     .B(T1332_Y), .Y(T12912_Y));
KC_AO22BB_X1 T12899 ( .D(T10254_Y), .A(T1571_Y), .C(T14990_Y),     .B(T4890_Y), .Y(T12899_Y));
KC_AO22BB_X1 T12898 ( .D(T10254_Y), .A(T1571_Y), .C(T14987_Y),     .B(T4880_Y), .Y(T12898_Y));
KC_AO22BB_X1 T12911 ( .D(T2492_Y), .A(T2475_Y), .C(T10918_Y),     .B(T1412_Y), .Y(T12911_Y));
KC_AO22BB_X1 T12894 ( .D(T10254_Y), .A(T1571_Y), .C(T10917_Y),     .B(T4891_Y), .Y(T12894_Y));
KC_AO22BB_X1 T12962 ( .D(T11032_Y), .A(T11551_Y), .C(T6101_Y),     .B(T8181_Y), .Y(T12962_Y));
KC_AO22BB_X1 T12958 ( .D(T11032_Y), .A(T15232_Y), .C(T16130_Y),     .B(T16073_Y), .Y(T12958_Y));
KC_AO22BB_X1 T12926 ( .D(T2477_Y), .A(T2450_Y), .C(T10883_Y),     .B(T9641_Y), .Y(T12926_Y));
KC_AO22BB_X1 T12925 ( .D(T2465_Y), .A(T2450_Y), .C(T10883_Y),     .B(T9639_Y), .Y(T12925_Y));
KC_AO22BB_X1 T12924 ( .D(T2465_Y), .A(T2450_Y), .C(T10912_Y),     .B(T2436_Y), .Y(T12924_Y));
KC_AO22BB_X1 T12961 ( .D(T5068_Y), .A(T3991_Y), .C(T6776_Co),     .B(T6776_S), .Y(T12961_Y));
KC_AO22BB_X1 T12944 ( .D(T13125_Y), .A(T2566_Y), .C(T2632_Y),     .B(T14951_Q), .Y(T12944_Y));
KC_AO22BB_X1 T12932 ( .D(T2465_Y), .A(T2475_Y), .C(T14987_Y),     .B(T3022_Y), .Y(T12932_Y));
KC_AO22BB_X1 T12931 ( .D(T2465_Y), .A(T2475_Y), .C(T15032_Y),     .B(T3021_Y), .Y(T12931_Y));
KC_AO22BB_X1 T12952 ( .D(T4452_Y), .A(T15907_Y), .C(T3857_Y),     .B(T11364_Y), .Y(T12952_Y));
KC_AO22BB_X1 T12564 ( .D(T2477_Y), .A(T2450_Y), .C(T10907_Y),     .B(T9672_Y), .Y(T12564_Y));
KC_AO22BB_X1 T12552 ( .D(T15032_Y), .A(T2450_Y), .C(T2477_Y),     .B(T10442_Y), .Y(T12552_Y));
KC_AO22BB_X1 T12545 ( .D(T2492_Y), .A(T2474_Y), .C(T10905_Y),     .B(T1424_Y), .Y(T12545_Y));
KC_AO22BB_X1 T12529 ( .D(T2492_Y), .A(T2474_Y), .C(T10916_Y),     .B(T1437_Y), .Y(T12529_Y));
KC_AO22BB_X1 T12595 ( .D(T16265_Y), .A(T2475_Y), .C(T14987_Y),     .B(T2489_Y), .Y(T12595_Y));
KC_AO22BB_X1 T12659 ( .D(T2508_Y), .A(T2475_Y), .C(T10912_Y),     .B(T4903_Y), .Y(T12659_Y));
KC_AO22BB_X1 T12627 ( .D(T10261_Y), .A(T1571_Y), .C(T11010_Y),     .B(T1474_Y), .Y(T12627_Y));
KC_AO22BB_X1 T12625 ( .D(T10261_Y), .A(T1571_Y), .C(T14990_Y),     .B(T1473_Y), .Y(T12625_Y));
KC_AO22BB_X1 T12886 ( .D(T967_Y), .A(T371_Y), .C(T8397_Y), .B(T8665_Y),     .Y(T12886_Y));
KC_AO22BB_X1 T12687 ( .D(T10254_Y), .A(T1571_Y), .C(T11011_Y),     .B(T1494_Y), .Y(T12687_Y));
KC_AO22BB_X1 T12723 ( .D(T254_Y), .A(T393_Y), .C(T15488_Y), .B(T254_Y),     .Y(T12723_Y));
KC_AO22BB_X1 T12766 ( .D(T16244_Y), .A(T2566_Y), .C(T10917_Y),     .B(T10180_Y), .Y(T12766_Y));
KC_AO22BB_X1 T12785 ( .D(T10936_Y), .A(T2566_Y), .C(T2632_Y),     .B(T14514_Q), .Y(T12785_Y));
KC_AO22BB_X1 T12782 ( .D(T15549_Y), .A(T10241_Y), .C(T5747_Y),     .B(T14477_Q), .Y(T12782_Y));
KC_AO22BB_X1 T12827 ( .D(T4991_Y), .A(T2381_Q), .C(T6040_Y),     .B(T16156_Y), .Y(T12827_Y));
KC_AO22BB_X1 T12830 ( .D(T16474_Y), .A(T12263_Y), .C(T12001_Y),     .B(T8258_Y), .Y(T12830_Y));
KC_AO22BB_X1 T12888 ( .D(T9012_Y), .A(T4821_Y), .C(T9012_Y),     .B(T1427_Y), .Y(T12888_Y));
KC_AOI211_X1 T15166 ( .C1(T15169_Y), .Y(T15166_Y), .B(T5624_Y),     .A(T9253_Y), .C0(T5633_Y));
KC_AOI211_X1 T12372 ( .C1(T83_Q), .Y(T12372_Y), .B(T5624_Y),     .A(T8548_Y), .C0(T5185_Q));
KC_AOI211_X1 T12370 ( .C1(T81_Q), .Y(T12370_Y), .B(T8549_Y),     .A(T5624_Y), .C0(T9253_Y));
KC_AOI211_X1 T12377 ( .C1(T15324_Y), .Y(T12377_Y), .B(T5624_Y),     .A(T8564_Y), .C0(T5634_Y));
KC_AOI211_X1 T12376 ( .C1(T127_Y), .Y(T12376_Y), .B(T15841_Y),     .A(T8537_Y), .C0(T119_Y));
KC_AOI211_X1 T12384 ( .C1(T9289_Y), .Y(T12384_Y), .B(T6934_Y),     .A(T133_Q), .C0(T9291_Y));
KC_AOI211_X1 T16316 ( .C1(T13241_Q), .Y(T16316_Y), .B(T15841_Y),     .A(T7698_Y), .C0(T8705_Y));
KC_AOI211_X1 T1364 ( .C1(T8993_S), .Y(T1364_Y), .B(T248_Y),     .A(T8992_Y), .C0(T8993_Co));
KC_AOI211_X1 T12373 ( .C1(T280_Y), .Y(T12373_Y), .B(T6859_Y),     .A(T275_Q), .C0(T433_Y));
KC_AOI211_X1 T12403 ( .C1(T9351_Q), .Y(T12403_Y), .B(T7275_Y),     .A(T340_Y), .C0(T569_Y));
KC_AOI211_X1 T16324 ( .C1(T7570_Y), .Y(T16324_Y), .B(T9385_Y),     .A(T16326_Y), .C0(T16331_Y));
KC_AOI211_X1 T1329 ( .C1(T7857_Y), .Y(T1329_Y), .B(T8965_Y),     .A(T8097_Y), .C0(T1334_Y));
KC_AOI211_X1 T12455 ( .C1(T1334_Y), .Y(T12455_Y), .B(T13253_Y),     .A(T13256_Y), .C0(T7909_Y));
KC_AOI211_X1 T12402 ( .C1(T15434_Y), .Y(T12402_Y), .B(T7397_Y),     .A(T11869_Y), .C0(T7421_Y));
KC_AOI211_X1 T12441 ( .C1(T529_Q), .Y(T12441_Y), .B(T16313_Y),     .A(T8751_Y), .C0(T915_Y));
KC_AOI211_X1 T12448 ( .C1(T9269_Y), .Y(T12448_Y), .B(T11230_Y),     .A(T15841_Y), .C0(T7844_Y));
KC_AOI211_X1 T12447 ( .C1(T933_Y), .Y(T12447_Y), .B(T538_Y),     .A(T8810_Y), .C0(T1095_Q));
KC_AOI211_X1 T16186 ( .C1(T9478_Y), .Y(T16186_Y), .B(T4814_Y),     .A(T9166_Y), .C0(T16187_Y));
KC_AOI211_X1 T12375 ( .C1(T5194_Q), .Y(T12375_Y), .B(T109_Y),     .A(T6861_Y), .C0(T108_Y));
KC_AOI211_X1 T12374 ( .C1(T621_Q), .Y(T12374_Y), .B(T9293_Y),     .A(T9292_Y), .C0(T15331_Y));
KC_AOI211_X1 T6272 ( .C1(T812_Q), .Y(T6272_Y), .B(T9274_Y), .A(T299_Y),     .C0(T15355_Y));
KC_AOI211_X1 T6270 ( .C1(T847_Q), .Y(T6270_Y), .B(T9263_Y),     .A(T9264_Y), .C0(T6288_Y));
KC_AOI211_X1 T12388 ( .C1(T446_Q), .Y(T12388_Y), .B(T15350_Y),     .A(T6965_Y), .C0(T250_Y));
KC_AOI211_X1 T12386 ( .C1(T5223_Q), .Y(T12386_Y), .B(T242_Y),     .A(T6942_Y), .C0(T249_Y));
KC_AOI211_X1 T12385 ( .C1(T649_Q), .Y(T12385_Y), .B(T8585_Y),     .A(T8593_Y), .C0(T15171_Y));
KC_AOI211_X1 T12381 ( .C1(T817_Q), .Y(T12381_Y), .B(T8571_Y),     .A(T8570_Y), .C0(T6289_Y));
KC_AOI211_X1 T12380 ( .C1(T5227_Q), .Y(T12380_Y), .B(T302_Y),     .A(T6943_Y), .C0(T304_Y));
KC_AOI211_X1 T12378 ( .C1(T5229_Q), .Y(T12378_Y), .B(T8566_Y),     .A(T8565_Y), .C0(T15349_Y));
KC_AOI211_X1 T6330 ( .C1(T4845_Q), .Y(T6330_Y), .B(T15648_Y),     .A(T7096_Y), .C0(T6332_Y));
KC_AOI211_X1 T12392 ( .C1(T653_Q), .Y(T12392_Y), .B(T8618_Y),     .A(T8617_Y), .C0(T333_Y));
KC_AOI211_X1 T12391 ( .C1(T5240_Q), .Y(T12391_Y), .B(T15367_Y),     .A(T7083_Y), .C0(T6266_Y));
KC_AOI211_X1 T12395 ( .C1(T7086_Y), .Y(T12395_Y), .B(T557_Y),     .A(T8643_Y), .C0(T6485_Y));
KC_AOI211_X1 T12438 ( .C1(T757_Y), .Y(T12438_Y), .B(T7366_Y),     .A(T7416_Y), .C0(T7653_Y));
KC_AOI211_X1 T12437 ( .C1(T8895_Y), .Y(T12437_Y), .B(T7565_Y),     .A(T11204_Y), .C0(T513_Y));
KC_AOI211_X1 T12456 ( .C1(T9242_Y), .Y(T12456_Y), .B(T12749_Y),     .A(T908_Y), .C0(T8066_Y));
KC_AOI211_X1 T12393 ( .C1(T16510_Y), .Y(T12393_Y), .B(T11085_Y),     .A(T4853_Y), .C0(T6250_Y));
KC_AOI211_X1 T6744 ( .C1(T9334_Y), .Y(T6744_Y), .B(T13273_Y),     .A(T734_Y), .C0(T7623_Y));
KC_AOI211_X1 T6743 ( .C1(T12401_Y), .Y(T6743_Y), .B(T13285_Y),     .A(T734_Y), .C0(T7623_Y));
KC_AOI211_X1 T6739 ( .C1(T12401_Y), .Y(T6739_Y), .B(T13272_Y),     .A(T734_Y), .C0(T15031_Y));
KC_AOI211_X1 T6738 ( .C1(T9334_Y), .Y(T6738_Y), .B(T13286_Y),     .A(T734_Y), .C0(T15031_Y));
KC_AOI211_X1 T6735 ( .C1(T9312_Y), .Y(T6735_Y), .B(T13275_Y),     .A(T734_Y), .C0(T15031_Y));
KC_AOI211_X1 T6734 ( .C1(T6805_Y), .Y(T6734_Y), .B(T13274_Y),     .A(T734_Y), .C0(T15031_Y));
KC_AOI211_X1 T6733 ( .C1(T6805_Y), .Y(T6733_Y), .B(T13287_Y),     .A(T734_Y), .C0(T7623_Y));
KC_AOI211_X1 T15748 ( .C1(T9507_Y), .Y(T15748_Y), .B(T10345_Y),     .A(T652_Y), .C0(T927_Y));
KC_AOI211_X1 T15744 ( .C1(T547_Y), .Y(T15744_Y), .B(T13233_Y),     .A(T5352_Y), .C0(T1724_Y));
KC_AOI211_X1 T12404 ( .C1(T552_Y), .Y(T12404_Y), .B(T15745_Y),     .A(T5352_Y), .C0(T9340_Q));
KC_AOI211_X1 T12397 ( .C1(T545_Y), .Y(T12397_Y), .B(T7435_Y),     .A(T5352_Y), .C0(T695_Q));
KC_AOI211_X1 T12396 ( .C1(T548_Y), .Y(T12396_Y), .B(T7356_Y),     .A(T5352_Y), .C0(T687_Q));
KC_AOI211_X1 T12436 ( .C1(T703_Y), .Y(T12436_Y), .B(T7631_Y),     .A(T5352_Y), .C0(T711_Q));
KC_AOI211_X1 T12434 ( .C1(T8719_Y), .Y(T12434_Y), .B(T652_Y),     .A(T7635_Y), .C0(T927_Y));
KC_AOI211_X1 T12433 ( .C1(T16163_Y), .Y(T12433_Y), .B(T7632_Y),     .A(T5352_Y), .C0(T5300_Q));
KC_AOI211_X1 T12431 ( .C1(T9505_Y), .Y(T12431_Y), .B(T639_Y),     .A(T652_Y), .C0(T927_Y));
KC_AOI211_X1 T12428 ( .C1(T9312_Y), .Y(T12428_Y), .B(T13237_Y),     .A(T734_Y), .C0(T7623_Y));
KC_AOI211_X1 T12422 ( .C1(T9714_Y), .Y(T12422_Y), .B(T7551_Y),     .A(T652_Y), .C0(T927_Y));
KC_AOI211_X1 T12421 ( .C1(T660_Y), .Y(T12421_Y), .B(T7587_Y),     .A(T5352_Y), .C0(T710_Q));
KC_AOI211_X1 T12420 ( .C1(T9504_Y), .Y(T12420_Y), .B(T15428_Y),     .A(T652_Y), .C0(T927_Y));
KC_AOI211_X1 T12445 ( .C1(T926_Y), .Y(T12445_Y), .B(T4353_Y),     .A(T7870_Y), .C0(T958_Y));
KC_AOI211_X1 T12453 ( .C1(T9420_Y), .Y(T12453_Y), .B(T965_Y),     .A(T16006_Y), .C0(T8058_Y));
KC_AOI211_X1 T12452 ( .C1(T953_Y), .Y(T12452_Y), .B(T5608_Y),     .A(T1134_Y), .C0(T15454_Y));
KC_AOI211_X1 T12419 ( .C1(T8683_Y), .Y(T12419_Y), .B(T11154_Y),     .A(T7588_Y), .C0(T7615_Y));
KC_AOI211_X1 T12444 ( .C1(T9915_Y), .Y(T12444_Y), .B(T1100_Q),     .A(T7840_Y), .C0(T15466_Y));
KC_AOI211_X1 T12095 ( .C1(T10169_Y), .Y(T12095_Y), .B(T11281_Y),     .A(T11280_Y), .C0(T8110_Y));
KC_AOI211_X1 T12114 ( .C1(T1174_Y), .Y(T12114_Y), .B(T1164_Y),     .A(T9187_Y), .C0(T15798_Q));
KC_AOI211_X1 T12100 ( .C1(T10106_Y), .Y(T12100_Y), .B(T10093_Y),     .A(T2035_Y), .C0(T15089_Y));
KC_AOI211_X1 T12097 ( .C1(T2625_Q), .Y(T12097_Y), .B(T4972_Y),     .A(T10065_Y), .C0(T10064_Y));
KC_AOI211_X1 T12096 ( .C1(T2625_Q), .Y(T12096_Y), .B(T16367_Y),     .A(T10062_Y), .C0(T12736_Y));
KC_AOI211_X1 T12211 ( .C1(T3411_Y), .Y(T12211_Y), .B(T6790_Y),     .A(T11492_Y), .C0(T16302_Y));
KC_AOI211_X1 T12198 ( .C1(T16156_Y), .Y(T12198_Y), .B(T6790_Y),     .A(T11501_Y), .C0(T5465_Q));
KC_AOI211_X1 T12350 ( .C1(T13127_Q), .Y(T12350_Y), .B(T4955_Y),     .A(T12824_Y), .C0(T12028_Y));
KC_AOI211_X1 T12234 ( .C1(T11551_Y), .Y(T12234_Y), .B(T15975_Y),     .A(T13178_Y), .C0(T8180_Y));
KC_AOI211_X1 T12231 ( .C1(T11551_Y), .Y(T12231_Y), .B(T11583_Y),     .A(T12821_Y), .C0(T8270_Y));
KC_AOI211_X1 T12230 ( .C1(T11551_Y), .Y(T12230_Y), .B(T12021_Y),     .A(T13149_Y), .C0(T15829_Y));
KC_AOI211_X1 T12228 ( .C1(T11551_Y), .Y(T12228_Y), .B(T2199_Y),     .A(T12820_Y), .C0(T11465_Y));
KC_AOI211_X1 T12220 ( .C1(T11551_Y), .Y(T12220_Y), .B(T11584_Y),     .A(T13322_Y), .C0(T2146_Y));
KC_AOI211_X1 T12219 ( .C1(T15232_Y), .Y(T12219_Y), .B(T2205_Y),     .A(T12819_Y), .C0(T2673_Y));
KC_AOI211_X1 T12218 ( .C1(T16270_Y), .Y(T12218_Y), .B(T12020_Y),     .A(T13144_Y), .C0(T2851_Y));
KC_AOI211_X1 T12217 ( .C1(T15232_Y), .Y(T12217_Y), .B(T12823_Y),     .A(T12962_Y), .C0(T16097_Y));
KC_AOI211_X1 T12245 ( .C1(T11613_Y), .Y(T12245_Y), .B(T8298_Y),     .A(T8466_Y), .C0(T2219_Y));
KC_AOI211_X1 T12301 ( .C1(T2355_Q), .Y(T12301_Y), .B(T11755_Y),     .A(T11754_Y), .C0(T11766_Y));
KC_AOI211_X1 T12319 ( .C1(T2956_Y), .Y(T12319_Y), .B(T2386_Y),     .A(T7836_Y), .C0(T2951_Y));
KC_AOI211_X1 T12080 ( .C1(T9745_Y), .Y(T12080_Y), .B(T12590_Y),     .A(T6849_Y), .C0(T9744_Y));
KC_AOI211_X1 T12090 ( .C1(T2957_Y), .Y(T12090_Y), .B(T1988_Y),     .A(T2571_Q), .C0(T15478_Y));
KC_AOI211_X1 T12098 ( .C1(T10526_Y), .Y(T12098_Y), .B(T11285_Y),     .A(T15501_Y), .C0(T2630_Y));
KC_AOI211_X1 T12128 ( .C1(T10278_Y), .Y(T12128_Y), .B(T10251_Y),     .A(T11960_Y), .C0(T5749_Y));
KC_AOI211_X1 T12334 ( .C1(T10243_Y), .Y(T12334_Y), .B(T4993_Y),     .A(T11963_Y), .C0(T15070_Y));
KC_AOI211_X1 T12141 ( .C1(T11964_Y), .Y(T12141_Y), .B(T10251_Y),     .A(T8187_Y), .C0(T5766_Y));
KC_AOI211_X1 T12136 ( .C1(T5773_Y), .Y(T12136_Y), .B(T15827_Y),     .A(T11960_Y), .C0(T11327_Y));
KC_AOI211_X1 T12155 ( .C1(T16082_Q), .Y(T12155_Y), .B(T2704_Y),     .A(T11431_Y), .C0(T2699_Y));
KC_AOI211_X1 T12189 ( .C1(T2751_Y), .Y(T12189_Y), .B(T2742_Y),     .A(T8234_Y), .C0(T13110_Q));
KC_AOI211_X1 T12203 ( .C1(T11448_Y), .Y(T12203_Y), .B(T15943_Y),     .A(T16302_Y), .C0(T11597_Y));
KC_AOI211_X1 T12291 ( .C1(T12102_Y), .Y(T12291_Y), .B(T2876_Y),     .A(T8503_Y), .C0(T10592_Y));
KC_AOI211_X1 T12285 ( .C1(T2870_Y), .Y(T12285_Y), .B(T16084_Y),     .A(T6144_Y), .C0(T3425_Y));
KC_AOI211_X1 T12275 ( .C1(T6237_Y), .Y(T12275_Y), .B(T2860_Y),     .A(T10604_Y), .C0(T6556_Y));
KC_AOI211_X1 T12267 ( .C1(T10583_Y), .Y(T12267_Y), .B(T11743_Y),     .A(T10589_Y), .C0(T12876_Y));
KC_AOI211_X1 T12266 ( .C1(T6140_Y), .Y(T12266_Y), .B(T3428_Y),     .A(T10552_Y), .C0(T2875_Y));
KC_AOI211_X1 T12259 ( .C1(T3517_Y), .Y(T12259_Y), .B(T3449_Y),     .A(T10569_Y), .C0(T11696_Y));
KC_AOI211_X1 T12312 ( .C1(T8261_Y), .Y(T12312_Y), .B(T2881_Y),     .A(T2897_Y), .C0(T5515_Y));
KC_AOI211_X1 T12311 ( .C1(T8261_Y), .Y(T12311_Y), .B(T4998_Y),     .A(T2891_Y), .C0(T6239_Y));
KC_AOI211_X1 T12306 ( .C1(T2833_Q), .Y(T12306_Y), .B(T2891_Y),     .A(T2900_Y), .C0(T6513_Y));
KC_AOI211_X1 T12305 ( .C1(T2316_Q), .Y(T12305_Y), .B(T3499_Y),     .A(T11782_Y), .C0(T10543_Y));
KC_AOI211_X1 T12296 ( .C1(T6195_Y), .Y(T12296_Y), .B(T11741_Y),     .A(T2865_Y), .C0(T2913_Y));
KC_AOI211_X1 T12126 ( .C1(T14520_Q), .Y(T12126_Y), .B(T10265_Y),     .A(T5748_Y), .C0(T10268_Y));
KC_AOI211_X1 T12147 ( .C1(T11370_Y), .Y(T12147_Y), .B(T5430_Y),     .A(T12148_Y), .C0(T11394_Y));
KC_AOI211_X1 T12146 ( .C1(T5428_Q), .Y(T12146_Y), .B(T11320_Y),     .A(T3201_Y), .C0(T3213_Q));
KC_AOI211_X1 T12140 ( .C1(T11394_Y), .Y(T12140_Y), .B(T3807_Y),     .A(T11319_Y), .C0(T3203_Y));
KC_AOI211_X1 T12135 ( .C1(T10241_Y), .Y(T12135_Y), .B(T11341_Y),     .A(T11960_Y), .C0(T14520_Q));
KC_AOI211_X1 T12131 ( .C1(T11410_Y), .Y(T12131_Y), .B(T15007_Y),     .A(T11319_Y), .C0(T11987_Y));
KC_AOI211_X1 T12168 ( .C1(T14546_Q), .Y(T12168_Y), .B(T11413_Y),     .A(T3855_Y), .C0(T11412_Y));
KC_AOI211_X1 T12201 ( .C1(T3303_Y), .Y(T12201_Y), .B(T11486_Y),     .A(T5890_Y), .C0(T8267_Y));
KC_AOI211_X1 T12240 ( .C1(T6320_Co), .Y(T12240_Y), .B(T7915_Y),     .A(T6335_Y), .C0(T3361_Y));
KC_AOI211_X1 T12254 ( .C1(T6842_S), .Y(T12254_Y), .B(T13160_Y),     .A(T11674_Y), .C0(T3381_Y));
KC_AOI211_X1 T12251 ( .C1(T11647_Y), .Y(T12251_Y), .B(T3410_Y),     .A(T5522_Y), .C0(T3468_Y));
KC_AOI211_X1 T12250 ( .C1(T11661_Y), .Y(T12250_Y), .B(T13161_Y),     .A(T3410_Y), .C0(T5492_Y));
KC_AOI211_X1 T12247 ( .C1(T15233_Y), .Y(T12247_Y), .B(T3395_Y),     .A(T3399_Y), .C0(T6081_Y));
KC_AOI211_X1 T12283 ( .C1(T6158_Y), .Y(T12283_Y), .B(T3461_Y),     .A(T3416_Y), .C0(T12877_Y));
KC_AOI211_X1 T12274 ( .C1(T2839_Y), .Y(T12274_Y), .B(T11694_Y),     .A(T12849_Y), .C0(T13175_Y));
KC_AOI211_X1 T12273 ( .C1(T12043_Y), .Y(T12273_Y), .B(T3441_Y),     .A(T3430_Y), .C0(T12040_Y));
KC_AOI211_X1 T12265 ( .C1(T12043_Y), .Y(T12265_Y), .B(T3440_Y),     .A(T12060_Y), .C0(T3371_Y));
KC_AOI211_X1 T12264 ( .C1(T15711_Y), .Y(T12264_Y), .B(T16136_Y),     .A(T10549_Y), .C0(T3453_Y));
KC_AOI211_X1 T12257 ( .C1(T12043_Y), .Y(T12257_Y), .B(T12057_Y),     .A(T10549_Y), .C0(T3446_Y));
KC_AOI211_X1 T12256 ( .C1(T6100_Y), .Y(T12256_Y), .B(T12846_Y),     .A(T3455_Y), .C0(T10552_Y));
KC_AOI211_X1 T12363 ( .C1(T12317_Y), .Y(T12363_Y), .B(T3462_Y),     .A(T6577_Y), .C0(T4094_Y));
KC_AOI211_X1 T12310 ( .C1(T11831_Y), .Y(T12310_Y), .B(T11797_Y),     .A(T13327_Y), .C0(T11697_Y));
KC_AOI211_X1 T12304 ( .C1(T16102_Y), .Y(T12304_Y), .B(T10990_Y),     .A(T10544_Y), .C0(T4098_Y));
KC_AOI211_X1 T12303 ( .C1(T2345_Q), .Y(T12303_Y), .B(T13188_Y),     .A(T8415_Y), .C0(T10543_Y));
KC_AOI211_X1 T12300 ( .C1(T11818_Y), .Y(T12300_Y), .B(T11800_Y),     .A(T13186_Y), .C0(T6585_Y));
KC_AOI211_X1 T12295 ( .C1(T6590_S), .Y(T12295_Y), .B(T11737_Y),     .A(T3497_Y), .C0(T3498_Y));
KC_AOI211_X1 T12294 ( .C1(T12103_Y), .Y(T12294_Y), .B(T11738_Y),     .A(T11765_Y), .C0(T10553_Y));
KC_AOI211_X1 T12293 ( .C1(T10571_Y), .Y(T12293_Y), .B(T8416_Y),     .A(T11765_Y), .C0(T6610_S));
KC_AOI211_X1 T5769 ( .C1(T15870_Y), .Y(T5769_Y), .B(T12134_Y),     .A(T6041_Y), .C0(T15865_Y));
KC_AOI211_X1 T5755 ( .C1(T15877_Y), .Y(T5755_Y), .B(T8192_Y),     .A(T6053_Y), .C0(T15852_Y));
KC_AOI211_X1 T12145 ( .C1(T11318_Y), .Y(T12145_Y), .B(T3798_Y),     .A(T13077_Y), .C0(T11984_Y));
KC_AOI211_X1 T12139 ( .C1(T11985_Y), .Y(T12139_Y), .B(T12793_Y),     .A(T11352_Y), .C0(T11336_Y));
KC_AOI211_X1 T12138 ( .C1(T4465_Q), .Y(T12138_Y), .B(T13086_Y),     .A(T12792_Y), .C0(T11350_Y));
KC_AOI211_X1 T12130 ( .C1(T11984_Y), .Y(T12130_Y), .B(T13066_Y),     .A(T13077_Y), .C0(T5815_Y));
KC_AOI211_X1 T12158 ( .C1(T16154_Y), .Y(T12158_Y), .B(T15887_Y),     .A(T8197_Y), .C0(T15889_Y));
KC_AOI211_X1 T12185 ( .C1(T3922_Y), .Y(T12185_Y), .B(T3265_Y),     .A(T3868_Y), .C0(T15939_Y));
KC_AOI211_X1 T12205 ( .C1(T11476_Y), .Y(T12205_Y), .B(T3906_Y),     .A(T11590_Y), .C0(T5986_Y));
KC_AOI211_X1 T12200 ( .C1(T11484_Y), .Y(T12200_Y), .B(T13313_Y),     .A(T12814_Y), .C0(T8237_Y));
KC_AOI211_X1 T12227 ( .C1(T3974_Q), .Y(T12227_Y), .B(T15589_Y),     .A(T3964_Q), .C0(T3965_Q));
KC_AOI211_X1 T12226 ( .C1(T15971_Y), .Y(T12226_Y), .B(T15588_Y),     .A(T5984_Y), .C0(T15589_Y));
KC_AOI211_X1 T12225 ( .C1(T5973_Y), .Y(T12225_Y), .B(T11576_Y),     .A(T5984_Y), .C0(T3947_Y));
KC_AOI211_X1 T12213 ( .C1(T5957_Y), .Y(T12213_Y), .B(T3981_Y),     .A(T6352_Y), .C0(T5459_Y));
KC_AOI211_X1 T12239 ( .C1(T15610_Y), .Y(T12239_Y), .B(T16029_Y),     .A(T4042_Y), .C0(T6033_Y));
KC_AOI211_X1 T12246 ( .C1(T12071_Y), .Y(T12246_Y), .B(T16030_Y),     .A(T4037_Y), .C0(T4928_Y));
KC_AOI211_X1 T12289 ( .C1(T16051_Y), .Y(T12289_Y), .B(T8503_Y),     .A(T8502_Y), .C0(T10615_Y));
KC_AOI211_X1 T12288 ( .C1(T4589_Y), .Y(T12288_Y), .B(T13176_Y),     .A(T11727_Y), .C0(T8502_Y));
KC_AOI211_X1 T12286 ( .C1(T10624_Y), .Y(T12286_Y), .B(T3431_Y),     .A(T11712_Y), .C0(T11715_Y));
KC_AOI211_X1 T12280 ( .C1(T4589_Y), .Y(T12280_Y), .B(T6162_Y),     .A(T11636_Y), .C0(T6157_Y));
KC_AOI211_X1 T12279 ( .C1(T6147_Y), .Y(T12279_Y), .B(T12851_Y),     .A(T10604_Y), .C0(T16148_Y));
KC_AOI211_X1 T12278 ( .C1(T10615_Y), .Y(T12278_Y), .B(T13174_Y),     .A(T8502_Y), .C0(T4075_Y));
KC_AOI211_X1 T12272 ( .C1(T10581_Y), .Y(T12272_Y), .B(T13173_Y),     .A(T8386_Y), .C0(T4086_Y));
KC_AOI211_X1 T12262 ( .C1(T10586_Y), .Y(T12262_Y), .B(T8381_Y),     .A(T3459_Y), .C0(T15619_Y));
KC_AOI211_X1 T12255 ( .C1(T11745_Y), .Y(T12255_Y), .B(T4102_Y),     .A(T4087_Y), .C0(T10583_Y));
KC_AOI211_X1 T12116 ( .C1(T4376_Q), .Y(T12116_Y), .B(T10246_Y),     .A(T10257_Y), .C0(T3185_Y));
KC_AOI211_X1 T12143 ( .C1(T11312_Y), .Y(T12143_Y), .B(T11344_Y),     .A(T8178_Y), .C0(T11348_Y));
KC_AOI211_X1 T12137 ( .C1(T11312_Y), .Y(T12137_Y), .B(T12787_Y),     .A(T8178_Y), .C0(T5777_Y));
KC_AOI211_X1 T12129 ( .C1(T5798_Y), .Y(T12129_Y), .B(T11371_Y),     .A(T6742_Y), .C0(T3826_Y));
KC_AOI211_X1 T12173 ( .C1(T14551_Q), .Y(T12173_Y), .B(T12799_Y),     .A(T4431_Y), .C0(T15870_Y));
KC_AOI211_X1 T12172 ( .C1(T5821_Y), .Y(T12172_Y), .B(T11423_Y),     .A(T8195_Y), .C0(T11419_Y));
KC_AOI211_X1 T12156 ( .C1(T11408_Y), .Y(T12156_Y), .B(T13084_Y),     .A(T143_Y), .C0(T11391_Y));
KC_AOI211_X1 T12183 ( .C1(T4477_Y), .Y(T12183_Y), .B(T15934_Y),     .A(T5141_Y), .C0(T12182_Y));
KC_AOI211_X1 T12180 ( .C1(T4479_Y), .Y(T12180_Y), .B(T5846_Y),     .A(T6136_Y), .C0(T4503_Y));
KC_AOI211_X1 T12207 ( .C1(T4534_Y), .Y(T12207_Y), .B(T4507_Y),     .A(T12196_Y), .C0(T12182_Y));
KC_AOI211_X1 T12193 ( .C1(T4528_Q), .Y(T12193_Y), .B(T11475_Y),     .A(T5139_Y), .C0(T15706_Y));
KC_AOI211_X1 T12233 ( .C1(T16013_Y), .Y(T12233_Y), .B(T4554_Y),     .A(T13134_Y), .C0(T4567_Y));
KC_AOI211_X1 T12232 ( .C1(T3870_Y), .Y(T12232_Y), .B(T5986_Y),     .A(T10951_Y), .C0(T6283_Y));
KC_AOI211_X1 T12229 ( .C1(T11572_Y), .Y(T12229_Y), .B(T11573_Y),     .A(T11573_Y), .C0(T11573_Y));
KC_AOI211_X1 T12224 ( .C1(T11574_Y), .Y(T12224_Y), .B(T10951_Y),     .A(T12024_Y), .C0(T4561_Y));
KC_AOI211_X1 T12223 ( .C1(T4514_Y), .Y(T12223_Y), .B(T4553_Y),     .A(T11539_Y), .C0(T5971_Y));
KC_AOI211_X1 T12222 ( .C1(T4561_Y), .Y(T12222_Y), .B(T2757_Y),     .A(T4577_Y), .C0(T8329_Y));
KC_AOI211_X1 T12221 ( .C1(T5971_Y), .Y(T12221_Y), .B(T5980_Y),     .A(T4577_Y), .C0(T4514_Y));
KC_AOI211_X1 T12345 ( .C1(T4688_Y), .Y(T12345_Y), .B(T15132_Y),     .A(T4692_Y), .C0(T16045_Y));
KC_AOI211_X1 T12261 ( .C1(T6102_Y), .Y(T12261_Y), .B(T15757_Y),     .A(T10575_Y), .C0(T6126_Y));
KC_AOI211_X1 T12260 ( .C1(T4720_Q), .Y(T12260_Y), .B(T10574_Y),     .A(T15757_Y), .C0(T10575_Y));
KC_AOI211_X1 T12360 ( .C1(T16146_Y), .Y(T12360_Y), .B(T10541_Y),     .A(T16144_Y), .C0(T12307_Y));
KC_AOI211_X1 T12307 ( .C1(T4750_Q), .Y(T12307_Y), .B(T11788_Y),     .A(T11787_Y), .C0(T4718_Q));
KC_AOI211_X1 T12302 ( .C1(T16145_Y), .Y(T12302_Y), .B(T6244_Y),     .A(T6234_Y), .C0(T6103_Y));
KC_AOI211_X1 T12298 ( .C1(T4749_Y), .Y(T12298_Y), .B(T4750_Q),     .A(T11758_Y), .C0(T6420_Co));
KC_AOI211_X1 T16320 ( .C1(T16331_Y), .Y(T16320_Y), .B(T13282_Y),     .A(T13283_Y), .C0(T7576_Y));
KC_AOI211_X1 T16288 ( .C1(T9085_Y), .Y(T16288_Y), .B(T9021_Y),     .A(T9027_Y), .C0(T9450_Y));
KC_AOI211_X1 T6258 ( .C1(T445_Q), .Y(T6258_Y), .B(T6300_Y),     .A(T6305_Y), .C0(T6264_Y));
KC_AOI211_X1 T15749 ( .C1(T9503_Y), .Y(T15749_Y), .B(T10344_Y),     .A(T652_Y), .C0(T927_Y));
KC_AOI211_X1 T15747 ( .C1(T9506_Y), .Y(T15747_Y), .B(T9332_Y),     .A(T652_Y), .C0(T927_Y));
KC_AOI211_X1 T15743 ( .C1(T6659_Y), .Y(T15743_Y), .B(T15746_Y),     .A(T5352_Y), .C0(T705_Q));
KC_AOI211_X1 T12347 ( .C1(T12009_Y), .Y(T12347_Y), .B(T11619_Y),     .A(T12007_Y), .C0(T8490_Y));
KC_AOI211_X1 T12340 ( .C1(T11499_Y), .Y(T12340_Y), .B(T15943_Y),     .A(T16033_Y), .C0(T11639_Y));
KC_AOI211_X1 T12335 ( .C1(T2655_Y), .Y(T12335_Y), .B(T2662_Y),     .A(T5766_Y), .C0(T10281_Y));
KC_AOI211_X1 T12069 ( .C1(T6545_Y), .Y(T12069_Y), .B(T1_Y),     .A(T6844_Y), .C0(T287_Y));
KC_AOI211_X1 T12364 ( .C1(T5491_Y), .Y(T12364_Y), .B(T5060_Y),     .A(T10552_Y), .C0(T10544_Y));
KC_AOI211_X1 T12358 ( .C1(T6082_Y), .Y(T12358_Y), .B(T13318_Y),     .A(T16104_Y), .C0(T6178_Y));
KC_AOI211_X1 T12333 ( .C1(T11337_Y), .Y(T12333_Y), .B(T15818_Y),     .A(T10239_Y), .C0(T5433_Y));
KC_AOI211_X1 T12362 ( .C1(T16142_Y), .Y(T12362_Y), .B(T10605_Y),     .A(T5116_Y), .C0(T4164_Q));
KC_AOI211_X1 T12361 ( .C1(T10566_Y), .Y(T12361_Y), .B(T13326_Y),     .A(T8385_Y), .C0(T6841_S));
KC_AOI211_X1 T12342 ( .C1(T15845_Y), .Y(T12342_Y), .B(T11389_Y),     .A(T11977_Y), .C0(T16153_Y));
KC_AOI211_X1 T12353 ( .C1(T15938_Y), .Y(T12353_Y), .B(T6194_S),     .A(T5154_Y), .C0(T4531_Y));
KC_AOI211_X1 T12351 ( .C1(T15964_Y), .Y(T12351_Y), .B(T5139_Y),     .A(T12023_Y), .C0(T4519_Y));
KC_AOI211_X1 T12341 ( .C1(T11984_Y), .Y(T12341_Y), .B(T4451_Y),     .A(T13083_Y), .C0(T15875_Y));
KC_AOI211_X1 T12337 ( .C1(T5789_Y), .Y(T12337_Y), .B(T5163_Y),     .A(T4465_Q), .C0(T11965_Y));
KC_AOI211_X1 T12394 ( .C1(T843_Q), .Y(T12394_Y), .B(T8634_Y),     .A(T8612_Y), .C0(T345_Y));
KC_AOI211_X1 T16335 ( .C1(T9387_Y), .Y(T16335_Y), .B(T13240_Y),     .A(T13281_Y), .C0(T12607_Y));
KC_AOI211_X1 T1423 ( .C1(T1427_Y), .Y(T1423_Y), .B(T4829_Y),     .A(T1422_Y), .C0(T1422_Y));
KC_AOI211_X1 T12458 ( .C1(T8082_Y), .Y(T12458_Y), .B(T13254_Y),     .A(T13255_Y), .C0(T12886_Y));
KC_AOI211_X1 T12099 ( .C1(T10070_Y), .Y(T12099_Y), .B(T10094_Y),     .A(T2035_Y), .C0(T15073_Y));
KC_AOI211_X1 T12109 ( .C1(T15999_Y), .Y(T12109_Y), .B(T1149_Y),     .A(T11913_Y), .C0(T10175_Y));
KC_AOI211_X1 T12127 ( .C1(T11337_Y), .Y(T12127_Y), .B(T2660_Y),     .A(T10242_Y), .C0(T3791_Y));
KC_AOI211_X1 T15755 ( .C1(T16160_Y), .Y(T15755_Y), .B(T2668_Y),     .A(T4994_Y), .C0(T11325_Y));
KC_AOI211_X1 T12157 ( .C1(T5795_Y), .Y(T12157_Y), .B(T13304_Y),     .A(T5437_Y), .C0(T15897_Y));
KC_AOI211_X1 T12354 ( .C1(T6219_Y), .Y(T12354_Y), .B(T12356_Y),     .A(T3903_Y), .C0(T3880_Y));
KC_AOI211_X1 T12214 ( .C1(T8289_Y), .Y(T12214_Y), .B(T11575_Y),     .A(T5022_Y), .C0(T15159_Y));
KC_AOI211_X1 T12287 ( .C1(T6178_Y), .Y(T12287_Y), .B(T13168_Y),     .A(T12036_Y), .C0(T11637_Y));
KC_AOI211_X1 T12271 ( .C1(T6842_S), .Y(T12271_Y), .B(T13166_Y),     .A(T12036_Y), .C0(T16125_Y));
KC_AOI211_X1 T12258 ( .C1(T10589_Y), .Y(T12258_Y), .B(T2859_Y),     .A(T10569_Y), .C0(T6193_Y));
KC_AOI211_X1 T12365 ( .C1(T10553_Y), .Y(T12365_Y), .B(T16136_Y),     .A(T10554_Y), .C0(T5523_Y));
KC_AOI211_X1 T12299 ( .C1(T10568_Y), .Y(T12299_Y), .B(T13180_Y),     .A(T2906_Y), .C0(T4609_Y));
KC_AOI211_X1 T12366 ( .C1(T3517_Y), .Y(T12366_Y), .B(T11723_Y),     .A(T10546_Y), .C0(T2852_Y));
KC_AOI211_X1 T12359 ( .C1(T2906_Y), .Y(T12359_Y), .B(T11672_Y),     .A(T3404_Y), .C0(T5491_Y));
KC_AOI211_X1 T12072 ( .C1(T15628_Y), .Y(T12072_Y), .B(T2374_Y),     .A(T6500_Y), .C0(T4978_Y));
KC_AOI32_X1 T11277 ( .B0(T9084_Y), .A0(T16286_Y), .A1(T16283_Y),     .Y(T11277_Y), .A2(T243_Y), .B1(T9030_Y));
KC_AOI32_X1 T11296 ( .B0(T9088_Y), .A0(T15092_Y), .A1(T9086_Y),     .Y(T11296_Y), .A2(T15091_Y), .B1(T9086_Y));
KC_AOI32_X1 T11209 ( .B0(T742_Y), .A0(T7821_Y), .A1(T7667_Y),     .Y(T11209_Y), .A2(T7626_Y), .B1(T7667_Y));
KC_AOI32_X1 T11208 ( .B0(T742_Y), .A0(T7823_Y), .A1(T7664_Y),     .Y(T11208_Y), .A2(T7662_Y), .B1(T7664_Y));
KC_AOI32_X1 T11198 ( .B0(T742_Y), .A0(T7627_Y), .A1(T7665_Y),     .Y(T11198_Y), .A2(T7819_Y), .B1(T7665_Y));
KC_AOI32_X1 T11238 ( .B0(T968_Y), .A0(T7911_Y), .A1(T7862_Y),     .Y(T11238_Y), .A2(T8140_Y), .B1(T7862_Y));
KC_AOI32_X1 T11237 ( .B0(T968_Y), .A0(T8137_Y), .A1(T7861_Y),     .Y(T11237_Y), .A2(T7860_Y), .B1(T7861_Y));
KC_AOI32_X1 T11236 ( .B0(T966_Y), .A0(T7900_Y), .A1(T7845_Y),     .Y(T11236_Y), .A2(T15453_Y), .B1(T7845_Y));
KC_AOI32_X1 T11235 ( .B0(T968_Y), .A0(T8139_Y), .A1(T7873_Y),     .Y(T11235_Y), .A2(T7817_Y), .B1(T7873_Y));
KC_AOI32_X1 T11227 ( .B0(T7628_Y), .A0(T7828_Y), .A1(T16321_Y),     .Y(T11227_Y), .A2(T917_Y), .B1(T16321_Y));
KC_AOI32_X1 T11271 ( .B0(T7858_Y), .A0(T8103_Y), .A1(T8105_Y),     .Y(T11271_Y), .A2(T1273_Y), .B1(T8105_Y));
KC_AOI32_X1 T11266 ( .B0(T7856_Y), .A0(T8916_Y), .A1(T8910_Y),     .Y(T11266_Y), .A2(T7917_Y), .B1(T8910_Y));
KC_AOI32_X1 T11304 ( .B0(T9496_Y), .A0(T9171_Y), .A1(T15525_Y),     .Y(T11304_Y), .A2(T16286_Y), .B1(T9172_Y));
KC_AOI32_X1 T11303 ( .B0(T9484_Y), .A0(T9170_Y), .A1(T16191_Y),     .Y(T11303_Y), .A2(T16286_Y), .B1(T9173_Y));
KC_AOI32_X1 T11294 ( .B0(T15816_Y), .A0(T9117_Y), .A1(T9119_Y),     .Y(T11294_Y), .A2(T9136_Y), .B1(T9119_Y));
KC_AOI32_X1 T11210 ( .B0(T742_Y), .A0(T7820_Y), .A1(T7663_Y),     .Y(T11210_Y), .A2(T7661_Y), .B1(T7663_Y));
KC_AOI32_X1 T11204 ( .B0(T13260_Y), .A0(T5346_Q), .A1(T12604_Y),     .Y(T11204_Y), .A2(T543_Q), .B1(T12604_Y));
KC_AOI32_X1 T11203 ( .B0(T8803_Y), .A0(T5356_Q), .A1(T5296_Y),     .Y(T11203_Y), .A2(T4827_Q), .B1(T5296_Y));
KC_AOI32_X1 T11233 ( .B0(T1095_Q), .A0(T16318_Y), .A1(T12448_Y),     .Y(T11233_Y), .A2(T928_Y), .B1(T12448_Y));
KC_AOI32_X1 T11276 ( .B0(T561_Q), .A0(T567_Q), .A1(T1352_Y),     .Y(T11276_Y), .A2(T8123_Y), .B1(T555_Y));
KC_AOI32_X1 T11273 ( .B0(T567_Q), .A0(T1593_Y), .A1(T1599_Y),     .Y(T11273_Y), .A2(T9418_Y), .B1(T8125_Y));
KC_AOI32_X1 T11272 ( .B0(T8980_Y), .A0(T750_Q), .A1(T8120_Y),     .Y(T11272_Y), .A2(T8116_Y), .B1(T8120_Y));
KC_AOI32_X1 T4806 ( .B0(T1593_Y), .A0(T9469_Q), .A1(T955_Y),     .Y(T4806_Y), .A2(T10140_Y), .B1(T955_Y));
KC_AOI32_X1 T11900 ( .B0(T4813_Y), .A0(T9477_Y), .A1(T16184_Y),     .Y(T11900_Y), .A2(T11306_Y), .B1(T9166_Y));
KC_AOI32_X1 T11301 ( .B0(T5406_Q), .A0(T8123_Y), .A1(T4815_Y),     .Y(T11301_Y), .A2(T9107_Y), .B1(T4806_Y));
KC_AOI32_X1 T11299 ( .B0(T9469_Q), .A0(T8123_Y), .A1(T1841_Y),     .Y(T11299_Y), .A2(T10140_Y), .B1(T599_Y));
KC_AOI32_X1 T11293 ( .B0(T1593_Y), .A0(T605_Q), .A1(T955_Y),     .Y(T11293_Y), .A2(T598_Y), .B1(T955_Y));
KC_AOI32_X1 T11292 ( .B0(T606_Q), .A0(T8123_Y), .A1(T1842_Y),     .Y(T11292_Y), .A2(T9109_Y), .B1(T11293_Y));
KC_AOI32_X1 T11308 ( .B0(T1599_Y), .A0(T216_Y), .A1(T11307_Y),     .Y(T11308_Y), .A2(T16189_Y), .B1(T11307_Y));
KC_AOI32_X1 T11307 ( .B0(T9475_Y), .A0(T16507_Y), .A1(T1352_Y),     .Y(T11307_Y), .A2(T5345_Y), .B1(T561_Q));
KC_AOI32_X1 T11306 ( .B0(T9243_Y), .A0(T605_Q), .A1(T1279_Y),     .Y(T11306_Y), .A2(T15538_Y), .B1(T1279_Y));
KC_AOI32_X1 T11183 ( .B0(T8939_Y), .A0(T725_Q), .A1(T6427_Y),     .Y(T11183_Y), .A2(T713_Q), .B1(T6427_Y));
KC_AOI32_X1 T11218 ( .B0(T930_Y), .A0(T907_Y), .A1(T8794_Y),     .Y(T11218_Y), .A2(T928_Y), .B1(T15454_Y));
KC_AOI32_X1 T11268 ( .B0(T8037_Y), .A0(T9096_Y), .A1(T8901_Y),     .Y(T11268_Y), .A2(T16420_Y), .B1(T8901_Y));
KC_AOI32_X1 T11085 ( .B0(T833_Y), .A0(T6250_Y), .A1(T16510_Y),     .Y(T11085_Y), .A2(T833_Y), .B1(T4853_Y));
KC_AOI32_X1 T11908 ( .B0(T700_Y), .A0(T9373_Y), .A1(T862_Q),     .Y(T11908_Y), .A2(T1049_Y), .B1(T862_Q));
KC_AOI32_X1 T11907 ( .B0(T542_Y), .A0(T6691_Y), .A1(T5264_Q),     .Y(T11907_Y), .A2(T1034_Y), .B1(T5264_Q));
KC_AOI32_X1 T11087 ( .B0(T9262_Y), .A0(T829_Q), .A1(T12904_Y),     .Y(T11087_Y), .A2(T380_Y), .B1(T12904_Y));
KC_AOI32_X1 T11874 ( .B0(T542_Y), .A0(T6691_Y), .A1(T4858_Q),     .Y(T11874_Y), .A2(T7630_Y), .B1(T4858_Q));
KC_AOI32_X1 T11864 ( .B0(T886_Y), .A0(T11140_Y), .A1(T7357_Y),     .Y(T11864_Y), .A2(T7418_Y), .B1(T7357_Y));
KC_AOI32_X1 T11863 ( .B0(T6650_Y), .A0(T637_Y), .A1(T865_Q),     .Y(T11863_Y), .A2(T4863_Y), .B1(T865_Q));
KC_AOI32_X1 T11861 ( .B0(T15432_Y), .A0(T9374_Y), .A1(T863_Q),     .Y(T11861_Y), .A2(T1056_Y), .B1(T863_Q));
KC_AOI32_X1 T11157 ( .B0(T726_Y), .A0(T727_Y), .A1(T696_Q),     .Y(T11157_Y), .A2(T1053_Y), .B1(T696_Q));
KC_AOI32_X1 T11202 ( .B0(T726_Y), .A0(T727_Y), .A1(T5308_Q),     .Y(T11202_Y), .A2(T7630_Y), .B1(T5308_Q));
KC_AOI32_X1 T11195 ( .B0(T8727_Y), .A0(T5302_Y), .A1(T8714_Q),     .Y(T11195_Y), .A2(T8716_Y), .B1(T8714_Q));
KC_AOI32_X1 T11194 ( .B0(T700_Y), .A0(T9373_Y), .A1(T5301_Q),     .Y(T11194_Y), .A2(T7630_Y), .B1(T5301_Q));
KC_AOI32_X1 T11181 ( .B0(T744_Y), .A0(T10942_Y), .A1(T755_Y),     .Y(T11181_Y), .A2(T15454_Y), .B1(T755_Y));
KC_AOI32_X1 T11180 ( .B0(T8727_Y), .A0(T719_Y), .A1(T709_Q),     .Y(T11180_Y), .A2(T8716_Y), .B1(T709_Q));
KC_AOI32_X1 T11179 ( .B0(T8727_Y), .A0(T934_Y), .A1(T935_Q),     .Y(T11179_Y), .A2(T8716_Y), .B1(T935_Q));
KC_AOI32_X1 T11178 ( .B0(T15432_Y), .A0(T9374_Y), .A1(T5309_Q),     .Y(T11178_Y), .A2(T7630_Y), .B1(T5309_Q));
KC_AOI32_X1 T11244 ( .B0(T5353_Q), .A0(T15466_Y), .A1(T951_Y),     .Y(T11244_Y), .A2(T7843_Y), .B1(T7878_Y));
KC_AOI32_X1 T11217 ( .B0(T8770_Y), .A0(T11218_Y), .A1(T783_Y),     .Y(T11217_Y), .A2(T908_Y), .B1(T783_Y));
KC_AOI32_X1 T11275 ( .B0(T8093_Y), .A0(T8060_Y), .A1(T1395_Y),     .Y(T11275_Y), .A2(T1551_Y), .B1(T9000_Y));
KC_AOI32_X1 T11909 ( .B0(T577_Y), .A0(T497_Y), .A1(T6486_Q),     .Y(T11909_Y), .A2(T4857_Y), .B1(T6486_Q));
KC_AOI32_X1 T11877 ( .B0(T8727_Y), .A0(T15750_Y), .A1(T1041_Q),     .Y(T11877_Y), .A2(T8716_Y), .B1(T1041_Q));
KC_AOI32_X1 T11876 ( .B0(T8727_Y), .A0(T6651_Y), .A1(T1040_Q),     .Y(T11876_Y), .A2(T8716_Y), .B1(T1040_Q));
KC_AOI32_X1 T11875 ( .B0(T8727_Y), .A0(T6652_Y), .A1(T1046_Q),     .Y(T11875_Y), .A2(T8716_Y), .B1(T1046_Q));
KC_AOI32_X1 T11862 ( .B0(T546_Y), .A0(T549_Y), .A1(T6487_Q),     .Y(T11862_Y), .A2(T6796_Y), .B1(T6487_Q));
KC_AOI32_X1 T11171 ( .B0(T1044_Q), .A0(T5297_Q), .A1(T596_Y),     .Y(T11171_Y), .A2(T7741_Y), .B1(T596_Y));
KC_AOI32_X1 T11165 ( .B0(T546_Y), .A0(T549_Y), .A1(T1037_Q),     .Y(T11165_Y), .A2(T7630_Y), .B1(T1037_Q));
KC_AOI32_X1 T11155 ( .B0(T7411_Y), .A0(T8657_Y), .A1(T1045_Q),     .Y(T11155_Y), .A2(T6694_Y), .B1(T1045_Q));
KC_AOI32_X1 T11154 ( .B0(T11171_Y), .A0(T9714_Y), .A1(T1043_Y),     .Y(T11154_Y), .A2(T854_Y), .B1(T1043_Y));
KC_AOI32_X1 T11142 ( .B0(T577_Y), .A0(T497_Y), .A1(T1044_Q),     .Y(T11142_Y), .A2(T7630_Y), .B1(T1044_Q));
KC_AOI32_X1 T11193 ( .B0(T1066_Q), .A0(T5561_Q), .A1(T656_Y),     .Y(T11193_Y), .A2(T7638_Y), .B1(T656_Y));
KC_AOI32_X1 T11245 ( .B0(T1127_Q), .A0(T1100_Q), .A1(T16384_Y),     .Y(T11245_Y), .A2(T16422_Q), .B1(T8800_Y));
KC_AOI32_X1 T11305 ( .B0(T1366_Y), .A0(T4868_Y), .A1(T1362_Y),     .Y(T11305_Y), .A2(T15529_Y), .B1(T1362_Y));
KC_AOI32_X1 T11596 ( .B0(T11481_Y), .A0(T10207_Y), .A1(T11594_Y),     .Y(T11596_Y), .A2(T10224_Y), .B1(T11594_Y));
KC_AOI32_X1 T11552 ( .B0(T15974_Y), .A0(T1749_Y), .A1(T10946_Y),     .Y(T11552_Y), .A2(T5966_Y), .B1(T10946_Y));
KC_AOI32_X1 T11840 ( .B0(T291_Y), .A0(T6498_Y), .A1(T11838_Y),     .Y(T11840_Y), .A2(T11827_Y), .B1(T11838_Y));
KC_AOI32_X1 T11827 ( .B0(T6543_Y), .A0(T11772_Y), .A1(T6542_Y),     .Y(T11827_Y), .A2(T6541_Y), .B1(T6542_Y));
KC_AOI32_X1 T11258 ( .B0(T1999_Y), .A0(T868_Y), .A1(T2028_Q),     .Y(T11258_Y), .A2(T11949_Y), .B1(T2028_Q));
KC_AOI32_X1 T11257 ( .B0(T10524_Y), .A0(T1990_Y), .A1(T2016_Q),     .Y(T11257_Y), .A2(T11949_Y), .B1(T2016_Q));
KC_AOI32_X1 T11256 ( .B0(T1993_Y), .A0(T1118_Y), .A1(T2015_Q),     .Y(T11256_Y), .A2(T1992_Y), .B1(T16378_Y));
KC_AOI32_X1 T11255 ( .B0(T9951_Y), .A0(T5881_Y), .A1(T2005_Q),     .Y(T11255_Y), .A2(T1991_Y), .B1(T868_Y));
KC_AOI32_X1 T11994 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T15860_Q),     .Y(T11994_Y), .A2(T2127_Y), .B1(T15860_Q));
KC_AOI32_X1 T11993 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T2689_Q),     .Y(T11993_Y), .A2(T15853_Y), .B1(T2689_Q));
KC_AOI32_X1 T11992 ( .B0(T2707_Y), .A0(T11432_Y), .A1(T15798_Q),     .Y(T11992_Y), .A2(T5759_Y), .B1(T15798_Q));
KC_AOI32_X1 T11417 ( .B0(T2707_Y), .A0(T11432_Y), .A1(T15809_Q),     .Y(T11417_Y), .A2(T5834_Y), .B1(T15809_Q));
KC_AOI32_X1 T11416 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T2114_Q),     .Y(T11416_Y), .A2(T15881_Y), .B1(T2114_Q));
KC_AOI32_X1 T11415 ( .B0(T2707_Y), .A0(T11432_Y), .A1(T15797_Q),     .Y(T11415_Y), .A2(T5833_Y), .B1(T15797_Q));
KC_AOI32_X1 T11386 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T5574_Q),     .Y(T11386_Y), .A2(T15912_Y), .B1(T5574_Q));
KC_AOI32_X1 T11385 ( .B0(T2707_Y), .A0(T11432_Y), .A1(T5380_Q),     .Y(T11385_Y), .A2(T15701_Y), .B1(T5380_Q));
KC_AOI32_X1 T11384 ( .B0(T2707_Y), .A0(T11432_Y), .A1(T15844_Q),     .Y(T11384_Y), .A2(T15859_Y), .B1(T15844_Q));
KC_AOI32_X1 T11529 ( .B0(T13132_Q), .A0(T15005_Y), .A1(T5943_Y),     .Y(T11529_Y), .A2(T3411_Y), .B1(T8316_Y));
KC_AOI32_X1 T11585 ( .B0(T6015_Y), .A0(T5967_Y), .A1(T16070_Y),     .Y(T11585_Y), .A2(T5982_Y), .B1(T16070_Y));
KC_AOI32_X1 T11569 ( .B0(T6015_Y), .A0(T5967_Y), .A1(T16072_Y),     .Y(T11569_Y), .A2(T5878_Y), .B1(T16072_Y));
KC_AOI32_X1 T11568 ( .B0(T6015_Y), .A0(T5967_Y), .A1(T16075_Y),     .Y(T11568_Y), .A2(T15590_Y), .B1(T16075_Y));
KC_AOI32_X1 T11550 ( .B0(T6015_Y), .A0(T5967_Y), .A1(T16071_Y),     .Y(T11550_Y), .A2(T6004_Y), .B1(T16071_Y));
KC_AOI32_X1 T11549 ( .B0(T6015_Y), .A0(T5967_Y), .A1(T16074_Y),     .Y(T11549_Y), .A2(T5902_Y), .B1(T16074_Y));
KC_AOI32_X1 T11621 ( .B0(T2854_Y), .A0(T16016_Y), .A1(T2232_Y),     .Y(T11621_Y), .A2(T5007_Y), .B1(T2232_Y));
KC_AOI32_X1 T12063 ( .B0(T12105_Y), .A0(T12101_Y), .A1(T6101_Y),     .Y(T12063_Y), .A2(T6225_Y), .B1(T6101_Y));
KC_AOI32_X1 T11812 ( .B0(T6232_Y), .A0(T12063_Y), .A1(T12108_Y),     .Y(T11812_Y), .A2(T16130_Y), .B1(T12108_Y));
KC_AOI32_X1 T11749 ( .B0(T11775_Y), .A0(T5527_Q), .A1(T2328_Y),     .Y(T11749_Y), .A2(T6523_Y), .B1(T2328_Y));
KC_AOI32_X1 T11748 ( .B0(T2326_Y), .A0(T5529_Q), .A1(T12301_Y),     .Y(T11748_Y), .A2(T2364_Q), .B1(T12301_Y));
KC_AOI32_X1 T11839 ( .B0(T8173_Y), .A0(T2362_Y), .A1(T11034_Y),     .Y(T11839_Y), .A2(T2363_Y), .B1(T11034_Y));
KC_AOI32_X1 T11033 ( .B0(T6521_Y), .A0(T12321_Y), .A1(T2363_Y),     .Y(T11033_Y), .A2(T2362_Y), .B1(T12321_Y));
KC_AOI32_X1 T11948 ( .B0(T9748_Y), .A0(T610_Y), .A1(T2460_Y),     .Y(T11948_Y), .A2(T2454_Y), .B1(T2460_Y));
KC_AOI32_X1 T11947 ( .B0(T9745_Y), .A0(T610_Y), .A1(T611_Y),     .Y(T11947_Y), .A2(T2482_Y), .B1(T2478_Y));
KC_AOI32_X1 T11361 ( .B0(T11321_Y), .A0(T14527_Q), .A1(T2682_Y),     .Y(T11361_Y), .A2(T2698_Y), .B1(T2682_Y));
KC_AOI32_X1 T11360 ( .B0(T11362_Y), .A0(T14537_Q), .A1(T2682_Y),     .Y(T11360_Y), .A2(T2788_Y), .B1(T2682_Y));
KC_AOI32_X1 T11340 ( .B0(T6063_Y), .A0(T2693_Y), .A1(T5776_Y),     .Y(T11340_Y), .A2(T5775_Y), .B1(T5776_Y));
KC_AOI32_X1 T11339 ( .B0(T11343_Y), .A0(T14535_Q), .A1(T15830_Y),     .Y(T11339_Y), .A2(T14536_Q), .B1(T15830_Y));
KC_AOI32_X1 T11338 ( .B0(T11342_Y), .A0(T14533_Q), .A1(T2682_Y),     .Y(T11338_Y), .A2(T5786_Y), .B1(T2682_Y));
KC_AOI32_X1 T11429 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T15891_Q),     .Y(T11429_Y), .A2(T15858_Y), .B1(T15891_Q));
KC_AOI32_X1 T11396 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T15879_Q),     .Y(T11396_Y), .A2(T15857_Y), .B1(T15879_Q));
KC_AOI32_X1 T11383 ( .B0(T2707_Y), .A0(T11432_Y), .A1(T16088_Q),     .Y(T11383_Y), .A2(T5812_Y), .B1(T16088_Q));
KC_AOI32_X1 T11368 ( .B0(T2707_Y), .A0(T11432_Y), .A1(T15005_Y),     .Y(T11368_Y), .A2(T2708_Y), .B1(T15005_Y));
KC_AOI32_X1 T11462 ( .B0(T13123_Y), .A0(T3411_Y), .A1(T13112_Q),     .Y(T11462_Y), .A2(T5896_Y), .B1(T13112_Q));
KC_AOI32_X1 T11461 ( .B0(T13123_Y), .A0(T3411_Y), .A1(T13111_Q),     .Y(T11461_Y), .A2(T11025_Y), .B1(T13111_Q));
KC_AOI32_X1 T11598 ( .B0(T16100_Y), .A0(T6007_Y), .A1(T2723_Y),     .Y(T11598_Y), .A2(T5944_Y), .B1(T6011_Y));
KC_AOI32_X1 T11678 ( .B0(T6088_Y), .A0(T16167_Y), .A1(T6085_Y),     .Y(T11678_Y), .A2(T3369_Y), .B1(T3379_Y));
KC_AOI32_X1 T11665 ( .B0(T11831_Y), .A0(T16102_Y), .A1(T6070_Y),     .Y(T11665_Y), .A2(T11647_Y), .B1(T6070_Y));
KC_AOI32_X1 T11649 ( .B0(T6054_Y), .A0(T2829_Y), .A1(T3398_Y),     .Y(T11649_Y), .A2(T15943_Y), .B1(T3398_Y));
KC_AOI32_X1 T11704 ( .B0(T11809_Y), .A0(T2906_Y), .A1(T12048_Y),     .Y(T11704_Y), .A2(T4748_Y), .B1(T12048_Y));
KC_AOI32_X1 T11699 ( .B0(T6145_Y), .A0(T6583_Y), .A1(T15622_Y),     .Y(T11699_Y), .A2(T6180_Y), .B1(T15622_Y));
KC_AOI32_X1 T12062 ( .B0(T4998_Y), .A0(T8261_Y), .A1(T11742_Y),     .Y(T12062_Y), .A2(T6573_Y), .B1(T11742_Y));
KC_AOI32_X1 T11807 ( .B0(T15255_Y), .A0(T2359_Q), .A1(T6214_Y),     .Y(T11807_Y), .A2(T6556_Y), .B1(T6214_Y));
KC_AOI32_X1 T11806 ( .B0(T12107_Y), .A0(T12102_Y), .A1(T10573_Y),     .Y(T11806_Y), .A2(T16131_Y), .B1(T6571_Y));
KC_AOI32_X1 T11768 ( .B0(T8409_Y), .A0(T6560_Y), .A1(T6225_Y),     .Y(T11768_Y), .A2(T12867_Y), .B1(T6225_Y));
KC_AOI32_X1 T11821 ( .B0(T12067_Y), .A0(T15643_Y), .A1(T12862_Y),     .Y(T11821_Y), .A2(T3436_Y), .B1(T12862_Y));
KC_AOI32_X1 T11309 ( .B0(T10268_Y), .A0(T14950_Q), .A1(T10241_Y),     .Y(T11309_Y), .A2(T5077_Y), .B1(T10241_Y));
KC_AOI32_X1 T11395 ( .B0(T3855_Y), .A0(T15010_Y), .A1(T10898_Y),     .Y(T11395_Y), .A2(T3224_Y), .B1(T10898_Y));
KC_AOI32_X1 T11382 ( .B0(T3855_Y), .A0(T3223_Y), .A1(T10898_Y),     .Y(T11382_Y), .A2(T5039_Y), .B1(T10898_Y));
KC_AOI32_X1 T11486 ( .B0(T3303_Y), .A0(T5894_Y), .A1(T8267_Y),     .Y(T11486_Y), .A2(T6231_Co), .B1(T6231_S));
KC_AOI32_X1 T11591 ( .B0(T15977_Y), .A0(T2719_Y), .A1(T3318_Y),     .Y(T11591_Y), .A2(T15978_Y), .B1(T15976_Y));
KC_AOI32_X1 T11610 ( .B0(T6320_S), .A0(T11609_Y), .A1(T4468_Y),     .Y(T11610_Y), .A2(T12240_Y), .B1(T15133_Y));
KC_AOI32_X1 T11609 ( .B0(T16015_Y), .A0(T6335_Y), .A1(T7915_Y),     .Y(T11609_Y), .A2(T16015_Y), .B1(T6024_Y));
KC_AOI32_X1 T11999 ( .B0(T3357_Y), .A0(T6036_Y), .A1(T10965_Y),     .Y(T11999_Y), .A2(T15613_Y), .B1(T10965_Y));
KC_AOI32_X1 T11998 ( .B0(T8228_Y), .A0(T12263_Y), .A1(T12043_Y),     .Y(T11998_Y), .A2(T16302_Y), .B1(T12043_Y));
KC_AOI32_X1 T11640 ( .B0(T12249_Y), .A0(T11664_Y), .A1(T16102_Y),     .Y(T11640_Y), .A2(T6052_Y), .B1(T16102_Y));
KC_AOI32_X1 T11723 ( .B0(T12322_Y), .A0(T3408_Y), .A1(T2919_Y),     .Y(T11723_Y), .A2(T5054_Y), .B1(T2919_Y));
KC_AOI32_X1 T11722 ( .B0(T11739_Y), .A0(T12044_Y), .A1(T11831_Y),     .Y(T11722_Y), .A2(T3418_Y), .B1(T11831_Y));
KC_AOI32_X1 T11703 ( .B0(T6147_Y), .A0(T15711_Y), .A1(T15233_Y),     .Y(T11703_Y), .A2(T8342_Y), .B1(T15233_Y));
KC_AOI32_X1 T11695 ( .B0(T15233_Y), .A0(T3426_Y), .A1(T6147_Y),     .Y(T11695_Y), .A2(T3424_Y), .B1(T6147_Y));
KC_AOI32_X1 T11684 ( .B0(T3442_Y), .A0(T6096_Y), .A1(T12317_Y),     .Y(T11684_Y), .A2(T10583_Y), .B1(T12317_Y));
KC_AOI32_X1 T12059 ( .B0(T3427_Y), .A0(T6575_Y), .A1(T12969_Y),     .Y(T12059_Y), .A2(T12283_Y), .B1(T12969_Y));
KC_AOI32_X1 T11800 ( .B0(T11796_Y), .A0(T11802_Y), .A1(T6549_Q),     .Y(T11800_Y), .A2(T5048_Y), .B1(T5072_Y));
KC_AOI32_X1 T11738 ( .B0(T15641_Y), .A0(T5047_Y), .A1(T5521_Y),     .Y(T11738_Y), .A2(T6215_Y), .B1(T5521_Y));
KC_AOI32_X1 T11980 ( .B0(T11983_Y), .A0(T11378_Y), .A1(T16154_Y),     .Y(T11980_Y), .A2(T15907_Y), .B1(T16154_Y));
KC_AOI32_X1 T11351 ( .B0(T11983_Y), .A0(T11365_Y), .A1(T11379_Y),     .Y(T11351_Y), .A2(T5802_Y), .B1(T11379_Y));
KC_AOI32_X1 T11334 ( .B0(T5788_Y), .A0(T3797_Y), .A1(T4465_Q),     .Y(T11334_Y), .A2(T3806_Y), .B1(T3809_Y));
KC_AOI32_X1 T11333 ( .B0(T4465_Q), .A0(T12137_Y), .A1(T5779_Y),     .Y(T11333_Y), .A2(T4420_Y), .B1(T5779_Y));
KC_AOI32_X1 T11331 ( .B0(T15821_Y), .A0(T11351_Y), .A1(T16160_Y),     .Y(T11331_Y), .A2(T12138_Y), .B1(T5774_Y));
KC_AOI32_X1 T11316 ( .B0(T11969_Y), .A0(T5816_Y), .A1(T3802_Y),     .Y(T11316_Y), .A2(T3788_Y), .B1(T3802_Y));
KC_AOI32_X1 T11425 ( .B0(T14494_Q), .A0(T16153_Y), .A1(T3856_Y),     .Y(T11425_Y), .A2(T14495_Q), .B1(T3856_Y));
KC_AOI32_X1 T11407 ( .B0(T5788_Y), .A0(T5842_Y), .A1(T11404_Y),     .Y(T11407_Y), .A2(T10911_Y), .B1(T11404_Y));
KC_AOI32_X1 T11406 ( .B0(T16153_Y), .A0(T3854_Y), .A1(T5815_Y),     .Y(T11406_Y), .A2(T15907_Y), .B1(T144_Q));
KC_AOI32_X1 T11405 ( .B0(T11379_Y), .A0(T11408_Y), .A1(T144_Q),     .Y(T11405_Y), .A2(T5788_Y), .B1(T144_Q));
KC_AOI32_X1 T11404 ( .B0(T11394_Y), .A0(T11381_Y), .A1(T15908_Y),     .Y(T11404_Y), .A2(T5823_Y), .B1(T15908_Y));
KC_AOI32_X1 T11392 ( .B0(T11375_Y), .A0(T15897_Y), .A1(T11428_Y),     .Y(T11392_Y), .A2(T5802_Y), .B1(T11428_Y));
KC_AOI32_X1 T11391 ( .B0(T5803_Y), .A0(T4486_Y), .A1(T8196_Y),     .Y(T11391_Y), .A2(T11406_Y), .B1(T8196_Y));
KC_AOI32_X1 T11390 ( .B0(T11392_Y), .A0(T11378_Y), .A1(T4465_Q),     .Y(T11390_Y), .A2(T3826_Y), .B1(T4465_Q));
KC_AOI32_X1 T11967 ( .B0(T4466_Y), .A0(T15897_Y), .A1(T15907_Y),     .Y(T11967_Y), .A2(T5852_Y), .B1(T15907_Y));
KC_AOI32_X1 T11514 ( .B0(T5981_Y), .A0(T8352_Q), .A1(T10937_Y),     .Y(T11514_Y), .A2(T3966_Y), .B1(T3968_Q));
KC_AOI32_X1 T11513 ( .B0(T11587_Y), .A0(T6204_Y), .A1(T12227_Y),     .Y(T11513_Y), .A2(T5989_Y), .B1(T12227_Y));
KC_AOI32_X1 T11512 ( .B0(T5919_Y), .A0(T11023_Y), .A1(T3907_Y),     .Y(T11512_Y), .A2(T10935_Y), .B1(T3907_Y));
KC_AOI32_X1 T11511 ( .B0(T5981_Y), .A0(T15138_Q), .A1(T10937_Y),     .Y(T11511_Y), .A2(T3966_Y), .B1(T3965_Q));
KC_AOI32_X1 T11635 ( .B0(T3530_Y), .A0(T13130_Q), .A1(T6060_Y),     .Y(T11635_Y), .A2(T15601_Y), .B1(T6060_Y));
KC_AOI32_X1 T11625 ( .B0(T4179_Q), .A0(T15760_Q), .A1(T4176_Q),     .Y(T11625_Y), .A2(T4035_Y), .B1(T4176_Q));
KC_AOI32_X1 T11708 ( .B0(T5568_Q), .A0(T11713_Y), .A1(T5135_Y),     .Y(T11708_Y), .A2(T6137_Y), .B1(T15619_Y));
KC_AOI32_X1 T11693 ( .B0(T5056_Y), .A0(T11657_Y), .A1(T4113_Y),     .Y(T11693_Y), .A2(T6046_Y), .B1(T4113_Y));
KC_AOI32_X1 T11794 ( .B0(T10983_Y), .A0(T6526_Q), .A1(T6547_Y),     .Y(T11794_Y), .A2(T3469_Y), .B1(T6547_Y));
KC_AOI32_X1 T11793 ( .B0(T10994_Y), .A0(T5525_Q), .A1(T6547_Y),     .Y(T11793_Y), .A2(T3469_Y), .B1(T6547_Y));
KC_AOI32_X1 T11762 ( .B0(T10982_Y), .A0(T6555_Q), .A1(T6547_Y),     .Y(T11762_Y), .A2(T3469_Y), .B1(T6547_Y));
KC_AOI32_X1 T11761 ( .B0(T11795_Y), .A0(T16102_Y), .A1(T4169_Q),     .Y(T11761_Y), .A2(T16142_Y), .B1(T4169_Q));
KC_AOI32_X1 T11829 ( .B0(T11813_Y), .A0(T4163_Q), .A1(T11817_Y),     .Y(T11829_Y), .A2(T4119_Y), .B1(T11817_Y));
KC_AOI32_X1 T11346 ( .B0(T4487_Q), .A0(T145_Q), .A1(T5789_Y),     .Y(T11346_Y), .A2(T5760_Y), .B1(T4389_Y));
KC_AOI32_X1 T11345 ( .B0(T15872_Y), .A0(T11976_Y), .A1(T12143_Y),     .Y(T11345_Y), .A2(T14523_Q), .B1(T12143_Y));
KC_AOI32_X1 T11419 ( .B0(T5823_Y), .A0(T16154_Y), .A1(T5789_Y),     .Y(T11419_Y), .A2(T5835_Y), .B1(T4487_Q));
KC_AOI32_X1 T11400 ( .B0(T4448_Y), .A0(T5789_Y), .A1(T5800_Y),     .Y(T11400_Y), .A2(T4478_Y), .B1(T5800_Y));
KC_AOI32_X1 T11369 ( .B0(T11421_Y), .A0(T11365_Y), .A1(T3856_Y),     .Y(T11369_Y), .A2(T3826_Y), .B1(T3856_Y));
KC_AOI32_X1 T11364 ( .B0(T3838_Y), .A0(T4487_Q), .A1(T3850_Y),     .Y(T11364_Y), .A2(T8442_Y), .B1(T3850_Y));
KC_AOI32_X1 T11966 ( .B0(T11422_Y), .A0(T11365_Y), .A1(T14549_Q),     .Y(T11966_Y), .A2(T15871_Y), .B1(T5854_Y));
KC_AOI32_X1 T11441 ( .B0(T8444_Y), .A0(T10922_Y), .A1(T5107_Y),     .Y(T11441_Y), .A2(T4499_Y), .B1(T5107_Y));
KC_AOI32_X1 T11440 ( .B0(T11442_Y), .A0(T14548_Q), .A1(T5851_Y),     .Y(T11440_Y), .A2(T14550_Q), .B1(T5851_Y));
KC_AOI32_X1 T11518 ( .B0(T12209_Y), .A0(T5884_Y), .A1(T4524_Y),     .Y(T11518_Y), .A2(T5934_Y), .B1(T11521_Y));
KC_AOI32_X1 T11504 ( .B0(T5459_Y), .A0(T4514_Y), .A1(T2073_Y),     .Y(T11504_Y), .A2(T15969_Y), .B1(T2073_Y));
KC_AOI32_X1 T11503 ( .B0(T15706_Y), .A0(T4528_Q), .A1(T5140_Y),     .Y(T11503_Y), .A2(T11507_Y), .B1(T5140_Y));
KC_AOI32_X1 T11606 ( .B0(T4612_Y), .A0(T9486_Y), .A1(T3973_Y),     .Y(T11606_Y), .A2(T4616_Y), .B1(T8312_Y));
KC_AOI32_X1 T6056 ( .B0(T16111_Y), .A0(T8355_Y), .A1(T4650_Y),     .Y(T6056_Y), .A2(T6057_Y), .B1(T4650_Y));
KC_AOI32_X1 T11670 ( .B0(T6076_Y), .A0(T8368_Y), .A1(T4651_Y),     .Y(T11670_Y), .A2(T6057_Y), .B1(T4651_Y));
KC_AOI32_X1 T11655 ( .B0(T6075_Y), .A0(T8369_Y), .A1(T4649_Y),     .Y(T11655_Y), .A2(T6057_Y), .B1(T4649_Y));
KC_AOI32_X1 T11681 ( .B0(T6091_Y), .A0(T4736_Y), .A1(T4707_Y),     .Y(T11681_Y), .A2(T15141_Y), .B1(T4707_Y));
KC_AOI32_X1 T11680 ( .B0(T4736_Y), .A0(T16460_Q), .A1(T15141_Y),     .Y(T11680_Y), .A2(T12033_Y), .B1(T15141_Y));
KC_AOI32_X1 T12053 ( .B0(T4739_Y), .A0(T16460_Q), .A1(T15634_Y),     .Y(T12053_Y), .A2(T10599_Y), .B1(T15634_Y));
KC_AOI32_X1 T11785 ( .B0(T5339_Y), .A0(T4739_Y), .A1(T4730_Y),     .Y(T11785_Y), .A2(T15634_Y), .B1(T4730_Y));
KC_AOI32_X1 T11759 ( .B0(T6203_Y), .A0(T4736_Y), .A1(T4752_Y),     .Y(T11759_Y), .A2(T12308_Y), .B1(T4752_Y));
KC_AOI32_X1 T11898 ( .B0(T9083_Y), .A0(T16286_Y), .A1(T1603_Y),     .Y(T11898_Y), .A2(T9453_Y), .B1(T9454_Y));
KC_AOI32_X1 T11893 ( .B0(T7673_Y), .A0(T9379_Y), .A1(T8778_Y),     .Y(T11893_Y), .A2(T9388_Y), .B1(T8778_Y));
KC_AOI32_X1 T11878 ( .B0(T6650_Y), .A0(T637_Y), .A1(T1066_Q),     .Y(T11878_Y), .A2(T7630_Y), .B1(T1066_Q));
KC_AOI32_X1 T11918 ( .B0(T1037_Q), .A0(T1084_Q), .A1(T15751_Y),     .Y(T11918_Y), .A2(T7719_Y), .B1(T15751_Y));
KC_AOI32_X1 T11880 ( .B0(T4858_Q), .A0(T5310_Q), .A1(T15665_Y),     .Y(T11880_Y), .A2(T7719_Y), .B1(T15665_Y));
KC_AOI32_X1 T11879 ( .B0(T8727_Y), .A0(T658_Y), .A1(T1068_Q),     .Y(T11879_Y), .A2(T8716_Y), .B1(T1068_Q));
KC_AOI32_X1 T11860 ( .B0(T7411_Y), .A0(T8716_Y), .A1(T5262_Q),     .Y(T11860_Y), .A2(T9723_Y), .B1(T5262_Q));
KC_AOI32_X1 T11914 ( .B0(T12109_Y), .A0(T10299_Y), .A1(T16276_Y),     .Y(T11914_Y), .A2(T16275_Y), .B1(T16276_Y));
KC_AOI32_X1 T12006 ( .B0(T8345_Y), .A0(T10584_Y), .A1(T15804_Q),     .Y(T12006_Y), .A2(T16036_Y), .B1(T15804_Q));
KC_AOI32_X1 T12005 ( .B0(T6006_Y), .A0(T5556_Y), .A1(T2805_Y),     .Y(T12005_Y), .A2(T11019_Y), .B1(T2805_Y));
KC_AOI32_X1 T12058 ( .B0(T3427_Y), .A0(T15257_Y), .A1(T12970_Y),     .Y(T12058_Y), .A2(T5507_Y), .B1(T12970_Y));
KC_AOI32_X1 T11986 ( .B0(T15864_Y), .A0(T5102_Y), .A1(T16160_Y),     .Y(T11986_Y), .A2(T11390_Y), .B1(T5774_Y));
KC_AOI32_X1 T11958 ( .B0(T5748_Y), .A0(T5077_Y), .A1(T5747_Y),     .Y(T11958_Y), .A2(T3211_Y), .B1(T5747_Y));
KC_AOI32_X1 T11036 ( .B0(T12069_Y), .A0(T12069_Y), .A1(T12070_Y),     .Y(T11036_Y), .A2(T6545_Y), .B1(T12070_Y));
KC_AOI32_X1 T12055 ( .B0(T11790_Y), .A0(T16102_Y), .A1(T6547_Y),     .Y(T12055_Y), .A2(T11693_Y), .B1(T6547_Y));
KC_AOI32_X1 T12037 ( .B0(T4058_Y), .A0(T16106_Y), .A1(T4065_Y),     .Y(T12037_Y), .A2(T4046_Y), .B1(T4065_Y));
KC_AOI32_X1 T12025 ( .B0(T11587_Y), .A0(T5905_Y), .A1(T12026_Y),     .Y(T12025_Y), .A2(T5989_Y), .B1(T12026_Y));
KC_AOI32_X1 T11974 ( .B0(T145_Q), .A0(T4404_Y), .A1(T4486_Y),     .Y(T11974_Y), .A2(T4452_Y), .B1(T8450_Y));
KC_AOI32_X1 T11332 ( .B0(T5764_Y), .A0(T11334_Y), .A1(T16160_Y),     .Y(T11332_Y), .A2(T3796_Y), .B1(T5774_Y));
KC_AOI32_X1 T11329 ( .B0(T11982_Y), .A0(T11365_Y), .A1(T11428_Y),     .Y(T11329_Y), .A2(T4394_Y), .B1(T11428_Y));
KC_AOI32_X1 T15041 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T15880_Q),     .Y(T15041_Y), .A2(T10245_Y), .B1(T15880_Q));
KC_AOI32_X1 T11430 ( .B0(T12340_Y), .A0(T11432_Y), .A1(T15894_Q),     .Y(T11430_Y), .A2(T16474_Y), .B1(T15894_Q));
KC_AOI32_X1 T11420 ( .B0(T3827_Y), .A0(T6114_Y), .A1(T12150_Y),     .Y(T11420_Y), .A2(T5446_Y), .B1(T12150_Y));
KC_AOI32_X1 T11611 ( .B0(T2854_Y), .A0(T12231_Y), .A1(T2282_Y),     .Y(T11611_Y), .A2(T2799_Y), .B1(T2282_Y));
KC_AOI32_X1 T11629 ( .B0(T3399_Y), .A0(T10961_Y), .A1(T8503_Y),     .Y(T11629_Y), .A2(T12830_Y), .B1(T8503_Y));
KC_AOI32_X1 T11971 ( .B0(T6737_Y), .A0(T5444_Y), .A1(T4931_Y),     .Y(T11971_Y), .A2(T15906_Y), .B1(T5793_Y));
KC_OAI112_X1 T12367 ( .A(T5602_Y), .B(T116_Y), .C0(T8554_Y),     .C1(T5631_Y), .Y(T12367_Y));
KC_OAI112_X1 T11274 ( .A(T15490_Y), .B(T8989_Y), .C0(T1367_Y),     .C1(T1367_Y), .Y(T11274_Y));
KC_OAI112_X1 T11295 ( .A(T4817_Y), .B(T4804_Y), .C0(T9135_Y),     .C1(T4818_Y), .Y(T11295_Y));
KC_OAI112_X1 T11048 ( .A(T6859_Y), .B(T12373_Y), .C0(T433_Y),     .C1(T12373_Y), .Y(T11048_Y));
KC_OAI112_X1 T12387 ( .A(T6966_Y), .B(T6315_Y), .C0(T6819_Y),     .C1(T10906_Y), .Y(T12387_Y));
KC_OAI112_X1 T11071 ( .A(T6930_Y), .B(T6962_Y), .C0(T15740_Y),     .C1(T10906_Y), .Y(T11071_Y));
KC_OAI112_X1 T11070 ( .A(T6941_Y), .B(T295_Y), .C0(T9316_Y),     .C1(T10906_Y), .Y(T11070_Y));
KC_OAI112_X1 T11062 ( .A(T268_Y), .B(T6963_Y), .C0(T15740_Y),     .C1(T10916_Y), .Y(T11062_Y));
KC_OAI112_X1 T11058 ( .A(T6314_Y), .B(T6928_Y), .C0(T896_Y),     .C1(T10906_Y), .Y(T11058_Y));
KC_OAI112_X1 T11086 ( .A(T269_Y), .B(T7059_Y), .C0(T6835_Y),     .C1(T10916_Y), .Y(T11086_Y));
KC_OAI112_X1 T11084 ( .A(T7258_Y), .B(T7098_Y), .C0(T6819_Y),     .C1(T11010_Y), .Y(T11084_Y));
KC_OAI112_X1 T11083 ( .A(T7107_Y), .B(T6473_Y), .C0(T124_Q),     .C1(T10916_Y), .Y(T11083_Y));
KC_OAI112_X1 T11082 ( .A(T7106_Y), .B(T7086_Y), .C0(T9317_Y),     .C1(T10916_Y), .Y(T11082_Y));
KC_OAI112_X1 T11081 ( .A(T7103_Y), .B(T7099_Y), .C0(T124_Q),     .C1(T10906_Y), .Y(T11081_Y));
KC_OAI112_X1 T11075 ( .A(T6316_Y), .B(T6268_Y), .C0(T896_Y),     .C1(T10916_Y), .Y(T11075_Y));
KC_OAI112_X1 T11074 ( .A(T7072_Y), .B(T7070_Y), .C0(T6819_Y),     .C1(T10916_Y), .Y(T11074_Y));
KC_OAI112_X1 T11912 ( .A(T6814_Y), .B(T6600_Y), .C0(T6819_Y),     .C1(T15032_Y), .Y(T11912_Y));
KC_OAI112_X1 T11911 ( .A(T6813_Y), .B(T6599_Y), .C0(T9317_Y),     .C1(T15032_Y), .Y(T11911_Y));
KC_OAI112_X1 T11108 ( .A(T7317_Y), .B(T7312_Y), .C0(T896_Y),     .C1(T11011_Y), .Y(T11108_Y));
KC_OAI112_X1 T11107 ( .A(T7311_Y), .B(T7309_Y), .C0(T15740_Y),     .C1(T11010_Y), .Y(T11107_Y));
KC_OAI112_X1 T11100 ( .A(T7314_Y), .B(T325_Y), .C0(T9317_Y),     .C1(T11011_Y), .Y(T11100_Y));
KC_OAI112_X1 T11099 ( .A(T7316_Y), .B(T7313_Y), .C0(T6819_Y),     .C1(T11011_Y), .Y(T11099_Y));
KC_OAI112_X1 T11098 ( .A(T7310_Y), .B(T328_Y), .C0(T15740_Y),     .C1(T11011_Y), .Y(T11098_Y));
KC_OAI112_X1 T11097 ( .A(T7315_Y), .B(T7274_Y), .C0(T124_Q),     .C1(T11011_Y), .Y(T11097_Y));
KC_OAI112_X1 T11089 ( .A(T7256_Y), .B(T6475_Y), .C0(T896_Y),     .C1(T11010_Y), .Y(T11089_Y));
KC_OAI112_X1 T11088 ( .A(T7253_Y), .B(T6474_Y), .C0(T124_Q),     .C1(T11010_Y), .Y(T11088_Y));
KC_OAI112_X1 T11883 ( .A(T7457_Y), .B(T7456_Y), .C0(T6819_Y),     .C1(T14990_Y), .Y(T11883_Y));
KC_OAI112_X1 T11871 ( .A(T7403_Y), .B(T6719_Y), .C0(T9317_Y),     .C1(T14989_Y), .Y(T11871_Y));
KC_OAI112_X1 T11169 ( .A(T7458_Y), .B(T7453_Y), .C0(T15740_Y),     .C1(T14987_Y), .Y(T11169_Y));
KC_OAI112_X1 T11168 ( .A(T7383_Y), .B(T6674_Y), .C0(T124_Q),     .C1(T14987_Y), .Y(T11168_Y));
KC_OAI112_X1 T11161 ( .A(T7426_Y), .B(T346_Y), .C0(T15740_Y),     .C1(T14989_Y), .Y(T11161_Y));
KC_OAI112_X1 T11160 ( .A(T7428_Y), .B(T7423_Y), .C0(T124_Q),     .C1(T14989_Y), .Y(T11160_Y));
KC_OAI112_X1 T11159 ( .A(T7427_Y), .B(T7399_Y), .C0(T6819_Y),     .C1(T14989_Y), .Y(T11159_Y));
KC_OAI112_X1 T11153 ( .A(T7404_Y), .B(T7402_Y), .C0(T896_Y),     .C1(T14989_Y), .Y(T11153_Y));
KC_OAI112_X1 T11151 ( .A(T7381_Y), .B(T7430_Y), .C0(T896_Y),     .C1(T14990_Y), .Y(T11151_Y));
KC_OAI112_X1 T11149 ( .A(T7384_Y), .B(T336_Y), .C0(T9317_Y),     .C1(T14990_Y), .Y(T11149_Y));
KC_OAI112_X1 T11148 ( .A(T7389_Y), .B(T7432_Y), .C0(T9317_Y),     .C1(T14987_Y), .Y(T11148_Y));
KC_OAI112_X1 T11147 ( .A(T7382_Y), .B(T7454_Y), .C0(T6819_Y),     .C1(T14987_Y), .Y(T11147_Y));
KC_OAI112_X1 T11214 ( .A(T7693_Y), .B(T16324_Y), .C0(T7826_Y),     .C1(T7672_Y), .Y(T11214_Y));
KC_OAI112_X1 T11213 ( .A(T7689_Y), .B(T9376_Y), .C0(T7574_Y),     .C1(T9380_Y), .Y(T11213_Y));
KC_OAI112_X1 T11207 ( .A(T8699_Y), .B(T7577_Y), .C0(T7674_Y),     .C1(T16330_Y), .Y(T11207_Y));
KC_OAI112_X1 T11206 ( .A(T7573_Y), .B(T7568_Y), .C0(T7669_Y),     .C1(T16330_Y), .Y(T11206_Y));
KC_OAI112_X1 T11205 ( .A(T7666_Y), .B(T8743_Y), .C0(T740_Y),     .C1(T11206_Y), .Y(T11205_Y));
KC_OAI112_X1 T11188 ( .A(T15764_Y), .B(T8700_Y), .C0(T7575_Y),     .C1(T9383_Y), .Y(T11188_Y));
KC_OAI112_X1 T11187 ( .A(T15771_Y), .B(T8702_Y), .C0(T7673_Y),     .C1(T9383_Y), .Y(T11187_Y));
KC_OAI112_X1 T11186 ( .A(T7572_Y), .B(T8701_Y), .C0(T7567_Y),     .C1(T9380_Y), .Y(T11186_Y));
KC_OAI112_X1 T11185 ( .A(T7571_Y), .B(T9377_Y), .C0(T12607_Y),     .C1(T9383_Y), .Y(T11185_Y));
KC_OAI112_X1 T11184 ( .A(T12606_Y), .B(T7679_Y), .C0(T7672_Y),     .C1(T16330_Y), .Y(T11184_Y));
KC_OAI112_X1 T11897 ( .A(T16360_Y), .B(T8870_Y), .C0(T16390_Y),     .C1(T9423_Y), .Y(T11897_Y));
KC_OAI112_X1 T11896 ( .A(T8048_Y), .B(T8914_Y), .C0(T12886_Y),     .C1(T9425_Y), .Y(T11896_Y));
KC_OAI112_X1 T11895 ( .A(T8050_Y), .B(T8912_Y), .C0(T7906_Y),     .C1(T9423_Y), .Y(T11895_Y));
KC_OAI112_X1 T11247 ( .A(T16389_Y), .B(T9422_Y), .C0(T7908_Y),     .C1(T9425_Y), .Y(T11247_Y));
KC_OAI112_X1 T11246 ( .A(T15791_Y), .B(T8911_Y), .C0(T7856_Y),     .C1(T9425_Y), .Y(T11246_Y));
KC_OAI112_X1 T11234 ( .A(T7907_Y), .B(T8815_Y), .C0(T936_Y),     .C1(T11265_Y), .Y(T11234_Y));
KC_OAI112_X1 T11270 ( .A(T8075_Y), .B(T1329_Y), .C0(T8079_Y),     .C1(T7903_Y), .Y(T11270_Y));
KC_OAI112_X1 T11269 ( .A(T12722_Y), .B(T8083_Y), .C0(T7903_Y),     .C1(T8076_Y), .Y(T11269_Y));
KC_OAI112_X1 T11265 ( .A(T8049_Y), .B(T8052_Y), .C0(T7910_Y),     .C1(T8076_Y), .Y(T11265_Y));
KC_OAI112_X1 T11264 ( .A(T8913_Y), .B(T8053_Y), .C0(T7904_Y),     .C1(T8076_Y), .Y(T11264_Y));
KC_OAI112_X1 T11858 ( .A(T6260_Y), .B(T6310_Y), .C0(T6835_Y),     .C1(T11016_Y), .Y(T11858_Y));
KC_OAI112_X1 T11069 ( .A(T6957_Y), .B(T6955_Y), .C0(T6819_Y),     .C1(T10884_Y), .Y(T11069_Y));
KC_OAI112_X1 T11068 ( .A(T6906_Y), .B(T6903_Y), .C0(T9316_Y),     .C1(T10884_Y), .Y(T11068_Y));
KC_OAI112_X1 T11067 ( .A(T6960_Y), .B(T6953_Y), .C0(T15740_Y),     .C1(T10884_Y), .Y(T11067_Y));
KC_OAI112_X1 T11061 ( .A(T6926_Y), .B(T6924_Y), .C0(T896_Y),     .C1(T10884_Y), .Y(T11061_Y));
KC_OAI112_X1 T11060 ( .A(T6958_Y), .B(T6940_Y), .C0(T6819_Y),     .C1(T11016_Y), .Y(T11060_Y));
KC_OAI112_X1 T11057 ( .A(T6927_Y), .B(T6920_Y), .C0(T896_Y),     .C1(T11016_Y), .Y(T11057_Y));
KC_OAI112_X1 T11054 ( .A(T6959_Y), .B(T6956_Y), .C0(T15740_Y),     .C1(T11016_Y), .Y(T11054_Y));
KC_OAI112_X1 T11053 ( .A(T6905_Y), .B(T454_Y), .C0(T9318_Y),     .C1(T10884_Y), .Y(T11053_Y));
KC_OAI112_X1 T11052 ( .A(T6907_Y), .B(T6902_Y), .C0(T9316_Y),     .C1(T11016_Y), .Y(T11052_Y));
KC_OAI112_X1 T11051 ( .A(T6908_Y), .B(T219_Y), .C0(T9318_Y),     .C1(T11016_Y), .Y(T11051_Y));
KC_OAI112_X1 T11080 ( .A(T7095_Y), .B(T7113_Y), .C0(T124_Q),     .C1(T10884_Y), .Y(T11080_Y));
KC_OAI112_X1 T11079 ( .A(T7102_Y), .B(T6338_Y), .C0(T10906_Y),     .C1(T6803_Y), .Y(T11079_Y));
KC_OAI112_X1 T11910 ( .A(T6732_Y), .B(T6641_Y), .C0(T11011_Y),     .C1(T6803_Y), .Y(T11910_Y));
KC_OAI112_X1 T11106 ( .A(T7305_Y), .B(T7302_Y), .C0(T9319_Y),     .C1(T11010_Y), .Y(T11106_Y));
KC_OAI112_X1 T11105 ( .A(T7248_Y), .B(T7246_Y), .C0(T10916_Y),     .C1(T6803_Y), .Y(T11105_Y));
KC_OAI112_X1 T11096 ( .A(T7286_Y), .B(T7266_Y), .C0(T6835_Y),     .C1(T11011_Y), .Y(T11096_Y));
KC_OAI112_X1 T11095 ( .A(T7282_Y), .B(T7284_Y), .C0(T6835_Y),     .C1(T11010_Y), .Y(T11095_Y));
KC_OAI112_X1 T11094 ( .A(T7287_Y), .B(T7303_Y), .C0(T11010_Y),     .C1(T6803_Y), .Y(T11094_Y));
KC_OAI112_X1 T11090 ( .A(T7267_Y), .B(T7264_Y), .C0(T9319_Y),     .C1(T11011_Y), .Y(T11090_Y));
KC_OAI112_X1 T11866 ( .A(T6807_Y), .B(T6709_Y), .C0(T6835_Y),     .C1(T15032_Y), .Y(T11866_Y));
KC_OAI112_X1 T11167 ( .A(T7444_Y), .B(T7448_Y), .C0(T9319_Y),     .C1(T14990_Y), .Y(T11167_Y));
KC_OAI112_X1 T11158 ( .A(T7375_Y), .B(T7369_Y), .C0(T9319_Y),     .C1(T14989_Y), .Y(T11158_Y));
KC_OAI112_X1 T11146 ( .A(T7450_Y), .B(T7372_Y), .C0(T9319_Y),     .C1(T14987_Y), .Y(T11146_Y));
KC_OAI112_X1 T11145 ( .A(T7449_Y), .B(T7371_Y), .C0(T6835_Y),     .C1(T14987_Y), .Y(T11145_Y));
KC_OAI112_X1 T11144 ( .A(T7374_Y), .B(T7420_Y), .C0(T6835_Y),     .C1(T14989_Y), .Y(T11144_Y));
KC_OAI112_X1 T11196 ( .A(T15728_Y), .B(T7601_Y), .C0(T14989_Y),     .C1(T6803_Y), .Y(T11196_Y));
KC_OAI112_X1 T11892 ( .A(T15789_Y), .B(T16342_Y), .C0(T8688_Y),     .C1(T11010_Y), .Y(T11892_Y));
KC_OAI112_X1 T11243 ( .A(T15785_Y), .B(T7891_Y), .C0(T16463_Y),     .C1(T912_Y), .Y(T11243_Y));
KC_OAI112_X1 T11242 ( .A(T15790_Y), .B(T7871_Y), .C0(T8773_Y),     .C1(T14987_Y), .Y(T11242_Y));
KC_OAI112_X1 T11241 ( .A(T15783_Y), .B(T7897_Y), .C0(T16463_Y),     .C1(T915_Y), .Y(T11241_Y));
KC_OAI112_X1 T11240 ( .A(T15787_Y), .B(T7896_Y), .C0(T16463_Y),     .C1(T914_Y), .Y(T11240_Y));
KC_OAI112_X1 T11232 ( .A(T15790_Y), .B(T7890_Y), .C0(T16463_Y),     .C1(T913_Y), .Y(T11232_Y));
KC_OAI112_X1 T11231 ( .A(T15789_Y), .B(T7849_Y), .C0(T8773_Y),     .C1(T11010_Y), .Y(T11231_Y));
KC_OAI112_X1 T11230 ( .A(T8838_Y), .B(T8067_Y), .C0(T16318_Y),     .C1(T933_Y), .Y(T11230_Y));
KC_OAI112_X1 T11229 ( .A(T15787_Y), .B(T7852_Y), .C0(T8773_Y),     .C1(T10916_Y), .Y(T11229_Y));
KC_OAI112_X1 T11226 ( .A(T15783_Y), .B(T7807_Y), .C0(T8773_Y),     .C1(T14989_Y), .Y(T11226_Y));
KC_OAI112_X1 T11224 ( .A(T15790_Y), .B(T16338_Y), .C0(T9372_Y),     .C1(T14987_Y), .Y(T11224_Y));
KC_OAI112_X1 T11223 ( .A(T15789_Y), .B(T16343_Y), .C0(T9372_Y),     .C1(T11010_Y), .Y(T11223_Y));
KC_OAI112_X1 T11220 ( .A(T15783_Y), .B(T16339_Y), .C0(T9372_Y),     .C1(T14989_Y), .Y(T11220_Y));
KC_OAI112_X1 T11219 ( .A(T15787_Y), .B(T7808_Y), .C0(T9372_Y),     .C1(T10916_Y), .Y(T11219_Y));
KC_OAI112_X1 T11899 ( .A(T4809_Y), .B(T590_Y), .C0(T9160_Y),     .C1(T604_Q), .Y(T11899_Y));
KC_OAI112_X1 T11300 ( .A(T1837_Y), .B(T11301_Y), .C0(T11233_Y),     .C1(T1265_Q), .Y(T11300_Y));
KC_OAI112_X1 T11298 ( .A(T1840_Y), .B(T11299_Y), .C0(T11233_Y),     .C1(T1264_Q), .Y(T11298_Y));
KC_OAI112_X1 T11297 ( .A(T1836_Y), .B(T11292_Y), .C0(T11233_Y),     .C1(T1271_Q), .Y(T11297_Y));
KC_OAI112_X1 T11291 ( .A(T1420_Y), .B(T1579_Y), .C0(T598_Y),     .C1(T1593_Y), .Y(T11291_Y));
KC_OAI112_X1 T11064 ( .A(T6952_Y), .B(T6946_Y), .C0(T9316_Y),     .C1(T10883_Y), .Y(T11064_Y));
KC_OAI112_X1 T11063 ( .A(T6951_Y), .B(T6947_Y), .C0(T15740_Y),     .C1(T10883_Y), .Y(T11063_Y));
KC_OAI112_X1 T11049 ( .A(T6900_Y), .B(T6898_Y), .C0(T9318_Y),     .C1(T10883_Y), .Y(T11049_Y));
KC_OAI112_X1 T11850 ( .A(T6339_Y), .B(T7079_Y), .C0(T124_Q),     .C1(T11016_Y), .Y(T11850_Y));
KC_OAI112_X1 T11848 ( .A(T6226_Y), .B(T6328_Y), .C0(T10883_Y),     .C1(T6803_Y), .Y(T11848_Y));
KC_OAI112_X1 T12439 ( .A(T15785_Y), .B(T7687_Y), .C0(T8688_Y),     .C1(T15032_Y), .Y(T12439_Y));
KC_OAI112_X1 T11212 ( .A(T15788_Y), .B(T7686_Y), .C0(T8688_Y),     .C1(T11011_Y), .Y(T11212_Y));
KC_OAI112_X1 T11211 ( .A(T15784_Y), .B(T16346_Y), .C0(T9372_Y),     .C1(T14990_Y), .Y(T11211_Y));
KC_OAI112_X1 T11182 ( .A(T15784_Y), .B(T7559_Y), .C0(T8688_Y),     .C1(T14990_Y), .Y(T11182_Y));
KC_OAI112_X1 T11888 ( .A(T8805_Y), .B(T7644_Y), .C0(T7801_Y),     .C1(T7868_Y), .Y(T11888_Y));
KC_OAI112_X1 T11887 ( .A(T8805_Y), .B(T7563_Y), .C0(T7801_Y),     .C1(T7867_Y), .Y(T11887_Y));
KC_OAI112_X1 T11239 ( .A(T15785_Y), .B(T7805_Y), .C0(T8773_Y),     .C1(T15032_Y), .Y(T11239_Y));
KC_OAI112_X1 T11228 ( .A(T15784_Y), .B(T7851_Y), .C0(T16463_Y),     .C1(T906_Y), .Y(T11228_Y));
KC_OAI112_X1 T11225 ( .A(T15788_Y), .B(T7850_Y), .C0(T16463_Y),     .C1(T9378_Y), .Y(T11225_Y));
KC_OAI112_X1 T11222 ( .A(T15788_Y), .B(T16345_Y), .C0(T9372_Y),     .C1(T11011_Y), .Y(T11222_Y));
KC_OAI112_X1 T11221 ( .A(T15785_Y), .B(T16344_Y), .C0(T9372_Y),     .C1(T15032_Y), .Y(T11221_Y));
KC_OAI112_X1 T11216 ( .A(T15788_Y), .B(T7806_Y), .C0(T8773_Y),     .C1(T11011_Y), .Y(T11216_Y));
KC_OAI112_X1 T11215 ( .A(T15784_Y), .B(T7804_Y), .C0(T8773_Y),     .C1(T14990_Y), .Y(T11215_Y));
KC_OAI112_X1 T11267 ( .A(T1197_Y), .B(T1196_Y), .C0(T941_Y),     .C1(T1255_Y), .Y(T11267_Y));
KC_OAI112_X1 T11263 ( .A(T12720_Y), .B(T1196_Y), .C0(T9419_Y),     .C1(T8064_Y), .Y(T11263_Y));
KC_OAI112_X1 T11262 ( .A(T12452_Y), .B(T8904_Y), .C0(T8905_Y),     .C1(T8944_Y), .Y(T11262_Y));
KC_OAI112_X1 T11857 ( .A(T6274_Y), .B(T6917_Y), .C0(T896_Y),     .C1(T10907_Y), .Y(T11857_Y));
KC_OAI112_X1 T11065 ( .A(T6937_Y), .B(T819_Y), .C0(T9316_Y),     .C1(T10907_Y), .Y(T11065_Y));
KC_OAI112_X1 T11059 ( .A(T6936_Y), .B(T6939_Y), .C0(T15740_Y),     .C1(T10907_Y), .Y(T11059_Y));
KC_OAI112_X1 T11056 ( .A(T6918_Y), .B(T6915_Y), .C0(T6819_Y),     .C1(T10907_Y), .Y(T11056_Y));
KC_OAI112_X1 T11050 ( .A(T6950_Y), .B(T6899_Y), .C0(T9318_Y),     .C1(T10907_Y), .Y(T11050_Y));
KC_OAI112_X1 T11847 ( .A(T7280_Y), .B(T6038_Y), .C0(T10905_Y),     .C1(T6803_Y), .Y(T11847_Y));
KC_OAI112_X1 T11078 ( .A(T7092_Y), .B(T7090_Y), .C0(T10907_Y),     .C1(T6803_Y), .Y(T11078_Y));
KC_OAI112_X1 T11077 ( .A(T7091_Y), .B(T842_Y), .C0(T124_Q),     .C1(T10883_Y), .Y(T11077_Y));
KC_OAI112_X1 T11076 ( .A(T7111_Y), .B(T839_Y), .C0(T124_Q),     .C1(T10907_Y), .Y(T11076_Y));
KC_OAI112_X1 T11073 ( .A(T7049_Y), .B(T7045_Y), .C0(T6835_Y),     .C1(T10883_Y), .Y(T11073_Y));
KC_OAI112_X1 T11072 ( .A(T6269_Y), .B(T7043_Y), .C0(T6835_Y),     .C1(T10907_Y), .Y(T11072_Y));
KC_OAI112_X1 T11905 ( .A(T6738_Y), .B(T11860_Y), .C0(T9306_Y),     .C1(T6619_Y), .Y(T11905_Y));
KC_OAI112_X1 T11902 ( .A(T6734_Y), .B(T11908_Y), .C0(T9305_Y),     .C1(T6620_Y), .Y(T11902_Y));
KC_OAI112_X1 T11901 ( .A(T6735_Y), .B(T11861_Y), .C0(T9304_Y),     .C1(T6621_Y), .Y(T11901_Y));
KC_OAI112_X1 T11104 ( .A(T7281_Y), .B(T7291_Y), .C0(T124_Q),     .C1(T10905_Y), .Y(T11104_Y));
KC_OAI112_X1 T11103 ( .A(T7259_Y), .B(T867_Y), .C0(T9316_Y),     .C1(T10905_Y), .Y(T11103_Y));
KC_OAI112_X1 T11102 ( .A(T7279_Y), .B(T7295_Y), .C0(T9318_Y),     .C1(T10905_Y), .Y(T11102_Y));
KC_OAI112_X1 T11101 ( .A(T7261_Y), .B(T7238_Y), .C0(T896_Y),     .C1(T10905_Y), .Y(T11101_Y));
KC_OAI112_X1 T11093 ( .A(T7278_Y), .B(T7297_Y), .C0(T6819_Y),     .C1(T10905_Y), .Y(T11093_Y));
KC_OAI112_X1 T11092 ( .A(T7260_Y), .B(T7276_Y), .C0(T15740_Y),     .C1(T10905_Y), .Y(T11092_Y));
KC_OAI112_X1 T11091 ( .A(T7262_Y), .B(T7292_Y), .C0(T6835_Y),     .C1(T10905_Y), .Y(T11091_Y));
KC_OAI112_X1 T11164 ( .A(T12404_Y), .B(T6647_Y), .C0(T731_Y),     .C1(T15413_Y), .Y(T11164_Y));
KC_OAI112_X1 T11163 ( .A(T12397_Y), .B(T7434_Y), .C0(T728_Y),     .C1(T573_Y), .Y(T11163_Y));
KC_OAI112_X1 T11162 ( .A(T15744_Y), .B(T11155_Y), .C0(T573_Y),     .C1(T731_Y), .Y(T11162_Y));
KC_OAI112_X1 T11156 ( .A(T12428_Y), .B(T11157_Y), .C0(T6803_Y),     .C1(T10918_Y), .Y(T11156_Y));
KC_OAI112_X1 T11143 ( .A(T9370_Y), .B(T549_Y), .C0(T15749_Y),     .C1(T7839_Y), .Y(T11143_Y));
KC_OAI112_X1 T11141 ( .A(T12396_Y), .B(T7354_Y), .C0(T728_Y),     .C1(T15413_Y), .Y(T11141_Y));
KC_OAI112_X1 T11140 ( .A(T8656_Y), .B(T15223_Y), .C0(T11087_Y),     .C1(T1131_Q), .Y(T11140_Y));
KC_OAI112_X1 T11139 ( .A(T9370_Y), .B(T6691_Y), .C0(T15748_Y),     .C1(T7839_Y), .Y(T11139_Y));
KC_OAI112_X1 T8396 ( .A(T8713_Y), .B(T8725_Y), .C0(T5343_Q),     .C1(T16091_Y), .Y(T8396_Y));
KC_OAI112_X1 T11201 ( .A(T12436_Y), .B(T7639_Y), .C0(T728_Y),     .C1(T702_Y), .Y(T11201_Y));
KC_OAI112_X1 T11200 ( .A(T8715_Y), .B(T8725_Y), .C0(T5360_Q),     .C1(T16092_Y), .Y(T11200_Y));
KC_OAI112_X1 T11199 ( .A(T727_Y), .B(T9370_Y), .C0(T12434_Y),     .C1(T7839_Y), .Y(T11199_Y));
KC_OAI112_X1 T11197 ( .A(T9370_Y), .B(T9374_Y), .C0(T12431_Y),     .C1(T7839_Y), .Y(T11197_Y));
KC_OAI112_X1 T11192 ( .A(T9370_Y), .B(T9373_Y), .C0(T12420_Y),     .C1(T7839_Y), .Y(T11192_Y));
KC_OAI112_X1 T11191 ( .A(T12421_Y), .B(T7586_Y), .C0(T731_Y),     .C1(T651_Y), .Y(T11191_Y));
KC_OAI112_X1 T11190 ( .A(T15743_Y), .B(T6649_Y), .C0(T728_Y),     .C1(T651_Y), .Y(T11190_Y));
KC_OAI112_X1 T11177 ( .A(T12433_Y), .B(T7552_Y), .C0(T731_Y),     .C1(T702_Y), .Y(T11177_Y));
KC_OAI112_X1 T11894 ( .A(T7876_Y), .B(T937_Y), .C0(T1458_Y),     .C1(T8938_Y), .Y(T11894_Y));
KC_OAI112_X1 T11906 ( .A(T6744_Y), .B(T11909_Y), .C0(T9309_Y),     .C1(T6795_Y), .Y(T11906_Y));
KC_OAI112_X1 T11903 ( .A(T6743_Y), .B(T11862_Y), .C0(T9508_Y),     .C1(T5703_Y), .Y(T11903_Y));
KC_OAI112_X1 T11917 ( .A(T9301_Y), .B(T8725_Y), .C0(T1084_Q),     .C1(T15779_Y), .Y(T11917_Y));
KC_OAI112_X1 T11170 ( .A(T8670_Y), .B(T8725_Y), .C0(T15775_Y),     .C1(T5359_Q), .Y(T11170_Y));
KC_OAI112_X1 T11138 ( .A(T6826_Y), .B(T8725_Y), .C0(T5297_Q),     .C1(T15777_Y), .Y(T11138_Y));
KC_OAI112_X1 T11281 ( .A(T10698_Y), .B(T10723_Y), .C0(T8974_Y),     .C1(T8032_Y), .Y(T11281_Y));
KC_OAI112_X1 T11280 ( .A(T1126_Y), .B(T1196_Y), .C0(T1458_Y),     .C1(T980_Q), .Y(T11280_Y));
KC_OAI112_X1 T6754 ( .A(T5028_Y), .B(T14940_Q), .C0(T6784_Y),     .C1(T6765_Y), .Y(T6754_Y));
KC_OAI112_X1 T11957 ( .A(T11945_Y), .B(T10484_Y), .C0(T6784_Y),     .C1(T15398_Y), .Y(T11957_Y));
KC_OAI112_X1 T11956 ( .A(T11922_Y), .B(T10355_Y), .C0(T6786_Y),     .C1(T15398_Y), .Y(T11956_Y));
KC_OAI112_X1 T11923 ( .A(T5649_Y), .B(T5028_Y), .C0(T13710_Q),     .C1(T1637_Y), .Y(T11923_Y));
KC_OAI112_X1 T11922 ( .A(T5028_Y), .B(T6594_Q), .C0(T6787_Y),     .C1(T6765_Y), .Y(T11922_Y));
KC_OAI112_X1 T11921 ( .A(T11920_Y), .B(T10354_Y), .C0(T6787_Y),     .C1(T15398_Y), .Y(T11921_Y));
KC_OAI112_X1 T11920 ( .A(T5028_Y), .B(T13732_Q), .C0(T15666_Y),     .C1(T6765_Y), .Y(T11920_Y));
KC_OAI112_X1 T11919 ( .A(T10412_Y), .B(T5647_Y), .C0(T15398_Y),     .C1(T15666_Y), .Y(T11919_Y));
KC_OAI112_X1 T11137 ( .A(T5028_Y), .B(T14773_Q), .C0(T457_Y),     .C1(T6765_Y), .Y(T11137_Y));
KC_OAI112_X1 T11136 ( .A(T5028_Y), .B(T14769_Q), .C0(T496_Y),     .C1(T6765_Y), .Y(T11136_Y));
KC_OAI112_X1 T11134 ( .A(T11137_Y), .B(T9658_Y), .C0(T496_Y),     .C1(T15398_Y), .Y(T11134_Y));
KC_OAI112_X1 T11128 ( .A(T11127_Y), .B(T9659_Y), .C0(T457_Y),     .C1(T15398_Y), .Y(T11128_Y));
KC_OAI112_X1 T11127 ( .A(T5028_Y), .B(T13777_Q), .C0(T15401_Y),     .C1(T6765_Y), .Y(T11127_Y));
KC_OAI112_X1 T11117 ( .A(T5028_Y), .B(T14939_Q), .C0(T417_Y),     .C1(T6765_Y), .Y(T11117_Y));
KC_OAI112_X1 T11915 ( .A(T10308_Y), .B(T13040_Y), .C0(T10032_Y),     .C1(T15087_Y), .Y(T11915_Y));
KC_OAI112_X1 T11261 ( .A(T15811_Y), .B(T7922_Y), .C0(T16371_Y),     .C1(T5364_Q), .Y(T11261_Y));
KC_OAI112_X1 T11254 ( .A(T15811_Y), .B(T7982_Y), .C0(T16371_Y),     .C1(T16433_Q), .Y(T11254_Y));
KC_OAI112_X1 T11253 ( .A(T15811_Y), .B(T7984_Y), .C0(T16371_Y),     .C1(T8877_Q), .Y(T11253_Y));
KC_OAI112_X1 T11252 ( .A(T10309_Y), .B(T13040_Y), .C0(T10305_Y),     .C1(T15069_Y), .Y(T11252_Y));
KC_OAI112_X1 T11251 ( .A(T15811_Y), .B(T7924_Y), .C0(T16371_Y),     .C1(T1707_Q), .Y(T11251_Y));
KC_OAI112_X1 T11250 ( .A(T15811_Y), .B(T7981_Y), .C0(T16371_Y),     .C1(T1717_Q), .Y(T11250_Y));
KC_OAI112_X1 T11249 ( .A(T15811_Y), .B(T7980_Y), .C0(T16371_Y),     .C1(T8880_Q), .Y(T11249_Y));
KC_OAI112_X1 T11248 ( .A(T15811_Y), .B(T7921_Y), .C0(T16371_Y),     .C1(T16413_Q), .Y(T11248_Y));
KC_OAI112_X1 T11289 ( .A(T15811_Y), .B(T10702_Y), .C0(T1533_Y),     .C1(T9970_Y), .Y(T11289_Y));
KC_OAI112_X1 T11288 ( .A(T15811_Y), .B(T10742_Y), .C0(T15519_Y),     .C1(T9970_Y), .Y(T11288_Y));
KC_OAI112_X1 T11286 ( .A(T15811_Y), .B(T10700_Y), .C0(T1532_Y),     .C1(T9970_Y), .Y(T11286_Y));
KC_OAI112_X1 T11279 ( .A(T15811_Y), .B(T7923_Y), .C0(T1517_Y),     .C1(T9970_Y), .Y(T11279_Y));
KC_OAI112_X1 T11278 ( .A(T15811_Y), .B(T10701_Y), .C0(T1519_Y),     .C1(T9970_Y), .Y(T11278_Y));
KC_OAI112_X1 T11481 ( .A(T10225_Y), .B(T16156_Y), .C0(T10207_Y),     .C1(T10224_Y), .Y(T11481_Y));
KC_OAI112_X1 T11602 ( .A(T5493_Y), .B(T6766_Y), .C0(T6121_Y),     .C1(T1786_Y), .Y(T11602_Y));
KC_OAI112_X1 T11601 ( .A(T8311_Y), .B(T1784_Y), .C0(T6121_Y),     .C1(T2246_Y), .Y(T11601_Y));
KC_OAI112_X1 T11600 ( .A(T4961_Y), .B(T2307_Y), .C0(T6005_Y),     .C1(T6121_Y), .Y(T11600_Y));
KC_OAI112_X1 T11669 ( .A(T8375_Y), .B(T1799_Y), .C0(T6121_Y),     .C1(T16042_Y), .Y(T11669_Y));
KC_OAI112_X1 T11668 ( .A(T1796_Y), .B(T6388_Y), .C0(T6121_Y),     .C1(T2250_Y), .Y(T11668_Y));
KC_OAI112_X1 T11667 ( .A(T1798_Y), .B(T6387_Y), .C0(T6121_Y),     .C1(T2279_Y), .Y(T11667_Y));
KC_OAI112_X1 T11654 ( .A(T8511_Y), .B(T1801_Y), .C0(T6121_Y),     .C1(T2245_Y), .Y(T11654_Y));
KC_OAI112_X1 T11653 ( .A(T1802_Y), .B(T1794_Y), .C0(T1805_Y),     .C1(T6184_Y), .Y(T11653_Y));
KC_OAI112_X1 T11701 ( .A(T1817_Y), .B(T1808_Y), .C0(T1804_Y),     .C1(T15618_Y), .Y(T11701_Y));
KC_OAI112_X1 T11691 ( .A(T5505_Y), .B(T1811_Y), .C0(T1805_Y),     .C1(T15618_Y), .Y(T11691_Y));
KC_OAI112_X1 T11954 ( .A(T2449_Y), .B(T14840_Q), .C0(T629_Y),     .C1(T2448_Y), .Y(T11954_Y));
KC_OAI112_X1 T11133 ( .A(T11121_Y), .B(T9682_Y), .C0(T487_Y),     .C1(T6592_Y), .Y(T11133_Y));
KC_OAI112_X1 T11126 ( .A(T11120_Y), .B(T9684_Y), .C0(T15405_Y),     .C1(T15398_Y), .Y(T11126_Y));
KC_OAI112_X1 T11125 ( .A(T2449_Y), .B(T13758_Q), .C0(T487_Y),     .C1(T2448_Y), .Y(T11125_Y));
KC_OAI112_X1 T11124 ( .A(T2449_Y), .B(T13771_Q), .C0(T484_Y),     .C1(T2448_Y), .Y(T11124_Y));
KC_OAI112_X1 T11123 ( .A(T11124_Y), .B(T9683_Y), .C0(T448_Y),     .C1(T6592_Y), .Y(T11123_Y));
KC_OAI112_X1 T11122 ( .A(T11119_Y), .B(T9685_Y), .C0(T493_Y),     .C1(T15398_Y), .Y(T11122_Y));
KC_OAI112_X1 T11121 ( .A(T5028_Y), .B(T13774_Q), .C0(T15405_Y),     .C1(T6765_Y), .Y(T11121_Y));
KC_OAI112_X1 T11120 ( .A(T5028_Y), .B(T13776_Q), .C0(T493_Y),     .C1(T6765_Y), .Y(T11120_Y));
KC_OAI112_X1 T11119 ( .A(T2449_Y), .B(T13775_Q), .C0(T448_Y),     .C1(T6765_Y), .Y(T11119_Y));
KC_OAI112_X1 T11113 ( .A(T2449_Y), .B(T14771_Q), .C0(T6460_Y),     .C1(T2448_Y), .Y(T11113_Y));
KC_OAI112_X1 T11112 ( .A(T2449_Y), .B(T13746_Q), .C0(T410_Y),     .C1(T2448_Y), .Y(T11112_Y));
KC_OAI112_X1 T11111 ( .A(T11114_Y), .B(T10441_Y), .C0(T484_Y),     .C1(T6592_Y), .Y(T11111_Y));
KC_OAI112_X1 T11943 ( .A(T11935_Y), .B(T10482_Y), .C0(T6783_Y),     .C1(T15398_Y), .Y(T11943_Y));
KC_OAI112_X1 T11941 ( .A(T5028_Y), .B(T14932_Q), .C0(T15421_Y),     .C1(T6765_Y), .Y(T11941_Y));
KC_OAI112_X1 T11940 ( .A(T11941_Y), .B(T9755_Y), .C0(T623_Y),     .C1(T15398_Y), .Y(T11940_Y));
KC_OAI112_X1 T11939 ( .A(T11937_Y), .B(T10481_Y), .C0(T15421_Y),     .C1(T15398_Y), .Y(T11939_Y));
KC_OAI112_X1 T11938 ( .A(T5028_Y), .B(T13896_Q), .C0(T6783_Y),     .C1(T6765_Y), .Y(T11938_Y));
KC_OAI112_X1 T11260 ( .A(T9966_Y), .B(T10515_Y), .C0(T2161_Q),     .C1(T868_Y), .Y(T11260_Y));
KC_OAI112_X1 T11290 ( .A(T2030_Y), .B(T16293_Y), .C0(T2031_Y),     .C1(T15814_Y), .Y(T11290_Y));
KC_OAI112_X1 T11287 ( .A(T15811_Y), .B(T4906_Y), .C0(T15512_Y),     .C1(T9970_Y), .Y(T11287_Y));
KC_OAI112_X1 T11284 ( .A(T10061_Y), .B(T12734_Y), .C0(T5369_Y),     .C1(T10078_Y), .Y(T11284_Y));
KC_OAI112_X1 T11283 ( .A(T15811_Y), .B(T1686_Y), .C0(T15511_Y),     .C1(T9970_Y), .Y(T11283_Y));
KC_OAI112_X1 T11282 ( .A(T2039_Y), .B(T2604_Y), .C0(T2036_Y),     .C1(T2001_Q), .Y(T11282_Y));
KC_OAI112_X1 T11465 ( .A(T2086_Y), .B(T2138_Y), .C0(T15574_Y),     .C1(T5898_Y), .Y(T11465_Y));
KC_OAI112_X1 T11435 ( .A(T2084_Y), .B(T2087_Y), .C0(T15566_Y),     .C1(T15574_Y), .Y(T11435_Y));
KC_OAI112_X1 T11528 ( .A(T12211_Y), .B(T2166_Y), .C0(T5898_Y),     .C1(T15942_Y), .Y(T11528_Y));
KC_OAI112_X1 T11595 ( .A(T5474_Q), .B(T15943_Y), .C0(T6515_Y),     .C1(T5902_Y), .Y(T11595_Y));
KC_OAI112_X1 T11594 ( .A(T1777_Q), .B(T15943_Y), .C0(T6515_Y),     .C1(T5878_Y), .Y(T11594_Y));
KC_OAI112_X1 T11584 ( .A(T2192_Y), .B(T2773_Y), .C0(T2802_Y),     .C1(T5982_Y), .Y(T11584_Y));
KC_OAI112_X1 T11583 ( .A(T2195_Y), .B(T11569_Y), .C0(T2250_Y),     .C1(T12064_Y), .Y(T11583_Y));
KC_OAI112_X1 T11599 ( .A(T2197_Y), .B(T2231_Y), .C0(T5902_Y),     .C1(T2802_Y), .Y(T11599_Y));
KC_OAI112_X1 T12050 ( .A(T2285_Y), .B(T6404_Y), .C0(T6185_Y),     .C1(T2280_Y), .Y(T12050_Y));
KC_OAI112_X1 T11634 ( .A(T2222_Y), .B(T2847_Y), .C0(T4968_Y),     .C1(T6000_Y), .Y(T11634_Y));
KC_OAI112_X1 T11732 ( .A(T2287_Y), .B(T6816_Y), .C0(T6185_Y),     .C1(T16042_Y), .Y(T11732_Y));
KC_OAI112_X1 T11690 ( .A(T2272_Y), .B(T2308_Y), .C0(T1805_Y),     .C1(T6121_Y), .Y(T11690_Y));
KC_OAI112_X1 T11811 ( .A(T12101_Y), .B(T12107_Y), .C0(T10573_Y),     .C1(T10558_Y), .Y(T11811_Y));
KC_OAI112_X1 T11824 ( .A(T6543_Y), .B(T11772_Y), .C0(T1856_Q),     .C1(T6542_Y), .Y(T11824_Y));
KC_OAI112_X1 T11034 ( .A(T2372_Y), .B(T2362_Y), .C0(T11775_Y),     .C1(T11826_Y), .Y(T11034_Y));
KC_OAI112_X1 T11924 ( .A(T11109_Y), .B(T10439_Y), .C0(T376_Y),     .C1(T6592_Y), .Y(T11924_Y));
KC_OAI112_X1 T11953 ( .A(T11927_Y), .B(T8528_Y), .C0(T6774_Y),     .C1(T6592_Y), .Y(T11953_Y));
KC_OAI112_X1 T11952 ( .A(T11950_Y), .B(T8529_Y), .C0(T6763_Y),     .C1(T6592_Y), .Y(T11952_Y));
KC_OAI112_X1 T11951 ( .A(T5028_Y), .B(T14936_Q), .C0(T6774_Y),     .C1(T6765_Y), .Y(T11951_Y));
KC_OAI112_X1 T11950 ( .A(T2449_Y), .B(T14935_Q), .C0(T6764_Y),     .C1(T2448_Y), .Y(T11950_Y));
KC_OAI112_X1 T11131 ( .A(T11118_Y), .B(T9676_Y), .C0(T15404_Y),     .C1(T6592_Y), .Y(T11131_Y));
KC_OAI112_X1 T11130 ( .A(T11115_Y), .B(T9675_Y), .C0(T405_Y),     .C1(T6592_Y), .Y(T11130_Y));
KC_OAI112_X1 T11118 ( .A(T2449_Y), .B(T13772_Q), .C0(T488_Y),     .C1(T2448_Y), .Y(T11118_Y));
KC_OAI112_X1 T11115 ( .A(T2449_Y), .B(T13773_Q), .C0(T15404_Y),     .C1(T2448_Y), .Y(T11115_Y));
KC_OAI112_X1 T11110 ( .A(T2449_Y), .B(T13654_Q), .C0(T376_Y),     .C1(T2448_Y), .Y(T11110_Y));
KC_OAI112_X1 T11109 ( .A(T2449_Y), .B(T13783_Q), .C0(T405_Y),     .C1(T2448_Y), .Y(T11109_Y));
KC_OAI112_X1 T11946 ( .A(T2674_Y), .B(T11948_Y), .C0(T16093_Y),     .C1(T610_Y), .Y(T11946_Y));
KC_OAI112_X1 T11932 ( .A(T2449_Y), .B(T14836_Q), .C0(T632_Y),     .C1(T2448_Y), .Y(T11932_Y));
KC_OAI112_X1 T11931 ( .A(T14933_Q), .B(T2449_Y), .C0(T6763_Y),     .C1(T2448_Y), .Y(T11931_Y));
KC_OAI112_X1 T11930 ( .A(T5028_Y), .B(T14838_Q), .C0(T623_Y),     .C1(T6765_Y), .Y(T11930_Y));
KC_OAI112_X1 T11176 ( .A(T2459_Y), .B(T2674_Y), .C0(T12080_Y),     .C1(T9774_Y), .Y(T11176_Y));
KC_OAI112_X1 T11174 ( .A(T9778_Y), .B(T11173_Y), .C0(T2480_Y),     .C1(T611_Y), .Y(T11174_Y));
KC_OAI112_X1 T11173 ( .A(T611_Y), .B(T4986_Y), .C0(T2454_Y),     .C1(T2476_Y), .Y(T11173_Y));
KC_OAI112_X1 T11172 ( .A(T2481_Y), .B(T2674_Y), .C0(T9772_Y),     .C1(T11174_Y), .Y(T11172_Y));
KC_OAI112_X1 T11359 ( .A(T11014_Y), .B(T15754_Y), .C0(T5427_Y),     .C1(T5758_Y), .Y(T11359_Y));
KC_OAI112_X1 T11327 ( .A(T2656_Y), .B(T6037_Y), .C0(T2675_Y),     .C1(T14954_Q), .Y(T11327_Y));
KC_OAI112_X1 T11471 ( .A(T2171_Y), .B(T2145_Y), .C0(T2754_Y),     .C1(T5875_Y), .Y(T11471_Y));
KC_OAI112_X1 T11470 ( .A(T2171_Y), .B(T2140_Y), .C0(T2754_Y),     .C1(T5908_Y), .Y(T11470_Y));
KC_OAI112_X1 T11478 ( .A(T2173_Y), .B(T2188_Y), .C0(T2189_Y),     .C1(T6212_Y), .Y(T11478_Y));
KC_OAI112_X1 T11619 ( .A(T2795_Y), .B(T4956_Y), .C0(T6055_Y),     .C1(T2802_Y), .Y(T11619_Y));
KC_OAI112_X1 T11648 ( .A(T2828_Y), .B(T2284_Y), .C0(T12347_Y),     .C1(T2854_Y), .Y(T11648_Y));
KC_OAI112_X1 T11726 ( .A(T12066_Y), .B(T10976_Y), .C0(T3408_Y),     .C1(T16105_Y), .Y(T11726_Y));
KC_OAI112_X1 T11698 ( .A(T12359_Y), .B(T2858_Y), .C0(T6161_Y),     .C1(T11598_Y), .Y(T11698_Y));
KC_OAI112_X1 T11697 ( .A(T6493_Y), .B(T6120_Y), .C0(T6140_Y),     .C1(T3429_Y), .Y(T11697_Y));
KC_OAI112_X1 T11696 ( .A(T12359_Y), .B(T6161_Y), .C0(T5523_Y),     .C1(T12039_Y), .Y(T11696_Y));
KC_OAI112_X1 T11686 ( .A(T12972_Y), .B(T5000_Y), .C0(T6087_Y),     .C1(T2863_Y), .Y(T11686_Y));
KC_OAI112_X1 T11685 ( .A(T10572_Y), .B(T6532_Y), .C0(T4705_Y),     .C1(T2866_Y), .Y(T11685_Y));
KC_OAI112_X1 T12061 ( .A(T11806_Y), .B(T10559_Y), .C0(T6101_Y),     .C1(T10561_Y), .Y(T12061_Y));
KC_OAI112_X1 T11805 ( .A(T12366_Y), .B(T6581_Y), .C0(T12064_Y),     .C1(T6120_Y), .Y(T11805_Y));
KC_OAI112_X1 T11783 ( .A(T12305_Y), .B(T4144_Y), .C0(T12871_Y),     .C1(T2865_Y), .Y(T11783_Y));
KC_OAI112_X1 T11767 ( .A(T6224_Y), .B(T2890_Y), .C0(T6229_Y),     .C1(T10988_Y), .Y(T11767_Y));
KC_OAI112_X1 T11740 ( .A(T2909_Y), .B(T2907_Y), .C0(T5518_Y),     .C1(T15633_Y), .Y(T11740_Y));
KC_OAI112_X1 T11040 ( .A(T6221_Y), .B(T6561_Y), .C0(T2912_Y),     .C1(T10986_Y), .Y(T11040_Y));
KC_OAI112_X1 T11039 ( .A(T2916_Y), .B(T12468_Y), .C0(T12067_Y),     .C1(T290_Y), .Y(T11039_Y));
KC_OAI112_X1 T11820 ( .A(T2916_Y), .B(T2928_Y), .C0(T2937_Y),     .C1(T6537_Y), .Y(T11820_Y));
KC_OAI112_X1 T11819 ( .A(T2939_Y), .B(T11040_Y), .C0(T2937_Y),     .C1(T6530_Y), .Y(T11819_Y));
KC_OAI112_X1 T11175 ( .A(T3045_Y), .B(T3045_Y), .C0(T15420_Y),     .C1(T2496_Y), .Y(T11175_Y));
KC_OAI112_X1 T11354 ( .A(T6059_Y), .B(T3819_Y), .C0(T3816_Y),     .C1(T3840_Y), .Y(T11354_Y));
KC_OAI112_X1 T11319 ( .A(T3823_Y), .B(T5435_Y), .C0(T5101_Y),     .C1(T11988_Y), .Y(T11319_Y));
KC_OAI112_X1 T11468 ( .A(T3250_Y), .B(T15129_Y), .C0(T3260_Y),     .C1(T15929_Y), .Y(T11468_Y));
KC_OAI112_X1 T11446 ( .A(T5445_Y), .B(T15945_Y), .C0(T4471_Y),     .C1(T5892_Y), .Y(T11446_Y));
KC_OAI112_X1 T11445 ( .A(T11522_Y), .B(T3247_Y), .C0(T4471_Y),     .C1(T5907_Y), .Y(T11445_Y));
KC_OAI112_X1 T11485 ( .A(T3314_Y), .B(T3292_Y), .C0(T2122_Y),     .C1(T11487_Y), .Y(T11485_Y));
KC_OAI112_X1 T11557 ( .A(T3326_Y), .B(T3323_Y), .C0(T3326_Y),     .C1(T15980_Y), .Y(T11557_Y));
KC_OAI112_X1 T11544 ( .A(T3332_Y), .B(T3343_Y), .C0(T3344_Y),     .C1(T3333_Y), .Y(T11544_Y));
KC_OAI112_X1 T11673 ( .A(T6393_Y), .B(T3392_Y), .C0(T3516_Y),     .C1(T11677_Y), .Y(T11673_Y));
KC_OAI112_X1 T11672 ( .A(T6086_Y), .B(T3386_Y), .C0(T3380_Y),     .C1(T5523_Y), .Y(T11672_Y));
KC_OAI112_X1 T11628 ( .A(T4179_Q), .B(T4176_Q), .C0(T4035_Y),     .C1(T15760_Q), .Y(T11628_Y));
KC_OAI112_X1 T11721 ( .A(T6177_Y), .B(T3422_Y), .C0(T10975_Y),     .C1(T6138_Y), .Y(T11721_Y));
KC_OAI112_X1 T11720 ( .A(T2878_Q), .B(T11002_Y), .C0(T16039_Y),     .C1(T16138_Y), .Y(T11720_Y));
KC_OAI112_X1 T11718 ( .A(T11720_Y), .B(T6179_Y), .C0(T3372_Y),     .C1(T15802_Q), .Y(T11718_Y));
KC_OAI112_X1 T11717 ( .A(T16107_Y), .B(T10610_Y), .C0(T6236_Y),     .C1(T5046_Y), .Y(T11717_Y));
KC_OAI112_X1 T11716 ( .A(T5522_Y), .B(T6160_Y), .C0(T4016_Y),     .C1(T6236_Y), .Y(T11716_Y));
KC_OAI112_X1 T11702 ( .A(T3420_Y), .B(T3450_Y), .C0(T5522_Y),     .C1(T3454_Y), .Y(T11702_Y));
KC_OAI112_X1 T11694 ( .A(T6532_Y), .B(T10611_Y), .C0(T6179_Y),     .C1(T12280_Y), .Y(T11694_Y));
KC_OAI112_X1 T11689 ( .A(T10609_Y), .B(T12848_Y), .C0(T6176_Y),     .C1(T10608_Y), .Y(T11689_Y));
KC_OAI112_X1 T11683 ( .A(T6831_Y), .B(T12257_Y), .C0(T3445_Y),     .C1(T12466_Y), .Y(T11683_Y));
KC_OAI112_X1 T11799 ( .A(T6584_Y), .B(T3472_Y), .C0(T12363_Y),     .C1(T2865_Y), .Y(T11799_Y));
KC_OAI112_X1 T11798 ( .A(T12309_Y), .B(T12872_Y), .C0(T10609_Y),     .C1(T6120_Y), .Y(T11798_Y));
KC_OAI112_X1 T11797 ( .A(T3444_Y), .B(T5521_Y), .C0(T3443_Y),     .C1(T6215_Y), .Y(T11797_Y));
KC_OAI112_X1 T11763 ( .A(T12300_Y), .B(T11684_Y), .C0(T6208_Y),     .C1(T3528_Q), .Y(T11763_Y));
KC_OAI112_X1 T11737 ( .A(T3491_Y), .B(T6213_Y), .C0(T8403_Y),     .C1(T2888_Y), .Y(T11737_Y));
KC_OAI112_X1 T11350 ( .A(T3842_Y), .B(T3800_Y), .C0(T4486_Y),     .C1(T15868_Y), .Y(T11350_Y));
KC_OAI112_X1 T11330 ( .A(T8185_Y), .B(T10885_Y), .C0(T3840_Y),     .C1(T3841_Y), .Y(T11330_Y));
KC_OAI112_X1 T11324 ( .A(T12788_Y), .B(T8179_Y), .C0(T5101_Y),     .C1(T145_Q), .Y(T11324_Y));
KC_OAI112_X1 T11323 ( .A(T10889_Y), .B(T3792_Y), .C0(T3840_Y),     .C1(T3802_Y), .Y(T11323_Y));
KC_OAI112_X1 T11315 ( .A(T12788_Y), .B(T10894_Y), .C0(T5840_Y),     .C1(T15869_Y), .Y(T11315_Y));
KC_OAI112_X1 T11314 ( .A(T3820_Y), .B(T3817_Y), .C0(T5789_Y),     .C1(T12129_Y), .Y(T11314_Y));
KC_OAI112_X1 T11424 ( .A(T11425_Y), .B(T15012_Y), .C0(T3850_Y),     .C1(T8188_Y), .Y(T11424_Y));
KC_OAI112_X1 T11423 ( .A(T6108_Y), .B(T3796_Y), .C0(T3825_Y),     .C1(T8204_Y), .Y(T11423_Y));
KC_OAI112_X1 T11374 ( .A(T11378_Y), .B(T16153_Y), .C0(T11381_Y),     .C1(T11428_Y), .Y(T11374_Y));
KC_OAI112_X1 T11373 ( .A(T8451_Y), .B(T12797_Y), .C0(T4461_Y),     .C1(T8193_Y), .Y(T11373_Y));
KC_OAI112_X1 T11366 ( .A(T5788_Y), .B(T3856_Y), .C0(T13296_Y),     .C1(T3837_Y), .Y(T11366_Y));
KC_OAI112_X1 T11467 ( .A(T3859_Y), .B(T6228_Y), .C0(T15571_Y),     .C1(T4471_Y), .Y(T11467_Y));
KC_OAI112_X1 T11443 ( .A(T5105_Y), .B(T10898_Y), .C0(T8213_Y),     .C1(T8445_Y), .Y(T11443_Y));
KC_OAI112_X1 T11434 ( .A(T11522_Y), .B(T3863_Y), .C0(T4968_Y),     .C1(T4471_Y), .Y(T11434_Y));
KC_OAI112_X1 T15956 ( .A(T3965_Q), .B(T11556_Y), .C0(T5989_Y),     .C1(T11587_Y), .Y(T15956_Y));
KC_OAI112_X1 T11510 ( .A(T3965_Q), .B(T11476_Y), .C0(T3919_Y),     .C1(T5986_Y), .Y(T11510_Y));
KC_OAI112_X1 T11509 ( .A(T11503_Y), .B(T3931_Y), .C0(T5120_Y),     .C1(T11514_Y), .Y(T11509_Y));
KC_OAI112_X1 T12017 ( .A(T3980_Y), .B(T3941_Y), .C0(T3975_Y),     .C1(T8290_Y), .Y(T12017_Y));
KC_OAI112_X1 T12035 ( .A(T2853_Y), .B(T3417_Y), .C0(T4058_Y),     .C1(T12039_Y), .Y(T12035_Y));
KC_OAI112_X1 T11688 ( .A(T10579_Y), .B(T10578_Y), .C0(T3458_Y),     .C1(T16141_Y), .Y(T11688_Y));
KC_OAI112_X1 T11687 ( .A(T10882_Y), .B(T4100_Y), .C0(T4074_Y),     .C1(T4083_Y), .Y(T11687_Y));
KC_OAI112_X1 T11682 ( .A(T4090_Y), .B(T5110_Y), .C0(T4076_Y),     .C1(T8373_Y), .Y(T11682_Y));
KC_OAI112_X1 T11792 ( .A(T12255_Y), .B(T4111_Y), .C0(T10580_Y),     .C1(T16143_Y), .Y(T11792_Y));
KC_OAI112_X1 T11791 ( .A(T4117_Y), .B(T12055_Y), .C0(T6155_Y),     .C1(T12361_Y), .Y(T11791_Y));
KC_OAI112_X1 T11790 ( .A(T2895_Y), .B(T4114_Y), .C0(T5049_Y),     .C1(T5135_Y), .Y(T11790_Y));
KC_OAI112_X1 T11789 ( .A(T11803_Y), .B(T4116_Y), .C0(T5051_Y),     .C1(T6175_Y), .Y(T11789_Y));
KC_OAI112_X1 T11780 ( .A(T11803_Y), .B(T6535_Y), .C0(T5051_Y),     .C1(T6043_Y), .Y(T11780_Y));
KC_OAI112_X1 T11760 ( .A(T4130_Y), .B(T12303_Y), .C0(T6557_Y),     .C1(T6549_Q), .Y(T11760_Y));
KC_OAI112_X1 T11735 ( .A(T4090_Y), .B(T4129_Y), .C0(T10580_Y),     .C1(T15640_Y), .Y(T11735_Y));
KC_OAI112_X1 T11035 ( .A(T3493_Y), .B(T4134_Y), .C0(T12295_Y),     .C1(T2865_Y), .Y(T11035_Y));
KC_OAI112_X1 T11972 ( .A(T4449_Y), .B(T15872_Y), .C0(T4383_Y),     .C1(T14942_Q), .Y(T11972_Y));
KC_OAI112_X1 T11344 ( .A(T12791_Y), .B(T11013_Y), .C0(T4387_Y),     .C1(T5824_Y), .Y(T11344_Y));
KC_OAI112_X1 T11311 ( .A(T11975_Y), .B(T3842_Y), .C0(T4383_Y),     .C1(T144_Q), .Y(T11311_Y));
KC_OAI112_X1 T11310 ( .A(T3825_Y), .B(T12953_Y), .C0(T5789_Y),     .C1(T14942_Q), .Y(T11310_Y));
KC_OAI112_X1 T11418 ( .A(T6117_Y), .B(T4434_Y), .C0(T5789_Y),     .C1(T12173_Y), .Y(T11418_Y));
KC_OAI112_X1 T11399 ( .A(T15872_Y), .B(T4437_Y), .C0(T4388_Y),     .C1(T4432_Y), .Y(T11399_Y));
KC_OAI112_X1 T11398 ( .A(T4444_Y), .B(T4383_Y), .C0(T4452_Y),     .C1(T4439_Y), .Y(T11398_Y));
KC_OAI112_X1 T11388 ( .A(T10914_Y), .B(T5816_Y), .C0(T5788_Y),     .C1(T4439_Y), .Y(T11388_Y));
KC_OAI112_X1 T11387 ( .A(T11369_Y), .B(T11013_Y), .C0(T4439_Y),     .C1(T15872_Y), .Y(T11387_Y));
KC_OAI112_X1 T11363 ( .A(T15900_Y), .B(T4453_Y), .C0(T5815_Y),     .C1(T12800_Y), .Y(T11363_Y));
KC_OAI112_X1 T11553 ( .A(T12212_Y), .B(T4560_Y), .C0(T5149_Y),     .C1(T4514_Y), .Y(T11553_Y));
KC_OAI112_X1 T11605 ( .A(T4597_Y), .B(T6010_Y), .C0(T6019_Y),     .C1(T6010_Y), .Y(T11605_Y));
KC_OAI112_X1 T11995 ( .A(T16112_Y), .B(T12345_Y), .C0(T11624_Y),     .C1(T4688_Y), .Y(T11995_Y));
KC_OAI112_X1 T11784 ( .A(T12360_Y), .B(T12308_Y), .C0(T4733_Y),     .C1(T4700_Y), .Y(T11784_Y));
KC_OAI112_X1 T11758 ( .A(T4749_Y), .B(T6420_Co), .C0(T6420_S),     .C1(T6420_Co), .Y(T11758_Y));
KC_OAI112_X1 T11733 ( .A(T4742_Y), .B(T4738_Y), .C0(T15629_Y),     .C1(T11777_Y), .Y(T11733_Y));
KC_OAI112_X1 T11885 ( .A(T15723_Y), .B(T6680_Y), .C0(T124_Q),     .C1(T14990_Y), .Y(T11885_Y));
KC_OAI112_X1 T11870 ( .A(T6812_Y), .B(T6725_Y), .C0(T896_Y),     .C1(T15032_Y), .Y(T11870_Y));
KC_OAI112_X1 T11868 ( .A(T6811_Y), .B(T6718_Y), .C0(T124_Q),     .C1(T15032_Y), .Y(T11868_Y));
KC_OAI112_X1 T11867 ( .A(T6810_Y), .B(T7272_Y), .C0(T15740_Y),     .C1(T15032_Y), .Y(T11867_Y));
KC_OAI112_X1 T11856 ( .A(T266_Y), .B(T6262_Y), .C0(T6835_Y),     .C1(T10906_Y), .Y(T11856_Y));
KC_OAI112_X1 T11853 ( .A(T7257_Y), .B(T6476_Y), .C0(T9317_Y),     .C1(T11010_Y), .Y(T11853_Y));
KC_OAI112_X1 T11891 ( .A(T15787_Y), .B(T16337_Y), .C0(T8688_Y),     .C1(T10916_Y), .Y(T11891_Y));
KC_OAI112_X1 T11890 ( .A(T15790_Y), .B(T16340_Y), .C0(T8688_Y),     .C1(T14987_Y), .Y(T11890_Y));
KC_OAI112_X1 T11889 ( .A(T15783_Y), .B(T16341_Y), .C0(T8688_Y),     .C1(T14989_Y), .Y(T11889_Y));
KC_OAI112_X1 T11884 ( .A(T15724_Y), .B(T12410_Y), .C0(T15740_Y),     .C1(T14990_Y), .Y(T11884_Y));
KC_OAI112_X1 T11882 ( .A(T15729_Y), .B(T6668_Y), .C0(T14987_Y),     .C1(T6803_Y), .Y(T11882_Y));
KC_OAI112_X1 T11869 ( .A(T12527_Y), .B(T12576_Y), .C0(T5256_Y),     .C1(T13260_Y), .Y(T11869_Y));
KC_OAI112_X1 T11865 ( .A(T6731_Y), .B(T6701_Y), .C0(T9319_Y),     .C1(T15032_Y), .Y(T11865_Y));
KC_OAI112_X1 T11855 ( .A(T520_Y), .B(T6311_Y), .C0(T6835_Y),     .C1(T10884_Y), .Y(T11855_Y));
KC_OAI112_X1 T11852 ( .A(T6345_Y), .B(T492_Y), .C0(T9319_Y),     .C1(T10916_Y), .Y(T11852_Y));
KC_OAI112_X1 T11851 ( .A(T6341_Y), .B(T6336_Y), .C0(T10884_Y),     .C1(T6803_Y), .Y(T11851_Y));
KC_OAI112_X1 T11886 ( .A(T8805_Y), .B(T7646_Y), .C0(T7801_Y),     .C1(T763_Y), .Y(T11886_Y));
KC_OAI112_X1 T11872 ( .A(T9370_Y), .B(T637_Y), .C0(T15747_Y),     .C1(T7839_Y), .Y(T11872_Y));
KC_OAI112_X1 T11859 ( .A(T6733_Y), .B(T11863_Y), .C0(T9308_Y),     .C1(T6690_Y), .Y(T11859_Y));
KC_OAI112_X1 T11854 ( .A(T6253_Y), .B(T6286_Y), .C0(T896_Y),     .C1(T10883_Y), .Y(T11854_Y));
KC_OAI112_X1 T11913 ( .A(T4872_Y), .B(T16274_Y), .C0(T10175_Y),     .C1(T15999_Y), .Y(T11913_Y));
KC_OAI112_X1 T11873 ( .A(T9303_Y), .B(T8725_Y), .C0(T5310_Q),     .C1(T15776_Y), .Y(T11873_Y));
KC_OAI112_X1 T12012 ( .A(T1800_Y), .B(T6370_Y), .C0(T6121_Y),     .C1(T1788_Y), .Y(T12012_Y));
KC_OAI112_X1 T12011 ( .A(T8364_Y), .B(T4915_Y), .C0(T6121_Y),     .C1(T2280_Y), .Y(T12011_Y));
KC_OAI112_X1 T11945 ( .A(T5028_Y), .B(T14941_Q), .C0(T6786_Y),     .C1(T6765_Y), .Y(T11945_Y));
KC_OAI112_X1 T11916 ( .A(T15811_Y), .B(T7983_Y), .C0(T16371_Y),     .C1(T1691_Q), .Y(T11916_Y));
KC_OAI112_X1 T12051 ( .A(T2296_Y), .B(T6817_Y), .C0(T6185_Y),     .C1(T2246_Y), .Y(T12051_Y));
KC_OAI112_X1 T12021 ( .A(T4954_Y), .B(T11550_Y), .C0(T6028_Y),     .C1(T12064_Y), .Y(T12021_Y));
KC_OAI112_X1 T12020 ( .A(T2216_Y), .B(T11549_Y), .C0(T2279_Y),     .C1(T12064_Y), .Y(T12020_Y));
KC_OAI112_X1 T12010 ( .A(T5555_Y), .B(T2251_Y), .C0(T16041_Y),     .C1(T6000_Y), .Y(T12010_Y));
KC_OAI112_X1 T11949 ( .A(T2041_Y), .B(T2060_Y), .C0(T10519_Y),     .C1(T16367_Y), .Y(T11949_Y));
KC_OAI112_X1 T11937 ( .A(T5028_Y), .B(T14937_Q), .C0(T15685_Y),     .C1(T6765_Y), .Y(T11937_Y));
KC_OAI112_X1 T11936 ( .A(T11934_Y), .B(T10479_Y), .C0(T6781_Y),     .C1(T15398_Y), .Y(T11936_Y));
KC_OAI112_X1 T11935 ( .A(T5028_Y), .B(T14938_Q), .C0(T6781_Y),     .C1(T6765_Y), .Y(T11935_Y));
KC_OAI112_X1 T11934 ( .A(T5028_Y), .B(T14934_Q), .C0(T15684_Y),     .C1(T2448_Y), .Y(T11934_Y));
KC_OAI112_X1 T11933 ( .A(T11954_Y), .B(T10480_Y), .C0(T15685_Y),     .C1(T15398_Y), .Y(T11933_Y));
KC_OAI112_X1 T11926 ( .A(T11112_Y), .B(T9643_Y), .C0(T6460_Y),     .C1(T6592_Y), .Y(T11926_Y));
KC_OAI112_X1 T16263 ( .A(T2593_Y), .B(T2596_Y), .C0(T2620_Y),     .C1(T4864_Y), .Y(T16263_Y));
KC_OAI112_X1 T12060 ( .A(T6831_Y), .B(T12973_Y), .C0(T6581_Y),     .C1(T2882_Y), .Y(T12060_Y));
KC_OAI112_X1 T11929 ( .A(T11931_Y), .B(T10473_Y), .C0(T632_Y),     .C1(T6592_Y), .Y(T11929_Y));
KC_OAI112_X1 T11928 ( .A(T2457_Y), .B(T2449_Y), .C0(T2464_Y),     .C1(T2458_Y), .Y(T11928_Y));
KC_OAI112_X1 T11927 ( .A(T5028_Y), .B(T14839_Q), .C0(T6773_Y),     .C1(T6765_Y), .Y(T11927_Y));
KC_OAI112_X1 T12057 ( .A(T5047_Y), .B(T11807_Y), .C0(T3439_Y),     .C1(T6039_Y), .Y(T12057_Y));
KC_OAI112_X1 T12056 ( .A(T12365_Y), .B(T11722_Y), .C0(T3467_Y),     .C1(T12250_Y), .Y(T12056_Y));
KC_OAI112_X1 T12041 ( .A(T3419_Y), .B(T5050_Y), .C0(T10979_Y),     .C1(T11677_Y), .Y(T12041_Y));
KC_OAI112_X1 T12040 ( .A(T11676_Y), .B(T12358_Y), .C0(T3383_Y),     .C1(T11764_Y), .Y(T12040_Y));
KC_OAI112_X1 T11997 ( .A(T5525_Q), .B(T3413_Y), .C0(T11604_Y),     .C1(T11641_Y), .Y(T11997_Y));
KC_OAI112_X1 T12054 ( .A(T12362_Y), .B(T4133_Y), .C0(T4062_Y),     .C1(T3368_Y), .Y(T12054_Y));
KC_OAI112_X1 T12019 ( .A(T15704_Y), .B(T10944_Y), .C0(T10958_Y),     .C1(T11577_Y), .Y(T12019_Y));
KC_OAI112_X1 T12018 ( .A(T11617_Y), .B(T8478_Y), .C0(T3975_Y),     .C1(T4569_Y), .Y(T12018_Y));
KC_OAI112_X1 T11979 ( .A(T8451_Y), .B(T12341_Y), .C0(T5756_Y),     .C1(T3827_Y), .Y(T11979_Y));
KC_OAI112_X1 T11978 ( .A(T3847_Y), .B(T12157_Y), .C0(T3856_Y),     .C1(T5103_Y), .Y(T11978_Y));
KC_OAI112_X1 T11965 ( .A(T15908_Y), .B(T4486_Y), .C0(T15697_Y),     .C1(T15907_Y), .Y(T11965_Y));
KC_OAI112_X1 T11066 ( .A(T6949_Y), .B(T6938_Y), .C0(T6819_Y),     .C1(T10883_Y), .Y(T11066_Y));
KC_OAI112_X1 T11055 ( .A(T6964_Y), .B(T218_Y), .C0(T9318_Y),     .C1(T10906_Y), .Y(T11055_Y));
KC_OAI112_X1 T11925 ( .A(T11110_Y), .B(T10440_Y), .C0(T6459_Y),     .C1(T6592_Y), .Y(T11925_Y));
KC_OAI112_X1 T11849 ( .A(T6343_Y), .B(T6337_Y), .C0(T11016_Y),     .C1(T6803_Y), .Y(T11849_Y));
KC_OAI112_X1 T6755 ( .A(T11938_Y), .B(T10485_Y), .C0(T417_Y),     .C1(T15398_Y), .Y(T6755_Y));
KC_OAI112_X1 T11955 ( .A(T11951_Y), .B(T10476_Y), .C0(T15684_Y),     .C1(T6592_Y), .Y(T11955_Y));
KC_OAI112_X1 T11904 ( .A(T6739_Y), .B(T11907_Y), .C0(T9307_Y),     .C1(T5702_Y), .Y(T11904_Y));
KC_OAI112_X1 T11135 ( .A(T11136_Y), .B(T9688_Y), .C0(T410_Y),     .C1(T15398_Y), .Y(T11135_Y));
KC_OAI112_X1 T11132 ( .A(T11113_Y), .B(T9674_Y), .C0(T488_Y),     .C1(T6592_Y), .Y(T11132_Y));
KC_OAI112_X1 T11129 ( .A(T11117_Y), .B(T9647_Y), .C0(T15401_Y),     .C1(T15398_Y), .Y(T11129_Y));
KC_OAI112_X1 T11116 ( .A(T11125_Y), .B(T9673_Y), .C0(T6764_Y),     .C1(T15398_Y), .Y(T11116_Y));
KC_OAI112_X1 T11114 ( .A(T2449_Y), .B(T13655_Q), .C0(T6459_Y),     .C1(T2448_Y), .Y(T11114_Y));
KC_OAI112_X1 T11942 ( .A(T11930_Y), .B(T9756_Y), .C0(T6773_Y),     .C1(T15398_Y), .Y(T11942_Y));
KC_OAI112_X1 T11166 ( .A(T15730_Y), .B(T7446_Y), .C0(T6835_Y),     .C1(T14990_Y), .Y(T11166_Y));
KC_OAI112_X1 T11152 ( .A(T7392_Y), .B(T7391_Y), .C0(T15032_Y),     .C1(T6803_Y), .Y(T11152_Y));
KC_OAI112_X1 T11150 ( .A(T7388_Y), .B(T7387_Y), .C0(T896_Y),     .C1(T14987_Y), .Y(T11150_Y));
KC_OAI112_X1 T11189 ( .A(T8707_Y), .B(T8725_Y), .C0(T5561_Q),     .C1(T15773_Y), .Y(T11189_Y));
KC_OAI112_X1 T11259 ( .A(T2014_Y), .B(T5366_Q), .C0(T1162_Y),     .C1(T1123_Y), .Y(T11259_Y));
KC_OAI112_X1 T11285 ( .A(T10056_Y), .B(T2036_Y), .C0(T1518_Y),     .C1(T10078_Y), .Y(T11285_Y));
KC_OAI112_X1 T11302 ( .A(T9132_Y), .B(T415_Y), .C0(T9182_Y),     .C1(T9150_Y), .Y(T11302_Y));
KC_OAI112_X1 T11973 ( .A(T5778_Y), .B(T3795_Y), .C0(T8184_Y),     .C1(T4436_Y), .Y(T11973_Y));
KC_OAI112_X1 T11328 ( .A(T3803_Y), .B(T3800_Y), .C0(T4388_Y),     .C1(T5760_Y), .Y(T11328_Y));
KC_OAI112_X1 T11326 ( .A(T12135_Y), .B(T12334_Y), .C0(T5774_Y),     .C1(T12140_Y), .Y(T11326_Y));
KC_OAI112_X1 T11403 ( .A(T3835_Y), .B(T10898_Y), .C0(T3855_Y),     .C1(T14543_Q), .Y(T11403_Y));
KC_OAI112_X1 T11469 ( .A(T3920_Y), .B(T3858_Y), .C0(T5870_Y),     .C1(T4471_Y), .Y(T11469_Y));
KC_OAI112_X1 T11447 ( .A(T3864_Y), .B(T6228_Y), .C0(T5874_Y),     .C1(T4471_Y), .Y(T11447_Y));
KC_OAI112_X1 T11439 ( .A(T5107_Y), .B(T11440_Y), .C0(T3849_Y),     .C1(T3800_Y), .Y(T11439_Y));
KC_OAI112_X1 T11623 ( .A(T12245_Y), .B(T2271_Y), .C0(T15611_Y),     .C1(T6000_Y), .Y(T11623_Y));
KC_OAI112_X1 T11612 ( .A(T2223_Y), .B(T2271_Y), .C0(T2246_Y),     .C1(T6000_Y), .Y(T11612_Y));
KC_OAI112_X1 T11719 ( .A(T10623_Y), .B(T12042_Y), .C0(T2879_Y),     .C1(T5523_Y), .Y(T11719_Y));
KC_OAI112_X1 T11700 ( .A(T6466_Y), .B(T1812_Y), .C0(T1804_Y),     .C1(T6184_Y), .Y(T11700_Y));
KC_OAI112_X1 T11692 ( .A(T2273_Y), .B(T1819_Y), .C0(T6125_Y),     .C1(T6121_Y), .Y(T11692_Y));
KC_OAI112_X1 T11734 ( .A(T4143_Y), .B(T11684_Y), .C0(T3481_Y),     .C1(T8403_Y), .Y(T11734_Y));
KC_OAI112_X1 T11841 ( .A(T5534_Y), .B(T10993_Y), .C0(T12864_Y),     .C1(T2865_Y), .Y(T11841_Y));
KC_OAI112_X1 T11838 ( .A(T11775_Y), .B(T6541_Y), .C0(T11772_Y),     .C1(T1856_Q), .Y(T11838_Y));
KC_OAI112_X1 T12036 ( .A(T3383_Y), .B(T3382_Y), .C0(T5056_Y),     .C1(T3409_Y), .Y(T12036_Y));
KC_OAI112_X1 T11944 ( .A(T6754_Y), .B(T10483_Y), .C0(T629_Y),     .C1(T15398_Y), .Y(T11944_Y));
KC_OAI112_X1 T11881 ( .A(T7451_Y), .B(T6661_Y), .C0(T6803_Y),     .C1(T14990_Y), .Y(T11881_Y));
KC_BUF_X6 T5608 ( .Y(T5608_Y), .A(T58_Y));
KC_BUF_X6 T7074 ( .Y(T7074_Y), .A(T869_Y));
KC_BUF_X6 T7073 ( .Y(T7073_Y), .A(T869_Y));
KC_BUF_X6 T7609 ( .Y(T7609_Y), .A(T7668_Y));
KC_BUF_X6 T7919 ( .Y(T7919_Y), .A(T16278_Y));
KC_BUF_X6 T1428 ( .Y(T1428_Y), .A(T11296_Y));
KC_BUF_X6 T8106 ( .Y(T8106_Y), .A(T8091_Y));
KC_BUF_X6 T1602 ( .Y(T1602_Y), .A(T9136_Y));
KC_BUF_X6 T5299 ( .Y(T5299_Y), .A(T16281_Y));
KC_BUF_X6 T34 ( .Y(T34_Y), .A(T271_Y));
KC_BUF_X6 T7108 ( .Y(T7108_Y), .A(T11209_Y));
KC_BUF_X6 T7318 ( .Y(T7318_Y), .A(T8723_Y));
KC_BUF_X6 T15722 ( .Y(T15722_Y), .A(T8836_Y));
KC_BUF_X6 T7385 ( .Y(T7385_Y), .A(T7950_Y));
KC_BUF_X6 T7675 ( .Y(T7675_Y), .A(T869_Y));
KC_BUF_X6 T7607 ( .Y(T7607_Y), .A(T11237_Y));
KC_BUF_X6 T6350 ( .Y(T6350_Y), .A(T8739_Y));
KC_BUF_X6 T7668 ( .Y(T7668_Y), .A(T15230_Y));
KC_BUF_X6 T7623 ( .Y(T7623_Y), .A(T8696_Y));
KC_BUF_X6 T7603 ( .Y(T7603_Y), .A(T8861_Y));
KC_BUF_X6 T7899 ( .Y(T7899_Y), .A(T16419_Y));
KC_BUF_X6 T7859 ( .Y(T7859_Y), .A(T8835_Y));
KC_BUF_X6 T7854 ( .Y(T7854_Y), .A(T16428_Y));
KC_BUF_X6 T7853 ( .Y(T7853_Y), .A(T8809_Y));
KC_BUF_X6 T7815 ( .Y(T7815_Y), .A(T16430_Y));
KC_BUF_X6 T7811 ( .Y(T7811_Y), .A(T5108_Y));
KC_BUF_X6 T7810 ( .Y(T7810_Y), .A(T8833_Y));
KC_BUF_X6 T7809 ( .Y(T7809_Y), .A(T5143_Y));
KC_BUF_X6 T7243 ( .Y(T7243_Y), .A(T7668_Y));
KC_BUF_X6 T7242 ( .Y(T7242_Y), .A(T7668_Y));
KC_BUF_X6 T7364 ( .Y(T7364_Y), .A(T12610_Y));
KC_BUF_X6 T7845 ( .Y(T7845_Y), .A(T14991_Y));
KC_BUF_X6 T7088 ( .Y(T7088_Y), .A(T9359_Y));
KC_BUF_X6 T8030 ( .Y(T8030_Y), .A(T1244_Y));
KC_BUF_X6 T16278 ( .Y(T16278_Y), .A(T9435_Y));
KC_BUF_X6 T10535 ( .Y(T10535_Y), .A(T1244_Y));
KC_BUF_X6 T7798 ( .Y(T7798_Y), .A(T1244_Y));
KC_BUF_X6 T7797 ( .Y(T7797_Y), .A(T1244_Y));
KC_BUF_X6 T7740 ( .Y(T7740_Y), .A(T1244_Y));
KC_BUF_X6 T10661 ( .Y(T10661_Y), .A(T1244_Y));
KC_BUF_X6 T10727 ( .Y(T10727_Y), .A(T1244_Y));
KC_BUF_X6 T10697 ( .Y(T10697_Y), .A(T1244_Y));
KC_BUF_X6 T1276 ( .Y(T1276_Y), .A(T12771_Y));
KC_BUF_X6 T7337 ( .Y(T7337_Y), .A(T16063_Y));
KC_BUF_X6 T7707 ( .Y(T7707_Y), .A(T16449_Y));
KC_BUF_X6 T6894 ( .Y(T6894_Y), .A(T9520_Y));
KC_BUF_X6 T7323 ( .Y(T7323_Y), .A(T16063_Y));
KC_BUF_X6 T7780 ( .Y(T7780_Y), .A(T12535_Y));
KC_BUF_X6 T7703 ( .Y(T7703_Y), .A(T16448_Y));
KC_BUF_X6 T10743 ( .Y(T10743_Y), .A(T8001_Y));
KC_BUF_X6 T8011 ( .Y(T8011_Y), .A(T16063_Y));
KC_BUF_X6 T8000 ( .Y(T8000_Y), .A(T2027_Y));
KC_BUF_X6 T7986 ( .Y(T7986_Y), .A(T10883_Y));
KC_BUF_X6 T7952 ( .Y(T7952_Y), .A(T16245_Y));
KC_BUF_X6 T1738 ( .Y(T1738_Y), .A(T5042_Y));
KC_BUF_X6 T6737 ( .Y(T6737_Y), .A(T16456_Y));
KC_BUF_X6 T1825 ( .Y(T1825_Y), .A(T11482_Y));
KC_BUF_X6 T1998 ( .Y(T1998_Y), .A(T4932_Q));
KC_BUF_X6 T2000 ( .Y(T2000_Y), .A(T1244_Y));
KC_BUF_X6 T2042 ( .Y(T2042_Y), .A(T2583_Q));
KC_BUF_X6 T2062 ( .Y(T2062_Y), .A(T1244_Y));
KC_BUF_X6 T2063 ( .Y(T2063_Y), .A(T1244_Y));
KC_BUF_X6 T2073 ( .Y(T2073_Y), .A(T15802_Q));
KC_BUF_X6 T2098 ( .Y(T2098_Y), .A(T15895_Y));
KC_BUF_X6 T2099 ( .Y(T2099_Y), .A(T13302_Y));
KC_BUF_X6 T2109 ( .Y(T2109_Y), .A(T2761_Y));
KC_BUF_X6 T2133 ( .Y(T2133_Y), .A(T12462_Y));
KC_BUF_X6 T2148 ( .Y(T2148_Y), .A(T2765_Y));
KC_BUF_X6 T2169 ( .Y(T2169_Y), .A(T2081_Y));
KC_BUF_X6 T2317 ( .Y(T2317_Y), .A(T8388_Y));
KC_BUF_X6 T2322 ( .Y(T2322_Y), .A(T2081_Y));
KC_BUF_X6 T2331 ( .Y(T2331_Y), .A(T11783_Y));
KC_BUF_X6 T2341 ( .Y(T2341_Y), .A(T8309_Y));
KC_BUF_X6 T2367 ( .Y(T2367_Y), .A(T2388_Q));
KC_BUF_X6 T2368 ( .Y(T2368_Y), .A(T12879_Y));
KC_BUF_X6 T2369 ( .Y(T2369_Y), .A(T11840_Y));
KC_BUF_X6 T2474 ( .Y(T2474_Y), .A(T10195_Y));
KC_BUF_X6 T2475 ( .Y(T2475_Y), .A(T10195_Y));
KC_BUF_X6 T2522 ( .Y(T2522_Y), .A(T1244_Y));
KC_BUF_X6 T2564 ( .Y(T2564_Y), .A(T16164_Y));
KC_BUF_X6 T2565 ( .Y(T2565_Y), .A(T9957_Y));
KC_BUF_X6 T2566 ( .Y(T2566_Y), .A(T10195_Y));
KC_BUF_X6 T2658 ( .Y(T2658_Y), .A(T4381_Q));
KC_BUF_X6 T2706 ( .Y(T2706_Y), .A(T12463_Y));
KC_BUF_X6 T2734 ( .Y(T2734_Y), .A(T3963_Y));
KC_BUF_X6 T2757 ( .Y(T2757_Y), .A(T16006_Y));
KC_BUF_X6 T2782 ( .Y(T2782_Y), .A(T3451_Y));
KC_BUF_X6 T2830 ( .Y(T2830_Y), .A(T12006_Y));
KC_BUF_X6 T2854 ( .Y(T2854_Y), .A(T2838_Y));
KC_BUF_X6 T2865 ( .Y(T2865_Y), .A(T2838_Y));
KC_BUF_X6 T2933 ( .Y(T2933_Y), .A(T5517_Y));
KC_BUF_X6 T3070 ( .Y(T3070_Y), .A(T422_Y));
KC_BUF_X6 T3071 ( .Y(T3071_Y), .A(T3781_Y));
KC_BUF_X6 T3072 ( .Y(T3072_Y), .A(T3780_Y));
KC_BUF_X6 T3073 ( .Y(T3073_Y), .A(T16448_Y));
KC_BUF_X6 T3222 ( .Y(T3222_Y), .A(T2668_Y));
KC_BUF_X6 T3250 ( .Y(T3250_Y), .A(T4410_Y));
KC_BUF_X6 T3252 ( .Y(T3252_Y), .A(T13055_Y));
KC_BUF_X6 T3288 ( .Y(T3288_Y), .A(T3331_Y));
KC_BUF_X6 T3292 ( .Y(T3292_Y), .A(T15981_Y));
KC_BUF_X6 T3294 ( .Y(T3294_Y), .A(T4532_Y));
KC_BUF_X6 T3295 ( .Y(T3295_Y), .A(T10641_Y));
KC_BUF_X6 T3296 ( .Y(T3296_Y), .A(T3329_Y));
KC_BUF_X6 T3298 ( .Y(T3298_Y), .A(T11477_Y));
KC_BUF_X6 T3299 ( .Y(T3299_Y), .A(T5061_Y));
KC_BUF_X6 T3322 ( .Y(T3322_Y), .A(T3318_Y));
KC_BUF_X6 T3323 ( .Y(T3323_Y), .A(T16503_Y));
KC_BUF_X6 T3324 ( .Y(T3324_Y), .A(T12461_Y));
KC_BUF_X6 T3326 ( .Y(T3326_Y), .A(T16202_Y));
KC_BUF_X6 T3327 ( .Y(T3327_Y), .A(T4411_Y));
KC_BUF_X6 T3347 ( .Y(T3347_Y), .A(T15912_Y));
KC_BUF_X6 T3351 ( .Y(T3351_Y), .A(T3268_Y));
KC_BUF_X6 T3358 ( .Y(T3358_Y), .A(T4028_Y));
KC_BUF_X6 T3359 ( .Y(T3359_Y), .A(T2239_Y));
KC_BUF_X6 T3425 ( .Y(T3425_Y), .A(T12244_Y));
KC_BUF_X6 T3610 ( .Y(T3610_Y), .A(T2027_Y));
KC_BUF_X6 T3635 ( .Y(T3635_Y), .A(T2027_Y));
KC_BUF_X6 T3650 ( .Y(T3650_Y), .A(T3774_Y));
KC_BUF_X6 T3653 ( .Y(T3653_Y), .A(T3775_Y));
KC_BUF_X6 T3707 ( .Y(T3707_Y), .A(T3706_Y));
KC_BUF_X6 T3728 ( .Y(T3728_Y), .A(T12785_Y));
KC_BUF_X6 T3830 ( .Y(T3830_Y), .A(T15864_Y));
KC_BUF_X6 T3868 ( .Y(T3868_Y), .A(T3883_Q));
KC_BUF_X6 T3904 ( .Y(T3904_Y), .A(T8263_Y));
KC_BUF_X6 T3940 ( .Y(T3940_Y), .A(T3334_Y));
KC_BUF_X6 T3942 ( .Y(T3942_Y), .A(T12214_Y));
KC_BUF_X6 T3950 ( .Y(T3950_Y), .A(T5963_Y));
KC_BUF_X6 T3982 ( .Y(T3982_Y), .A(T13150_Q));
KC_BUF_X6 T4037 ( .Y(T4037_Y), .A(T5111_Y));
KC_BUF_X6 T4071 ( .Y(T4071_Y), .A(T11558_Y));
KC_BUF_X6 T4151 ( .Y(T4151_Y), .A(T12842_Y));
KC_BUF_X6 T4156 ( .Y(T4156_Y), .A(T4019_Y));
KC_BUF_X6 T4272 ( .Y(T4272_Y), .A(T9852_Y));
KC_BUF_X6 T4386 ( .Y(T4386_Y), .A(T5044_Y));
KC_BUF_X6 T4402 ( .Y(T4402_Y), .A(T2709_Y));
KC_BUF_X6 T4447 ( .Y(T4447_Y), .A(T10914_Y));
KC_BUF_X6 T4470 ( .Y(T4470_Y), .A(T10228_Y));
KC_BUF_X6 T4479 ( .Y(T4479_Y), .A(T4435_Y));
KC_BUF_X6 T4594 ( .Y(T4594_Y), .A(T12244_Y));
KC_BUF_X6 T4638 ( .Y(T4638_Y), .A(T241_Y));
KC_BUF_X6 T4661 ( .Y(T4661_Y), .A(T12463_Y));
KC_BUF_X6 T4697 ( .Y(T4697_Y), .A(T4637_Y));
KC_BUF_X6 T4741 ( .Y(T4741_Y), .A(T4754_Y));
KC_BUF_X6 T4761 ( .Y(T4761_Y), .A(T5511_Q));
KC_BUF_X6 T15721 ( .Y(T15721_Y), .A(T7668_Y));
KC_BUF_X6 T15731 ( .Y(T15731_Y), .A(T11210_Y));
KC_BUF_X6 T10788 ( .Y(T10788_Y), .A(T16063_Y));
KC_BUF_X6 T4937 ( .Y(T4937_Y), .A(T9642_Y));
KC_BUF_X6 T4963 ( .Y(T4963_Y), .A(T8428_Y));
KC_BUF_X6 T4983 ( .Y(T4983_Y), .A(T10509_Y));
KC_BUF_X6 T4997 ( .Y(T4997_Y), .A(T2652_Y));
KC_BUF_X6 T5009 ( .Y(T5009_Y), .A(T12220_Y));
KC_BUF_X6 T5040 ( .Y(T5040_Y), .A(T5077_Y));
KC_BUF_X6 T5088 ( .Y(T5088_Y), .A(T16063_Y));
KC_BUF_X6 T5141 ( .Y(T5141_Y), .A(T4517_Y));
KC_BUF_X6 T5142 ( .Y(T5142_Y), .A(T4554_Y));
KC_BUF_X6 T7606 ( .Y(T7606_Y), .A(T8837_Y));
KC_BUF_X6 T16382 ( .Y(T16382_Y), .A(T8814_Y));
KC_BUF_X6 T5331 ( .Y(T5331_Y), .A(T3779_Y));
KC_BUF_X6 T5444 ( .Y(T5444_Y), .A(T3963_Y));
KC_BUF_X6 T5504 ( .Y(T5504_Y), .A(T1708_Y));
KC_BUF_X6 T10757 ( .Y(T10757_Y), .A(T15467_Y));
KC_AND2_X2 T8538 ( .B(T8537_Y), .A(T8543_Y), .Y(T8538_Y));
KC_AND2_X2 T9297 ( .B(T878_Y), .A(T6913_Y), .Y(T9297_Y));
KC_AND2_X2 T8960 ( .B(T8089_Y), .A(T8993_Co), .Y(T8960_Y));
KC_AND2_X2 T9123 ( .B(T15093_Y), .A(T15109_Y), .Y(T9123_Y));
KC_AND2_X2 T9072 ( .B(T2390_Y), .A(T15109_Y), .Y(T9072_Y));
KC_AND2_X2 T9071 ( .B(T9118_Y), .A(T9117_Y), .Y(T9071_Y));
KC_AND2_X2 T8983 ( .B(T1594_Y), .A(T7872_Y), .Y(T8983_Y));
KC_AND2_X2 T8903 ( .B(T1199_Y), .A(T756_Y), .Y(T8903_Y));
KC_AND2_X2 T9109 ( .B(T605_Q), .A(T598_Y), .Y(T9109_Y));
KC_AND2_X2 T9293 ( .B(T110_Y), .A(T826_Q), .Y(T9293_Y));
KC_AND2_X2 T8585 ( .B(T245_Y), .A(T820_Q), .Y(T8585_Y));
KC_AND2_X2 T8571 ( .B(T301_Y), .A(T823_Q), .Y(T8571_Y));
KC_AND2_X2 T8566 ( .B(T244_Y), .A(T815_Q), .Y(T8566_Y));
KC_AND2_X2 T9263 ( .B(T315_Y), .A(T848_Q), .Y(T9263_Y));
KC_AND2_X2 T8618 ( .B(T334_Y), .A(T838_Q), .Y(T8618_Y));
KC_AND2_X2 T9417 ( .B(T15485_Y), .A(T15660_Y), .Y(T9417_Y));
KC_AND2_X2 T8857 ( .B(T15485_Y), .A(T975_Y), .Y(T8857_Y));
KC_AND2_X2 T8856 ( .B(T15485_Y), .A(T15463_Y), .Y(T8856_Y));
KC_AND2_X2 T8806 ( .B(T15485_Y), .A(T1059_Y), .Y(T8806_Y));
KC_AND2_X2 T9140 ( .B(T977_Q), .A(T1001_Q), .Y(T9140_Y));
KC_AND2_X2 T9034 ( .B(T972_Y), .A(T9033_Y), .Y(T9034_Y));
KC_AND2_X2 T8634 ( .B(T317_Y), .A(T834_Q), .Y(T8634_Y));
KC_AND2_X2 T9506 ( .B(T6373_Y), .A(T15781_Y), .Y(T9506_Y));
KC_AND2_X2 T9505 ( .B(T6374_Y), .A(T15772_Y), .Y(T9505_Y));
KC_AND2_X2 T9504 ( .B(T6372_Y), .A(T15780_Y), .Y(T9504_Y));
KC_AND2_X2 T8719 ( .B(T5804_Y), .A(T16090_Y), .Y(T8719_Y));
KC_AND2_X2 T9413 ( .B(T15485_Y), .A(T1709_Y), .Y(T9413_Y));
KC_AND2_X2 T8858 ( .B(T15485_Y), .A(T1578_Y), .Y(T8858_Y));
KC_AND2_X2 T8848 ( .B(T15458_Y), .A(T949_Q), .Y(T8848_Y));
KC_AND2_X2 T8832 ( .B(T8794_Y), .A(T9402_Y), .Y(T8832_Y));
KC_AND2_X2 T8772 ( .B(T903_Y), .A(T1249_Q), .Y(T8772_Y));
KC_AND2_X2 T8764 ( .B(T5376_Q), .A(T8938_Y), .Y(T8764_Y));
KC_AND2_X2 T9002 ( .B(T972_Y), .A(T9431_Y), .Y(T9002_Y));
KC_AND2_X2 T8976 ( .B(T9056_Y), .A(T5386_Q), .Y(T8976_Y));
KC_AND2_X2 T9463 ( .B(T977_Q), .A(T998_Q), .Y(T9463_Y));
KC_AND2_X2 T9033 ( .B(T10298_Y), .A(T9031_Y), .Y(T9033_Y));
KC_AND2_X2 T9507 ( .B(T6220_Y), .A(T15778_Y), .Y(T9507_Y));
KC_AND2_X2 T9503 ( .B(T5782_Y), .A(T15774_Y), .Y(T9503_Y));
KC_AND2_X2 T9714 ( .B(T2391_Y), .A(T12706_Y), .Y(T9714_Y));
KC_AND2_X2 T8657 ( .B(T498_Y), .A(T8656_Y), .Y(T8657_Y));
KC_AND2_X2 T9816 ( .B(T7845_Y), .A(T7385_Y), .Y(T9816_Y));
KC_AND2_X2 T8728 ( .B(T715_Y), .A(T12690_Y), .Y(T8728_Y));
KC_AND2_X2 T10330 ( .B(T7845_Y), .A(T15722_Y), .Y(T10330_Y));
KC_AND2_X2 T9918 ( .B(T16422_Q), .A(T1095_Q), .Y(T9918_Y));
KC_AND2_X2 T9985 ( .B(T15485_Y), .A(T1450_Y), .Y(T9985_Y));
KC_AND2_X2 T10168 ( .B(T15485_Y), .A(T16271_Y), .Y(T10168_Y));
KC_AND2_X2 T10167 ( .B(T15485_Y), .A(T1456_Y), .Y(T10167_Y));
KC_AND2_X2 T10166 ( .B(T15485_Y), .A(T15531_Y), .Y(T10166_Y));
KC_AND2_X2 T10165 ( .B(T972_Y), .A(T1472_Y), .Y(T10165_Y));
KC_AND2_X2 T10164 ( .B(T15485_Y), .A(T1058_Y), .Y(T10164_Y));
KC_AND2_X2 T9982 ( .B(T10163_Y), .A(T10293_Y), .Y(T9982_Y));
KC_AND2_X2 T10157 ( .B(T4902_Y), .A(T1365_Y), .Y(T10157_Y));
KC_AND2_X2 T9608 ( .B(T12529_Y), .A(T1431_Y), .Y(T9608_Y));
KC_AND2_X2 T9696 ( .B(T12583_Y), .A(T4885_Y), .Y(T9696_Y));
KC_AND2_X2 T9812 ( .B(T12639_Y), .A(T4885_Y), .Y(T9812_Y));
KC_AND2_X2 T9811 ( .B(T12640_Y), .A(T4885_Y), .Y(T9811_Y));
KC_AND2_X2 T9803 ( .B(T12629_Y), .A(T4885_Y), .Y(T9803_Y));
KC_AND2_X2 T9793 ( .B(T12626_Y), .A(T4885_Y), .Y(T9793_Y));
KC_AND2_X2 T9792 ( .B(T12625_Y), .A(T4885_Y), .Y(T9792_Y));
KC_AND2_X2 T9789 ( .B(T12624_Y), .A(T4885_Y), .Y(T9789_Y));
KC_AND2_X2 T9788 ( .B(T12627_Y), .A(T4885_Y), .Y(T9788_Y));
KC_AND2_X2 T10325 ( .B(T12899_Y), .A(T1491_Y), .Y(T10325_Y));
KC_AND2_X2 T10324 ( .B(T12897_Y), .A(T1491_Y), .Y(T10324_Y));
KC_AND2_X2 T9913 ( .B(T12688_Y), .A(T1491_Y), .Y(T9913_Y));
KC_AND2_X2 T9912 ( .B(T12687_Y), .A(T1491_Y), .Y(T9912_Y));
KC_AND2_X2 T9911 ( .B(T12686_Y), .A(T1491_Y), .Y(T9911_Y));
KC_AND2_X2 T9910 ( .B(T12680_Y), .A(T1491_Y), .Y(T9910_Y));
KC_AND2_X2 T9888 ( .B(T12689_Y), .A(T1491_Y), .Y(T9888_Y));
KC_AND2_X2 T10207 ( .B(T10005_Y), .A(T2073_Y), .Y(T10207_Y));
KC_AND2_X2 T10417 ( .B(T6750_Y), .A(T4885_Y), .Y(T10417_Y));
KC_AND2_X2 T10416 ( .B(T12922_Y), .A(T4885_Y), .Y(T10416_Y));
KC_AND2_X2 T9700 ( .B(T12600_Y), .A(T1453_Y), .Y(T9700_Y));
KC_AND2_X2 T9699 ( .B(T12596_Y), .A(T1453_Y), .Y(T9699_Y));
KC_AND2_X2 T9698 ( .B(T12599_Y), .A(T1453_Y), .Y(T9698_Y));
KC_AND2_X2 T9907 ( .B(T12679_Y), .A(T1491_Y), .Y(T9907_Y));
KC_AND2_X2 T9906 ( .B(T12894_Y), .A(T1491_Y), .Y(T9906_Y));
KC_AND2_X2 T9905 ( .B(T12684_Y), .A(T1491_Y), .Y(T9905_Y));
KC_AND2_X2 T9903 ( .B(T12683_Y), .A(T1491_Y), .Y(T9903_Y));
KC_AND2_X2 T10225 ( .B(T10003_Y), .A(T2073_Y), .Y(T10225_Y));
KC_AND2_X2 T9808 ( .B(T12937_Y), .A(T1492_Y), .Y(T9808_Y));
KC_AND2_X2 T9782 ( .B(T7780_Y), .A(T15662_Y), .Y(T9782_Y));
KC_AND2_X2 T9904 ( .B(T12682_Y), .A(T1491_Y), .Y(T9904_Y));
KC_AND2_X2 T10224 ( .B(T9981_Y), .A(T2073_Y), .Y(T10224_Y));
KC_AND2_X2 T10445 ( .B(T12551_Y), .A(T2452_Y), .Y(T10445_Y));
KC_AND2_X2 T9687 ( .B(T12572_Y), .A(T1930_Y), .Y(T9687_Y));
KC_AND2_X2 T9618 ( .B(T12540_Y), .A(T1930_Y), .Y(T9618_Y));
KC_AND2_X2 T9617 ( .B(T12532_Y), .A(T1930_Y), .Y(T9617_Y));
KC_AND2_X2 T9609 ( .B(T12534_Y), .A(T1930_Y), .Y(T9609_Y));
KC_AND2_X2 T9606 ( .B(T12533_Y), .A(T1930_Y), .Y(T9606_Y));
KC_AND2_X2 T9605 ( .B(T12528_Y), .A(T1930_Y), .Y(T9605_Y));
KC_AND2_X2 T8420 ( .B(T15515_Y), .A(T6216_Y), .Y(T8420_Y));
KC_AND2_X2 T10443 ( .B(T12570_Y), .A(T2452_Y), .Y(T10443_Y));
KC_AND2_X2 T9601 ( .B(T12569_Y), .A(T2452_Y), .Y(T9601_Y));
KC_AND2_X2 T8533 ( .B(T12949_Y), .A(T1930_Y), .Y(T8533_Y));
KC_AND2_X2 T9760 ( .B(T12593_Y), .A(T1930_Y), .Y(T9760_Y));
KC_AND2_X2 T9759 ( .B(T12935_Y), .A(T1930_Y), .Y(T9759_Y));
KC_AND2_X2 T9758 ( .B(T12554_Y), .A(T1930_Y), .Y(T9758_Y));
KC_AND2_X2 T9757 ( .B(T12597_Y), .A(T1930_Y), .Y(T9757_Y));
KC_AND2_X2 T9749 ( .B(T12594_Y), .A(T1930_Y), .Y(T9749_Y));
KC_AND2_X2 T10083 ( .B(T2057_Y), .A(T15003_Y), .Y(T10083_Y));
KC_AND2_X2 T10065 ( .B(T5906_Y), .A(T10100_Y), .Y(T10065_Y));
KC_AND2_X2 T10062 ( .B(T15506_Y), .A(T9974_Y), .Y(T10062_Y));
KC_AND2_X2 T10205 ( .B(T5731_Y), .A(T2717_Y), .Y(T10205_Y));
KC_AND2_X2 T10185 ( .B(T16237_Y), .A(T16234_Y), .Y(T10185_Y));
KC_AND2_X2 T8423 ( .B(T2347_Y), .A(T12316_Y), .Y(T8423_Y));
KC_AND2_X2 T8418 ( .B(T12313_Y), .A(T15140_Y), .Y(T8418_Y));
KC_AND2_X2 T8410 ( .B(T11770_Y), .A(T2331_Y), .Y(T8410_Y));
KC_AND2_X2 T8433 ( .B(T2951_Y), .A(T2956_Y), .Y(T8433_Y));
KC_AND2_X2 T8432 ( .B(T8433_Y), .A(T8433_Y), .Y(T8432_Y));
KC_AND2_X2 T8156 ( .B(T4979_Y), .A(T6605_Y), .Y(T8156_Y));
KC_AND2_X2 T10456 ( .B(T12560_Y), .A(T2452_Y), .Y(T10456_Y));
KC_AND2_X2 T10455 ( .B(T12564_Y), .A(T2452_Y), .Y(T10455_Y));
KC_AND2_X2 T10454 ( .B(T12568_Y), .A(T2452_Y), .Y(T10454_Y));
KC_AND2_X2 T10453 ( .B(T12571_Y), .A(T2452_Y), .Y(T10453_Y));
KC_AND2_X2 T9600 ( .B(T12928_Y), .A(T2452_Y), .Y(T9600_Y));
KC_AND2_X2 T9599 ( .B(T12553_Y), .A(T2452_Y), .Y(T9599_Y));
KC_AND2_X2 T9593 ( .B(T12550_Y), .A(T2452_Y), .Y(T9593_Y));
KC_AND2_X2 T9592 ( .B(T12549_Y), .A(T2452_Y), .Y(T9592_Y));
KC_AND2_X2 T9589 ( .B(T12924_Y), .A(T2452_Y), .Y(T9589_Y));
KC_AND2_X2 T9588 ( .B(T12925_Y), .A(T2452_Y), .Y(T9588_Y));
KC_AND2_X2 T10475 ( .B(T16079_Q), .A(T13710_Q), .Y(T10475_Y));
KC_AND2_X2 T9855 ( .B(T9873_Y), .A(T2529_Y), .Y(T9855_Y));
KC_AND2_X2 T10187 ( .B(T12759_Y), .A(T2651_Y), .Y(T10187_Y));
KC_AND2_X2 T10280 ( .B(T5751_Y), .A(T10278_Y), .Y(T10280_Y));
KC_AND2_X2 T8447 ( .B(T2748_Q), .A(T2738_Q), .Y(T8447_Y));
KC_AND2_X2 T8286 ( .B(T6297_Y), .A(T2783_Y), .Y(T8286_Y));
KC_AND2_X2 T8280 ( .B(T2810_Y), .A(T2810_Y), .Y(T8280_Y));
KC_AND2_X2 T8334 ( .B(T14571_Q), .A(T14572_Q), .Y(T8334_Y));
KC_AND2_X2 T8325 ( .B(T3351_Y), .A(T6024_Y), .Y(T8325_Y));
KC_AND2_X2 T8510 ( .B(T3517_Y), .A(T2618_Q), .Y(T8510_Y));
KC_AND2_X2 T8435 ( .B(T8161_Y), .A(T8162_Y), .Y(T8435_Y));
KC_AND2_X2 T9591 ( .B(T12927_Y), .A(T3025_Y), .Y(T9591_Y));
KC_AND2_X2 T9587 ( .B(T12565_Y), .A(T3025_Y), .Y(T9587_Y));
KC_AND2_X2 T9648 ( .B(T12934_Y), .A(T3025_Y), .Y(T9648_Y));
KC_AND2_X2 T9644 ( .B(T12932_Y), .A(T3025_Y), .Y(T9644_Y));
KC_AND2_X2 T8522 ( .B(T12931_Y), .A(T3025_Y), .Y(T8522_Y));
KC_AND2_X2 T9773 ( .B(T16201_Y), .A(T16201_Y), .Y(T9773_Y));
KC_AND2_X2 T9742 ( .B(T9739_Y), .A(T3678_Y), .Y(T9742_Y));
KC_AND2_X2 T9741 ( .B(T12598_Y), .A(T3678_Y), .Y(T9741_Y));
KC_AND2_X2 T9879 ( .B(T12674_Y), .A(T2651_Y), .Y(T9879_Y));
KC_AND2_X2 T9844 ( .B(T12652_Y), .A(T3678_Y), .Y(T9844_Y));
KC_AND2_X2 T9964 ( .B(T12707_Y), .A(T2651_Y), .Y(T9964_Y));
KC_AND2_X2 T9939 ( .B(T12938_Y), .A(T2651_Y), .Y(T9939_Y));
KC_AND2_X2 T10087 ( .B(T12739_Y), .A(T2651_Y), .Y(T10087_Y));
KC_AND2_X2 T10055 ( .B(T12731_Y), .A(T2651_Y), .Y(T10055_Y));
KC_AND2_X2 T8206 ( .B(T11458_Y), .A(T3282_Y), .Y(T8206_Y));
KC_AND2_X2 T8267 ( .B(T3303_Y), .A(T3295_Y), .Y(T8267_Y));
KC_AND2_X2 T8275 ( .B(T3324_Y), .A(T3332_Y), .Y(T8275_Y));
KC_AND2_X2 T8333 ( .B(T3347_Y), .A(T3349_Y), .Y(T8333_Y));
KC_AND2_X2 T8348 ( .B(T6365_Y), .A(T3414_Y), .Y(T8348_Y));
KC_AND2_X2 T9602 ( .B(T12557_Y), .A(T3025_Y), .Y(T9602_Y));
KC_AND2_X2 T9590 ( .B(T12558_Y), .A(T3025_Y), .Y(T9590_Y));
KC_AND2_X2 T9735 ( .B(T12602_Y), .A(T3682_Y), .Y(T9735_Y));
KC_AND2_X2 T9734 ( .B(T12654_Y), .A(T3682_Y), .Y(T9734_Y));
KC_AND2_X2 T9733 ( .B(T12589_Y), .A(T3682_Y), .Y(T9733_Y));
KC_AND2_X2 T9727 ( .B(T12588_Y), .A(T3682_Y), .Y(T9727_Y));
KC_AND2_X2 T9876 ( .B(T12976_Y), .A(T3682_Y), .Y(T9876_Y));
KC_AND2_X2 T9875 ( .B(T12647_Y), .A(T3682_Y), .Y(T9875_Y));
KC_AND2_X2 T9869 ( .B(T16230_Y), .A(T6846_Y), .Y(T9869_Y));
KC_AND2_X2 T9853 ( .B(T12651_Y), .A(T3682_Y), .Y(T9853_Y));
KC_AND2_X2 T9852 ( .B(T12658_Y), .A(T3682_Y), .Y(T9852_Y));
KC_AND2_X2 T9826 ( .B(T12648_Y), .A(T3682_Y), .Y(T9826_Y));
KC_AND2_X2 T9962 ( .B(T12710_Y), .A(T3682_Y), .Y(T9962_Y));
KC_AND2_X2 T9954 ( .B(T12940_Y), .A(T3682_Y), .Y(T9954_Y));
KC_AND2_X2 T9953 ( .B(T12712_Y), .A(T3682_Y), .Y(T9953_Y));
KC_AND2_X2 T9943 ( .B(T12711_Y), .A(T3682_Y), .Y(T9943_Y));
KC_AND2_X2 T9933 ( .B(T12939_Y), .A(T3682_Y), .Y(T9933_Y));
KC_AND2_X2 T8197 ( .B(T11393_Y), .A(T11375_Y), .Y(T8197_Y));
KC_AND2_X2 T8264 ( .B(T3934_Y), .A(T5937_Y), .Y(T8264_Y));
KC_AND2_X2 T8290 ( .B(T4569_Y), .A(T6265_Y), .Y(T8290_Y));
KC_AND2_X2 T8313 ( .B(T13167_Q), .A(T13145_Q), .Y(T8313_Y));
KC_AND2_X2 T8305 ( .B(T4732_Y), .A(T5573_Q), .Y(T8305_Y));
KC_AND2_X2 T9564 ( .B(T4191_Y), .A(T15365_Y), .Y(T9564_Y));
KC_AND2_X2 T9563 ( .B(T4191_Y), .A(T15365_Y), .Y(T9563_Y));
KC_AND2_X2 T8244 ( .B(T8247_Y), .A(T5885_Y), .Y(T8244_Y));
KC_AND2_X2 T8236 ( .B(T4542_Y), .A(T4539_Y), .Y(T8236_Y));
KC_AND2_X2 T8475 ( .B(T5946_Y), .A(T3953_Y), .Y(T8475_Y));
KC_AND2_X2 T8331 ( .B(T4594_Y), .A(T4605_Y), .Y(T8331_Y));
KC_AND2_X2 T8330 ( .B(T12242_Y), .A(T13153_Y), .Y(T8330_Y));
KC_AND2_X2 T8329 ( .B(T4587_Y), .A(T6344_Y), .Y(T8329_Y));
KC_AND2_X2 T8304 ( .B(T4732_Y), .A(T4629_Q), .Y(T8304_Y));
KC_AND2_X2 T8303 ( .B(T4732_Y), .A(T4626_Q), .Y(T8303_Y));
KC_AND2_X2 T8302 ( .B(T4732_Y), .A(T4628_Q), .Y(T8302_Y));
KC_AND2_X2 T8370 ( .B(T8367_Y), .A(T4661_Y), .Y(T8370_Y));
KC_AND2_X2 T8369 ( .B(T4631_Y), .A(T6166_Y), .Y(T8369_Y));
KC_AND2_X2 T8368 ( .B(T4635_Y), .A(T6166_Y), .Y(T8368_Y));
KC_AND2_X2 T8355 ( .B(T4636_Y), .A(T6166_Y), .Y(T8355_Y));
KC_AND2_X2 T8390 ( .B(T4697_Y), .A(T16122_Y), .Y(T8390_Y));
KC_AND2_X2 T9467 ( .B(T977_Q), .A(T9461_Q), .Y(T9467_Y));
KC_AND2_X2 T9466 ( .B(T977_Q), .A(T9460_Q), .Y(T9466_Y));
KC_AND2_X2 T9465 ( .B(T977_Q), .A(T770_Q), .Y(T9465_Y));
KC_AND2_X2 T9464 ( .B(T977_Q), .A(T780_Q), .Y(T9464_Y));
KC_AND2_X2 T9442 ( .B(T972_Y), .A(T9439_Y), .Y(T9442_Y));
KC_AND2_X2 T9441 ( .B(T972_Y), .A(T10297_Y), .Y(T9441_Y));
KC_AND2_X2 T9468 ( .B(T977_Q), .A(T5407_Q), .Y(T9468_Y));
KC_AND2_X2 T9434 ( .B(T972_Y), .A(T9032_Y), .Y(T9434_Y));
KC_AND2_X2 T9433 ( .B(T972_Y), .A(T8997_Y), .Y(T9433_Y));
KC_AND2_X2 T10402 ( .B(T12531_Y), .A(T1431_Y), .Y(T10402_Y));
KC_AND2_X2 T10401 ( .B(T12546_Y), .A(T1431_Y), .Y(T10401_Y));
KC_AND2_X2 T10323 ( .B(T12898_Y), .A(T1491_Y), .Y(T10323_Y));
KC_AND2_X2 T10394 ( .B(T12916_Y), .A(T1418_Y), .Y(T10394_Y));
KC_AND2_X2 T10349 ( .B(T12918_Y), .A(T1930_Y), .Y(T10349_Y));
KC_AND2_X2 T10348 ( .B(T12555_Y), .A(T1930_Y), .Y(T10348_Y));
KC_AND2_X2 T10444 ( .B(T12573_Y), .A(T2452_Y), .Y(T10444_Y));
KC_AND2_X2 T10448 ( .B(T12562_Y), .A(T2452_Y), .Y(T10448_Y));
KC_AND2_X2 T10447 ( .B(T12563_Y), .A(T2452_Y), .Y(T10447_Y));
KC_AND2_X2 T10446 ( .B(T12561_Y), .A(T2452_Y), .Y(T10446_Y));
KC_AND2_X2 T8446 ( .B(T2749_Q), .A(T2737_Q), .Y(T8446_Y));
KC_AND2_X2 T16260 ( .B(T16254_Y), .A(T2651_Y), .Y(T16260_Y));
KC_AND2_X2 T10508 ( .B(T12673_Y), .A(T2651_Y), .Y(T10508_Y));
KC_AND2_X2 T8488 ( .B(T5064_Y), .A(T3299_Y), .Y(T8488_Y));
KC_AND2_X2 T10492 ( .B(T12653_Y), .A(T3682_Y), .Y(T10492_Y));
KC_AND2_X2 T10491 ( .B(T12659_Y), .A(T3682_Y), .Y(T10491_Y));
KC_AND2_X2 T8465 ( .B(T4732_Y), .A(T15815_Q), .Y(T8465_Y));
KC_AND2_X2 T8464 ( .B(T4732_Y), .A(T4627_Q), .Y(T8464_Y));
KC_AND2_X2 T8463 ( .B(T4732_Y), .A(T4630_Q), .Y(T8463_Y));
KC_AND2_X2 T10409 ( .B(T12946_Y), .A(T1930_Y), .Y(T10409_Y));
KC_AND2_X2 T10351 ( .B(T12592_Y), .A(T1930_Y), .Y(T10351_Y));
KC_AND2_X2 T9740 ( .B(T12595_Y), .A(T3678_Y), .Y(T9740_Y));
KC_AND2_X2 T9713 ( .B(T12538_Y), .A(T1453_Y), .Y(T9713_Y));
KC_AND2_X2 T8937 ( .B(T972_Y), .A(T1471_Y), .Y(T8937_Y));
KC_AND2_X2 T10285 ( .B(T10725_Y), .A(T1372_Y), .Y(T10285_Y));
KC_AND2_X2 T10193 ( .B(T12764_Y), .A(T2651_Y), .Y(T10193_Y));
KC_AND2_X2 T10186 ( .B(T12766_Y), .A(T2651_Y), .Y(T10186_Y));
KC_AND2_X2 T10182 ( .B(T12765_Y), .A(T2651_Y), .Y(T10182_Y));
KC_AND2_X2 T10181 ( .B(T12767_Y), .A(T2651_Y), .Y(T10181_Y));
KC_AND2_X2 T8301 ( .B(T4732_Y), .A(T5488_Q), .Y(T8301_Y));
KC_AND2_X2 T8436 ( .B(T6495_Y), .A(T6544_Y), .Y(T8436_Y));
KC_AND2_X2 T8426 ( .B(T4096_Y), .A(T11043_Y), .Y(T8426_Y));
KC_AND2_X2 T16255 ( .B(T12748_Y), .A(T2651_Y), .Y(T16255_Y));
KC_AND2_X2 T10350 ( .B(T12948_Y), .A(T1930_Y), .Y(T10350_Y));
KC_AOI21B_X2 T9012 ( .A0(T9014_Y), .BN(T1423_Y), .Y(T9012_Y),     .A1(T15097_Y));
KC_AOI21B_X2 T8982 ( .A0(T9442_Y), .BN(T7898_Y), .Y(T8982_Y),     .A1(T9017_Y));
KC_AOI21B_X2 T10646 ( .A0(T15244_Y), .BN(T10842_Y), .Y(T10646_Y),     .A1(T13432_Q));
KC_AOI21B_X2 T10645 ( .A0(T13438_Q), .BN(T10845_Y), .Y(T10645_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T10644 ( .A0(T13432_Q), .BN(T6885_Y), .Y(T10644_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9562 ( .A0(T15244_Y), .BN(T7041_Y), .Y(T9562_Y),     .A1(T13438_Q));
KC_AOI21B_X2 T9561 ( .A0(T13435_Q), .BN(T6897_Y), .Y(T9561_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9560 ( .A0(T15244_Y), .BN(T7042_Y), .Y(T9560_Y),     .A1(T13337_Q));
KC_AOI21B_X2 T9559 ( .A0(T15244_Y), .BN(T10843_Y), .Y(T9559_Y),     .A1(T13435_Q));
KC_AOI21B_X2 T9558 ( .A0(T14587_Q), .BN(T6884_Y), .Y(T9558_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9555 ( .A0(T15244_Y), .BN(T6888_Y), .Y(T9555_Y),     .A1(T14587_Q));
KC_AOI21B_X2 T9554 ( .A0(T15244_Y), .BN(T6896_Y), .Y(T9554_Y),     .A1(T13434_Q));
KC_AOI21B_X2 T9553 ( .A0(T13434_Q), .BN(T10844_Y), .Y(T9553_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9538 ( .A0(T13337_Q), .BN(T10846_Y), .Y(T9538_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T10430 ( .A0(T13727_Q), .BN(T7333_Y), .Y(T10430_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T10429 ( .A0(T13740_Q), .BN(T7331_Y), .Y(T10429_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9628 ( .A0(T1337_Y), .BN(T7343_Y), .Y(T9628_Y),     .A1(T13727_Q));
KC_AOI21B_X2 T9627 ( .A0(T1337_Y), .BN(T7332_Y), .Y(T9627_Y),     .A1(T13740_Q));
KC_AOI21B_X2 T9702 ( .A0(T1337_Y), .BN(T5697_Y), .Y(T9702_Y),     .A1(T13840_Q));
KC_AOI21B_X2 T9701 ( .A0(T13840_Q), .BN(T5698_Y), .Y(T9701_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T8934 ( .A0(T8032_Y), .BN(T8938_Y), .Y(T8934_Y),     .A1(T139_Y));
KC_AOI21B_X2 T10383 ( .A0(T15244_Y), .BN(T6883_Y), .Y(T10383_Y),     .A1(T13502_Q));
KC_AOI21B_X2 T9557 ( .A0(T13502_Q), .BN(T6887_Y), .Y(T9557_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9556 ( .A0(T13352_Q), .BN(T6886_Y), .Y(T9556_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9552 ( .A0(T15244_Y), .BN(T6880_Y), .Y(T9552_Y),     .A1(T13503_Q));
KC_AOI21B_X2 T9550 ( .A0(T15244_Y), .BN(T6877_Y), .Y(T9550_Y),     .A1(T14680_Q));
KC_AOI21B_X2 T9549 ( .A0(T15244_Y), .BN(T6875_Y), .Y(T9549_Y),     .A1(T13350_Q));
KC_AOI21B_X2 T9548 ( .A0(T14680_Q), .BN(T6895_Y), .Y(T9548_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9547 ( .A0(T15244_Y), .BN(T6879_Y), .Y(T9547_Y),     .A1(T13501_Q));
KC_AOI21B_X2 T9537 ( .A0(T13501_Q), .BN(T6878_Y), .Y(T9537_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9535 ( .A0(T13350_Q), .BN(T6881_Y), .Y(T9535_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9534 ( .A0(T13503_Q), .BN(T6882_Y), .Y(T9534_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9625 ( .A0(T13723_Q), .BN(T7330_Y), .Y(T9625_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9616 ( .A0(T1337_Y), .BN(T7352_Y), .Y(T9616_Y),     .A1(T13729_Q));
KC_AOI21B_X2 T9615 ( .A0(T1337_Y), .BN(T7321_Y), .Y(T9615_Y),     .A1(T13723_Q));
KC_AOI21B_X2 T10340 ( .A0(T1337_Y), .BN(T7473_Y), .Y(T10340_Y),     .A1(T13866_Q));
KC_AOI21B_X2 T9722 ( .A0(T13870_Q), .BN(T7498_Y), .Y(T9722_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9703 ( .A0(T1337_Y), .BN(T7497_Y), .Y(T9703_Y),     .A1(T13870_Q));
KC_AOI21B_X2 T9807 ( .A0(T14004_Q), .BN(T10795_Y), .Y(T9807_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9806 ( .A0(T1337_Y), .BN(T7768_Y), .Y(T9806_Y),     .A1(T14004_Q));
KC_AOI21B_X2 T9805 ( .A0(T1337_Y), .BN(T10794_Y), .Y(T9805_Y),     .A1(T14007_Q));
KC_AOI21B_X2 T10381 ( .A0(T15244_Y), .BN(T10837_Y), .Y(T10381_Y),     .A1(T13498_Q));
KC_AOI21B_X2 T9551 ( .A0(T15244_Y), .BN(T10838_Y), .Y(T9551_Y),     .A1(T14681_Q));
KC_AOI21B_X2 T9546 ( .A0(T14679_Q), .BN(T10840_Y), .Y(T9546_Y),     .A1(T15244_Y));
KC_AOI21B_X2 T9545 ( .A0(T15244_Y), .BN(T7040_Y), .Y(T9545_Y),     .A1(T13499_Q));
KC_AOI21B_X2 T9544 ( .A0(T13499_Q), .BN(T10839_Y), .Y(T9544_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9536 ( .A0(T14681_Q), .BN(T6874_Y), .Y(T9536_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9533 ( .A0(T13498_Q), .BN(T6872_Y), .Y(T9533_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9532 ( .A0(T14679_Q), .BN(T6876_Y), .Y(T9532_Y),     .A1(T15198_Y));
KC_AOI21B_X2 T9624 ( .A0(T13721_Q), .BN(T7326_Y), .Y(T9624_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9623 ( .A0(T1337_Y), .BN(T7328_Y), .Y(T9623_Y),     .A1(T13724_Q));
KC_AOI21B_X2 T9622 ( .A0(T13724_Q), .BN(T7329_Y), .Y(T9622_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9621 ( .A0(T1337_Y), .BN(T7327_Y), .Y(T9621_Y),     .A1(T13721_Q));
KC_AOI21B_X2 T9620 ( .A0(T1337_Y), .BN(T7325_Y), .Y(T9620_Y),     .A1(T13695_Q));
KC_AOI21B_X2 T9619 ( .A0(T13695_Q), .BN(T7324_Y), .Y(T9619_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T10339 ( .A0(T14648_Q), .BN(T7758_Y), .Y(T10339_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T10337 ( .A0(T1337_Y), .BN(T10789_Y), .Y(T10337_Y),     .A1(T14648_Q));
KC_AOI21B_X2 T9804 ( .A0(T1337_Y), .BN(T7763_Y), .Y(T9804_Y),     .A1(T13982_Q));
KC_AOI21B_X2 T9802 ( .A0(T14001_Q), .BN(T7759_Y), .Y(T9802_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9801 ( .A0(T13997_Q), .BN(T10786_Y), .Y(T9801_Y),     .A1(T1337_Y));
KC_AOI21B_X2 T9800 ( .A0(T13997_Q), .BN(T10784_Y), .Y(T9800_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9799 ( .A0(T13982_Q), .BN(T7764_Y), .Y(T9799_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9798 ( .A0(T1337_Y), .BN(T10785_Y), .Y(T9798_Y),     .A1(T14001_Q));
KC_AOI21B_X2 T10312 ( .A0(T10743_Y), .BN(T10716_Y), .Y(T10312_Y),     .A1(T14282_Q));
KC_AOI21B_X2 T9909 ( .A0(T10743_Y), .BN(T7946_Y), .Y(T9909_Y),     .A1(T14122_Q));
KC_AOI21B_X2 T9908 ( .A0(T14122_Q), .BN(T7947_Y), .Y(T9908_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T9887 ( .A0(T14110_Q), .BN(T10753_Y), .Y(T9887_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T9886 ( .A0(T14282_Q), .BN(T10689_Y), .Y(T9886_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T9885 ( .A0(T10743_Y), .BN(T10751_Y), .Y(T9885_Y),     .A1(T14110_Q));
KC_AOI21B_X2 T10036 ( .A0(T14258_Q), .BN(T10695_Y), .Y(T10036_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10019 ( .A0(T10743_Y), .BN(T10692_Y), .Y(T10019_Y),     .A1(T14258_Q));
KC_AOI21B_X2 T9979 ( .A0(T10743_Y), .BN(T10657_Y), .Y(T9979_Y),     .A1(T14598_Q));
KC_AOI21B_X2 T9978 ( .A0(T10743_Y), .BN(T4832_Y), .Y(T9978_Y),     .A1(T14386_Q));
KC_AOI21B_X2 T10151 ( .A0(T14386_Q), .BN(T10732_Y), .Y(T10151_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10122 ( .A0(T10724_Y), .BN(T10285_Y), .Y(T10122_Y),     .A1(T1738_Y));
KC_AOI21B_X2 T10357 ( .A0(T14660_Q), .BN(T7535_Y), .Y(T10357_Y),     .A1(T15235_Y));
KC_AOI21B_X2 T9709 ( .A0(T13814_Q), .BN(T7538_Y), .Y(T9709_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9708 ( .A0(T14660_Q), .BN(T7487_Y), .Y(T9708_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9697 ( .A0(T13834_Q), .BN(T7536_Y), .Y(T9697_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9797 ( .A0(T13994_Q), .BN(T7755_Y), .Y(T9797_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9796 ( .A0(T15235_Y), .BN(T7756_Y), .Y(T9796_Y),     .A1(T13956_Q));
KC_AOI21B_X2 T10311 ( .A0(T10743_Y), .BN(T10712_Y), .Y(T10311_Y),     .A1(T14271_Q));
KC_AOI21B_X2 T9884 ( .A0(T14271_Q), .BN(T10747_Y), .Y(T9884_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10150 ( .A0(T10743_Y), .BN(T10730_Y), .Y(T10150_Y),     .A1(T14385_Q));
KC_AOI21B_X2 T10149 ( .A0(T14385_Q), .BN(T10731_Y), .Y(T10149_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10148 ( .A0(T10743_Y), .BN(T5399_Y), .Y(T10148_Y),     .A1(T14380_Q));
KC_AOI21B_X2 T10126 ( .A0(T10743_Y), .BN(T1512_Y), .Y(T10126_Y),     .A1(T14592_Q));
KC_AOI21B_X2 T10376 ( .A0(T15201_Y), .BN(T6864_Y), .Y(T10376_Y),     .A1(T13342_Q));
KC_AOI21B_X2 T10375 ( .A0(T13342_Q), .BN(T6863_Y), .Y(T10375_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T10385 ( .A0(T15201_Y), .BN(T10867_Y), .Y(T10385_Y),     .A1(T14687_Q));
KC_AOI21B_X2 T10384 ( .A0(T14687_Q), .BN(T10848_Y), .Y(T10384_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9629 ( .A0(T15201_Y), .BN(T10870_Y), .Y(T9629_Y),     .A1(T13689_Q));
KC_AOI21B_X2 T9717 ( .A0(T15235_Y), .BN(T7532_Y), .Y(T9717_Y),     .A1(T13806_Q));
KC_AOI21B_X2 T9716 ( .A0(T13805_Q), .BN(T7521_Y), .Y(T9716_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9715 ( .A0(T15235_Y), .BN(T7524_Y), .Y(T9715_Y),     .A1(T13805_Q));
KC_AOI21B_X2 T9711 ( .A0(T15235_Y), .BN(T7537_Y), .Y(T9711_Y),     .A1(T13834_Q));
KC_AOI21B_X2 T9710 ( .A0(T15235_Y), .BN(T7529_Y), .Y(T9710_Y),     .A1(T13814_Q));
KC_AOI21B_X2 T9695 ( .A0(T13784_Q), .BN(T10766_Y), .Y(T9695_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9795 ( .A0(T15235_Y), .BN(T7743_Y), .Y(T9795_Y),     .A1(T13994_Q));
KC_AOI21B_X2 T10728 ( .A0(T14594_Q), .BN(T4893_Y), .Y(T10728_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10147 ( .A0(T14378_Q), .BN(T10729_Y), .Y(T10147_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10145 ( .A0(T14377_Q), .BN(T5400_Y), .Y(T10145_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10133 ( .A0(T10743_Y), .BN(T1606_Y), .Y(T10133_Y),     .A1(T14377_Q));
KC_AOI21B_X2 T10125 ( .A0(T10743_Y), .BN(T10726_Y), .Y(T10125_Y),     .A1(T14372_Q));
KC_AOI21B_X2 T10121 ( .A0(T10743_Y), .BN(T1607_Y), .Y(T10121_Y),     .A1(T14594_Q));
KC_AOI21B_X2 T10464 ( .A0(T15201_Y), .BN(T5178_Y), .Y(T10464_Y),     .A1(T13431_Q));
KC_AOI21B_X2 T10379 ( .A0(T15201_Y), .BN(T6892_Y), .Y(T10379_Y),     .A1(T14676_Q));
KC_AOI21B_X2 T10378 ( .A0(T15201_Y), .BN(T6869_Y), .Y(T10378_Y),     .A1(T13344_Q));
KC_AOI21B_X2 T10377 ( .A0(T13344_Q), .BN(T10835_Y), .Y(T10377_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9531 ( .A0(T13431_Q), .BN(T1618_Y), .Y(T9531_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9521 ( .A0(T13339_Q), .BN(T6865_Y), .Y(T9521_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9520 ( .A0(T14676_Q), .BN(T6867_Y), .Y(T9520_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9519 ( .A0(T15201_Y), .BN(T6893_Y), .Y(T9519_Y),     .A1(T13339_Q));
KC_AOI21B_X2 T9518 ( .A0(T13371_Q), .BN(T6868_Y), .Y(T9518_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9517 ( .A0(T15201_Y), .BN(T6866_Y), .Y(T9517_Y),     .A1(T13371_Q));
KC_AOI21B_X2 T9584 ( .A0(T13580_Q), .BN(T7170_Y), .Y(T9584_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9583 ( .A0(T15201_Y), .BN(T7169_Y), .Y(T9583_Y),     .A1(T13580_Q));
KC_AOI21B_X2 T10497 ( .A0(T15235_Y), .BN(T10769_Y), .Y(T10497_Y),     .A1(T13986_Q));
KC_AOI21B_X2 T9751 ( .A0(T13986_Q), .BN(T1639_Y), .Y(T9751_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9750 ( .A0(T15235_Y), .BN(T10768_Y), .Y(T9750_Y),     .A1(T13931_Q));
KC_AOI21B_X2 T9694 ( .A0(T13931_Q), .BN(T7462_Y), .Y(T9694_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9693 ( .A0(T13973_Q), .BN(T10767_Y), .Y(T9693_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9692 ( .A0(T15235_Y), .BN(T10763_Y), .Y(T9692_Y),     .A1(T13973_Q));
KC_AOI21B_X2 T9691 ( .A0(T14628_Q), .BN(T7460_Y), .Y(T9691_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9690 ( .A0(T15235_Y), .BN(T10764_Y), .Y(T9690_Y),     .A1(T14628_Q));
KC_AOI21B_X2 T9689 ( .A0(T15235_Y), .BN(T10770_Y), .Y(T9689_Y),     .A1(T13784_Q));
KC_AOI21B_X2 T8311 ( .A0(T11728_Y), .BN(T2266_Y), .Y(T8311_Y),     .A1(T1790_Q));
KC_AOI21B_X2 T8375 ( .A0(T4965_Y), .BN(T2283_Y), .Y(T8375_Y),     .A1(T4925_Q));
KC_AOI21B_X2 T8364 ( .A0(T4965_Y), .BN(T2268_Y), .Y(T8364_Y),     .A1(T1823_Q));
KC_AOI21B_X2 T8434 ( .A0(T2400_Y), .BN(T2339_Y), .Y(T8434_Y),     .A1(T1847_Y));
KC_AOI21B_X2 T10463 ( .A0(T15201_Y), .BN(T1861_Y), .Y(T10463_Y),     .A1(T13429_Q));
KC_AOI21B_X2 T10462 ( .A0(T15201_Y), .BN(T1860_Y), .Y(T10462_Y),     .A1(T13430_Q));
KC_AOI21B_X2 T9530 ( .A0(T13430_Q), .BN(T1859_Y), .Y(T9530_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9603 ( .A0(T13641_Q), .BN(T1909_Y), .Y(T9603_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9598 ( .A0(T13659_Q), .BN(T1911_Y), .Y(T9598_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9597 ( .A0(T15201_Y), .BN(T1910_Y), .Y(T9597_Y),     .A1(T13659_Q));
KC_AOI21B_X2 T9596 ( .A0(T15201_Y), .BN(T5739_Y), .Y(T9596_Y),     .A1(T13641_Q));
KC_AOI21B_X2 T9595 ( .A0(T15201_Y), .BN(T1908_Y), .Y(T9595_Y),     .A1(T13643_Q));
KC_AOI21B_X2 T9594 ( .A0(T13643_Q), .BN(T1912_Y), .Y(T9594_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9851 ( .A0(T15235_Y), .BN(T1968_Y), .Y(T9851_Y),     .A1(T14053_Q));
KC_AOI21B_X2 T9850 ( .A0(T14053_Q), .BN(T5286_Y), .Y(T9850_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T8297 ( .A0(T11620_Y), .BN(T2208_Y), .Y(T8297_Y),     .A1(T5463_Q));
KC_AOI21B_X2 T8173 ( .A0(T5527_Q), .BN(T2335_Y), .Y(T8173_Y),     .A1(T2364_Q));
KC_AOI21B_X2 T8160 ( .A0(T2376_Y), .BN(T2947_Y), .Y(T8160_Y),     .A1(T2947_Y));
KC_AOI21B_X2 T9848 ( .A0(T2535_Y), .BN(T3064_Y), .Y(T9848_Y),     .A1(T7346_Y));
KC_AOI21B_X2 T9847 ( .A0(T2535_Y), .BN(T3063_Y), .Y(T9847_Y),     .A1(T10398_Y));
KC_AOI21B_X2 T9846 ( .A0(T2535_Y), .BN(T3067_Y), .Y(T9846_Y),     .A1(T7039_Y));
KC_AOI21B_X2 T9845 ( .A0(T2535_Y), .BN(T3065_Y), .Y(T9845_Y),     .A1(T7126_Y));
KC_AOI21B_X2 T9947 ( .A0(T2577_Y), .BN(T5869_S), .Y(T9947_Y),     .A1(T2577_Y));
KC_AOI21B_X2 T10537 ( .A0(T15689_Y), .BN(T10536_Y), .Y(T10537_Y),     .A1(T2649_Y));
KC_AOI21B_X2 T8269 ( .A0(T5456_Y), .BN(T5941_Y), .Y(T8269_Y),     .A1(T2734_Y));
KC_AOI21B_X2 T10461 ( .A0(T15251_Y), .BN(T2968_Y), .Y(T10461_Y),     .A1(T13508_Q));
KC_AOI21B_X2 T10460 ( .A0(T13508_Q), .BN(T5177_Y), .Y(T10460_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9529 ( .A0(T15251_Y), .BN(T2969_Y), .Y(T9529_Y),     .A1(T13391_Q));
KC_AOI21B_X2 T9528 ( .A0(T15251_Y), .BN(T5179_Y), .Y(T9528_Y),     .A1(T13407_Q));
KC_AOI21B_X2 T9527 ( .A0(T13407_Q), .BN(T5181_Y), .Y(T9527_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9526 ( .A0(T13391_Q), .BN(T5180_Y), .Y(T9526_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9572 ( .A0(T15251_Y), .BN(T5210_Y), .Y(T9572_Y),     .A1(T13542_Q));
KC_AOI21B_X2 T9571 ( .A0(T13424_Q), .BN(T5216_Y), .Y(T9571_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9570 ( .A0(T15251_Y), .BN(T2993_Y), .Y(T9570_Y),     .A1(T13424_Q));
KC_AOI21B_X2 T9569 ( .A0(T13542_Q), .BN(T5215_Y), .Y(T9569_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9568 ( .A0(T13525_Q), .BN(T2988_Y), .Y(T9568_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9567 ( .A0(T15251_Y), .BN(T2982_Y), .Y(T9567_Y),     .A1(T13525_Q));
KC_AOI21B_X2 T10488 ( .A0(T14854_Q), .BN(T3028_Y), .Y(T10488_Y),     .A1(T3636_Y));
KC_AOI21B_X2 T10487 ( .A0(T14854_Q), .BN(T3066_Y), .Y(T10487_Y),     .A1(T3054_Y));
KC_AOI21B_X2 T10486 ( .A0(T3636_Y), .BN(T3029_Y), .Y(T10486_Y),     .A1(T14050_Q));
KC_AOI21B_X2 T9777 ( .A0(T13928_Q), .BN(T5266_Y), .Y(T9777_Y),     .A1(T3054_Y));
KC_AOI21B_X2 T9776 ( .A0(T3636_Y), .BN(T3612_Y), .Y(T9776_Y),     .A1(T13928_Q));
KC_AOI21B_X2 T9934 ( .A0(T14182_Q), .BN(T3715_Y), .Y(T9934_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T8230 ( .A0(T15129_Y), .BN(T3250_Y), .Y(T8230_Y),     .A1(T15929_Y));
KC_AOI21B_X2 T8215 ( .A0(T4384_Y), .BN(T8206_Y), .Y(T8215_Y),     .A1(T4384_Y));
KC_AOI21B_X2 T8323 ( .A0(T15134_Y), .BN(T8333_Y), .Y(T8323_Y),     .A1(T8322_Y));
KC_AOI21B_X2 T8393 ( .A0(T12284_Y), .BN(T12284_Y), .Y(T8393_Y),     .A1(T12284_Y));
KC_AOI21B_X2 T10459 ( .A0(T15251_Y), .BN(T3539_Y), .Y(T10459_Y),     .A1(T14812_Q));
KC_AOI21B_X2 T10458 ( .A0(T14812_Q), .BN(T4183_Y), .Y(T10458_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9525 ( .A0(T13421_Q), .BN(T5182_Y), .Y(T9525_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9524 ( .A0(T15251_Y), .BN(T4182_Y), .Y(T9524_Y),     .A1(T13421_Q));
KC_AOI21B_X2 T9523 ( .A0(T13389_Q), .BN(T3542_Y), .Y(T9523_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9522 ( .A0(T15251_Y), .BN(T3543_Y), .Y(T9522_Y),     .A1(T13389_Q));
KC_AOI21B_X2 T10450 ( .A0(T15251_Y), .BN(T3559_Y), .Y(T10450_Y),     .A1(T14792_Q));
KC_AOI21B_X2 T10449 ( .A0(T15251_Y), .BN(T3557_Y), .Y(T10449_Y),     .A1(T14793_Q));
KC_AOI21B_X2 T9566 ( .A0(T14792_Q), .BN(T3560_Y), .Y(T9566_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9565 ( .A0(T14793_Q), .BN(T3562_Y), .Y(T9565_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T474 ( .A0(T15251_Y), .BN(T3591_Y), .Y(T474_Y),     .A1(T14757_Q));
KC_AOI21B_X2 T473 ( .A0(T13753_Q), .BN(T5248_Y), .Y(T473_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9662 ( .A0(T15251_Y), .BN(T3592_Y), .Y(T9662_Y),     .A1(T13752_Q));
KC_AOI21B_X2 T9661 ( .A0(T15251_Y), .BN(T5247_Y), .Y(T9661_Y),     .A1(T13753_Q));
KC_AOI21B_X2 T9660 ( .A0(T13752_Q), .BN(T3599_Y), .Y(T9660_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T9634 ( .A0(T14757_Q), .BN(T3593_Y), .Y(T9634_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T10513 ( .A0(T15253_Y), .BN(T3733_Y), .Y(T10513_Y),     .A1(T14301_Q));
KC_AOI21B_X2 T9963 ( .A0(T14301_Q), .BN(T3694_Y), .Y(T9963_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T9956 ( .A0(T14170_Q), .BN(T3703_Y), .Y(T9956_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T9955 ( .A0(T15253_Y), .BN(T3704_Y), .Y(T9955_Y),     .A1(T14170_Q));
KC_AOI21B_X2 T9945 ( .A0(T14195_Q), .BN(T3699_Y), .Y(T9945_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T9944 ( .A0(T14195_Q), .BN(T3698_Y), .Y(T9944_Y),     .A1(T15253_Y));
KC_AOI21B_X2 T9935 ( .A0(T15253_Y), .BN(T3718_Y), .Y(T9935_Y),     .A1(T14182_Q));
KC_AOI21B_X2 T10117 ( .A0(T15253_Y), .BN(T3722_Y), .Y(T10117_Y),     .A1(T14356_Q));
KC_AOI21B_X2 T10116 ( .A0(T14356_Q), .BN(T3723_Y), .Y(T10116_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10098 ( .A0(T15253_Y), .BN(T3727_Y), .Y(T10098_Y),     .A1(T14324_Q));
KC_AOI21B_X2 T10097 ( .A0(T14324_Q), .BN(T3726_Y), .Y(T10097_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10076 ( .A0(T14297_Q), .BN(T3732_Y), .Y(T10076_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10075 ( .A0(T14314_Q), .BN(T3729_Y), .Y(T10075_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10074 ( .A0(T15253_Y), .BN(T3730_Y), .Y(T10074_Y),     .A1(T14314_Q));
KC_AOI21B_X2 T10053 ( .A0(T15253_Y), .BN(T3734_Y), .Y(T10053_Y),     .A1(T14297_Q));
KC_AOI21B_X2 T8507 ( .A0(T6077_Y), .BN(T12291_Y), .Y(T8507_Y),     .A1(T12965_Y));
KC_AOI21B_X2 T8386 ( .A0(T15623_Y), .BN(T12268_Y), .Y(T8386_Y),     .A1(T3443_Y));
KC_AOI21B_X2 T8380 ( .A0(T8382_Y), .BN(T10563_Y), .Y(T8380_Y),     .A1(T4077_Y));
KC_AOI21B_X2 T8519 ( .A0(T14914_Q), .BN(T4218_Y), .Y(T8519_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T8518 ( .A0(T14912_Q), .BN(T4221_Y), .Y(T8518_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T8517 ( .A0(T15214_Y), .BN(T4220_Y), .Y(T8517_Y),     .A1(T13748_Q));
KC_AOI21B_X2 T8516 ( .A0(T13748_Q), .BN(T4217_Y), .Y(T8516_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9775 ( .A0(T13924_Q), .BN(T4233_Y), .Y(T9775_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9762 ( .A0(T13890_Q), .BN(T4244_Y), .Y(T9762_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9761 ( .A0(T15214_Y), .BN(T4248_Y), .Y(T9761_Y),     .A1(T13890_Q));
KC_AOI21B_X2 T9726 ( .A0(T15214_Y), .BN(T4234_Y), .Y(T9726_Y),     .A1(T13924_Q));
KC_AOI21B_X2 T9725 ( .A0(T15214_Y), .BN(T4256_Y), .Y(T9725_Y),     .A1(T13873_Q));
KC_AOI21B_X2 T9724 ( .A0(T13873_Q), .BN(T4257_Y), .Y(T9724_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9857 ( .A0(T15214_Y), .BN(T4269_Y), .Y(T9857_Y),     .A1(T14039_Q));
KC_AOI21B_X2 T9856 ( .A0(T14039_Q), .BN(T4270_Y), .Y(T9856_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9821 ( .A0(T14086_Q), .BN(T4263_Y), .Y(T9821_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9820 ( .A0(T15214_Y), .BN(T4264_Y), .Y(T9820_Y),     .A1(T14086_Q));
KC_AOI21B_X2 T10512 ( .A0(T14284_Q), .BN(T4293_Y), .Y(T10512_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T10499 ( .A0(T14873_Q), .BN(T4315_Y), .Y(T10499_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9961 ( .A0(T15214_Y), .BN(T4304_Y), .Y(T9961_Y),     .A1(T4317_Y));
KC_AOI21B_X2 T9960 ( .A0(T15214_Y), .BN(T4295_Y), .Y(T9960_Y),     .A1(T14187_Q));
KC_AOI21B_X2 T9959 ( .A0(T14187_Q), .BN(T4294_Y), .Y(T9959_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9952 ( .A0(T4317_Y), .BN(T4300_Y), .Y(T9952_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9931 ( .A0(T15214_Y), .BN(T4310_Y), .Y(T9931_Y),     .A1(T14141_Q));
KC_AOI21B_X2 T9930 ( .A0(T14141_Q), .BN(T4311_Y), .Y(T9930_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T9929 ( .A0(T15214_Y), .BN(T4316_Y), .Y(T9929_Y),     .A1(T14873_Q));
KC_AOI21B_X2 T10114 ( .A0(T15253_Y), .BN(T4319_Y), .Y(T10114_Y),     .A1(T14348_Q));
KC_AOI21B_X2 T10073 ( .A0(T14319_Q), .BN(T4323_Y), .Y(T10073_Y),     .A1(T15214_Y));
KC_AOI21B_X2 T10072 ( .A0(T14319_Q), .BN(T4321_Y), .Y(T10072_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T10052 ( .A0(T14305_Q), .BN(T4322_Y), .Y(T10052_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T10051 ( .A0(T15214_Y), .BN(T4324_Y), .Y(T10051_Y),     .A1(T14284_Q));
KC_AOI21B_X2 T10050 ( .A0(T15214_Y), .BN(T4325_Y), .Y(T10050_Y),     .A1(T14305_Q));
KC_AOI21B_X2 T10533 ( .A0(T14897_Q), .BN(T4338_Y), .Y(T10533_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10200 ( .A0(T15253_Y), .BN(T5975_Y), .Y(T10200_Y),     .A1(T14502_Q));
KC_AOI21B_X2 T10199 ( .A0(T15253_Y), .BN(T4339_Y), .Y(T10199_Y),     .A1(T14897_Q));
KC_AOI21B_X2 T10198 ( .A0(T15253_Y), .BN(T4340_Y), .Y(T10198_Y),     .A1(T14899_Q));
KC_AOI21B_X2 T10197 ( .A0(T14436_Q), .BN(T4342_Y), .Y(T10197_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10196 ( .A0(T15253_Y), .BN(T4343_Y), .Y(T10196_Y),     .A1(T14436_Q));
KC_AOI21B_X2 T10192 ( .A0(T14428_Q), .BN(T4344_Y), .Y(T10192_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10190 ( .A0(T15253_Y), .BN(T4345_Y), .Y(T10190_Y),     .A1(T14428_Q));
KC_AOI21B_X2 T10189 ( .A0(T14502_Q), .BN(T5974_Y), .Y(T10189_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10179 ( .A0(T14409_Q), .BN(T4346_Y), .Y(T10179_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10178 ( .A0(T15253_Y), .BN(T4348_Y), .Y(T10178_Y),     .A1(T14409_Q));
KC_AOI21B_X2 T10177 ( .A0(T14408_Q), .BN(T4347_Y), .Y(T10177_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10176 ( .A0(T15253_Y), .BN(T4349_Y), .Y(T10176_Y),     .A1(T14408_Q));
KC_AOI21B_X2 T8178 ( .A0(T16241_Y), .BN(T11381_Y), .Y(T8178_Y),     .A1(T11365_Y));
KC_AOI21B_X2 T8321 ( .A0(T6327_Y), .BN(T6023_Y), .Y(T8321_Y),     .A1(T6009_Y));
KC_AOI21B_X2 T8300 ( .A0(T4623_Y), .BN(T13309_Y), .Y(T8300_Y),     .A1(T8455_Y));
KC_AOI21B_X2 T8367 ( .A0(T4690_Y), .BN(T4665_Y), .Y(T8367_Y),     .A1(T4668_Y));
KC_AOI21B_X2 T10342 ( .A0(T14007_Q), .BN(T10793_Y), .Y(T10342_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T10292 ( .A0(T14388_Q), .BN(T10735_Y), .Y(T10292_Y),     .A1(T10743_Y));
KC_AOI21B_X2 T10291 ( .A0(T14598_Q), .BN(T10741_Y), .Y(T10291_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10290 ( .A0(T14388_Q), .BN(T10736_Y), .Y(T10290_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10395 ( .A0(T14722_Q), .BN(T10871_Y), .Y(T10395_Y),     .A1(T15201_Y));
KC_AOI21B_X2 T10289 ( .A0(T10743_Y), .BN(T10733_Y), .Y(T10289_Y),     .A1(T14384_Q));
KC_AOI21B_X2 T10288 ( .A0(T14384_Q), .BN(T10734_Y), .Y(T10288_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10393 ( .A0(T15201_Y), .BN(T7208_Y), .Y(T10393_Y),     .A1(T14684_Q));
KC_AOI21B_X2 T10392 ( .A0(T14684_Q), .BN(T10866_Y), .Y(T10392_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T8511 ( .A0(T4965_Y), .BN(T2282_Y), .Y(T8511_Y),     .A1(T1826_Q));
KC_AOI21B_X2 T10496 ( .A0(T15235_Y), .BN(T1652_Y), .Y(T10496_Y),     .A1(T14862_Q));
KC_AOI21B_X2 T10495 ( .A0(T15235_Y), .BN(T4908_Y), .Y(T10495_Y),     .A1(T14074_Q));
KC_AOI21B_X2 T10494 ( .A0(T14074_Q), .BN(T4907_Y), .Y(T10494_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T8492 ( .A0(T11491_Y), .BN(T5877_Y), .Y(T8492_Y),     .A1(T2791_Y));
KC_AOI21B_X2 T10490 ( .A0(T14050_Q), .BN(T5032_Y), .Y(T10490_Y),     .A1(T3054_Y));
KC_AOI21B_X2 T10489 ( .A0(T14855_Q), .BN(T5031_Y), .Y(T10489_Y),     .A1(T3054_Y));
KC_AOI21B_X2 T8486 ( .A0(T3297_Y), .BN(T12981_Y), .Y(T8486_Y),     .A1(T5062_Y));
KC_AOI21B_X2 T10435 ( .A0(T13648_Q), .BN(T5250_Y), .Y(T10435_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T10434 ( .A0(T13648_Q), .BN(T3594_Y), .Y(T10434_Y),     .A1(T15251_Y));
KC_AOI21B_X2 T16249 ( .A0(T14348_Q), .BN(T4320_Y), .Y(T16249_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10469 ( .A0(T15214_Y), .BN(T5137_Y), .Y(T10469_Y),     .A1(T14912_Q));
KC_AOI21B_X2 T10468 ( .A0(T14821_Q), .BN(T5138_Y), .Y(T10468_Y),     .A1(T15216_Y));
KC_AOI21B_X2 T10467 ( .A0(T15214_Y), .BN(T4219_Y), .Y(T10467_Y),     .A1(T14821_Q));
KC_AOI21B_X2 T10466 ( .A0(T15214_Y), .BN(T4222_Y), .Y(T10466_Y),     .A1(T14914_Q));
KC_AOI21B_X2 T8450 ( .A0(T3826_Y), .BN(T4382_Y), .Y(T8450_Y),     .A1(T3856_Y));
KC_AOI21B_X2 T10465 ( .A0(T13429_Q), .BN(T1858_Y), .Y(T10465_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T10382 ( .A0(T15244_Y), .BN(T10841_Y), .Y(T10382_Y),     .A1(T13352_Q));
KC_AOI21B_X2 T10452 ( .A0(T14796_Q), .BN(T5213_Y), .Y(T10452_Y),     .A1(T15212_Y));
KC_AOI21B_X2 T10451 ( .A0(T15251_Y), .BN(T5214_Y), .Y(T10451_Y),     .A1(T14796_Q));
KC_AOI21B_X2 T9630 ( .A0(T13689_Q), .BN(T10877_Y), .Y(T9630_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T9626 ( .A0(T13729_Q), .BN(T10649_Y), .Y(T9626_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T10341 ( .A0(T13866_Q), .BN(T10792_Y), .Y(T10341_Y),     .A1(T15207_Y));
KC_AOI21B_X2 T9718 ( .A0(T13806_Q), .BN(T7531_Y), .Y(T9718_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9794 ( .A0(T14635_Q), .BN(T10783_Y), .Y(T9794_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T9791 ( .A0(T13956_Q), .BN(T7720_Y), .Y(T9791_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T10191 ( .A0(T14899_Q), .BN(T4341_Y), .Y(T10191_Y),     .A1(T15217_Y));
KC_AOI21B_X2 T10146 ( .A0(T10743_Y), .BN(T1605_Y), .Y(T10146_Y),     .A1(T14378_Q));
KC_AOI21B_X2 T10135 ( .A0(T14592_Q), .BN(T1511_Y), .Y(T10135_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10134 ( .A0(T14380_Q), .BN(T1513_Y), .Y(T10134_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10132 ( .A0(T14372_Q), .BN(T4830_Y), .Y(T10132_Y),     .A1(T15224_Y));
KC_AOI21B_X2 T10498 ( .A0(T14862_Q), .BN(T1967_Y), .Y(T10498_Y),     .A1(T15246_Y));
KC_AOI21B_X2 T10396 ( .A0(T14722_Q), .BN(T7175_Y), .Y(T10396_Y),     .A1(T15205_Y));
KC_AOI21B_X2 T10332 ( .A0(T15235_Y), .BN(T10771_Y), .Y(T10332_Y),     .A1(T14635_Q));
KC_MXI2_X1 T8591 ( .Y(T8591_Y), .A(T6321_Y), .B(T9289_Y), .S0(T236_Y));
KC_MXI2_X1 T8886 ( .Y(T8886_Y), .A(T3926_Y), .B(T6358_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8884 ( .Y(T8884_Y), .A(T1617_Y), .B(T6364_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8883 ( .Y(T8883_Y), .A(T12331_Y), .B(T6415_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8882 ( .Y(T8882_Y), .A(T12344_Y), .B(T15313_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8881 ( .Y(T8881_Y), .A(T12125_Y), .B(T6430_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8879 ( .Y(T8879_Y), .A(T12112_Y), .B(T5349_Y),     .S0(T7919_Y));
KC_MXI2_X1 T8878 ( .Y(T8878_Y), .A(T12122_Y), .B(T6426_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8843 ( .Y(T8843_Y), .A(T619_Y), .B(T6411_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8842 ( .Y(T8842_Y), .A(T5418_Y), .B(T6357_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8841 ( .Y(T8841_Y), .A(T430_Y), .B(T6423_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8840 ( .Y(T8840_Y), .A(T12332_Y), .B(T6361_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8826 ( .Y(T8826_Y), .A(T617_Y), .B(T6401_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8824 ( .Y(T8824_Y), .A(T12190_Y), .B(T6730_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8823 ( .Y(T8823_Y), .A(T615_Y), .B(T6418_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8788 ( .Y(T8788_Y), .A(T12166_Y), .B(T6412_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8787 ( .Y(T8787_Y), .A(T5732_Y), .B(T16085_Q),     .S0(T16278_Y));
KC_MXI2_X1 T8786 ( .Y(T8786_Y), .A(T12443_Y), .B(T229_Y), .S0(T235_Q));
KC_MXI2_X1 T8990 ( .Y(T8990_Y), .A(T9203_Y), .B(T16287_Y),     .S0(T1339_Y));
KC_MXI2_X1 T8972 ( .Y(T8972_Y), .A(T12113_Y), .B(T2319_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8971 ( .Y(T8971_Y), .A(T12187_Y), .B(T6369_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8970 ( .Y(T8970_Y), .A(T10223_Y), .B(T6479_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8969 ( .Y(T8969_Y), .A(T12192_Y), .B(T6425_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8968 ( .Y(T8968_Y), .A(T12188_Y), .B(T6362_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8967 ( .Y(T8967_Y), .A(T1281_Y), .B(T6422_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8966 ( .Y(T8966_Y), .A(T618_Y), .B(T6379_Q), .S0(T7919_Y));
KC_MXI2_X1 T8959 ( .Y(T8959_Y), .A(T12120_Y), .B(T6391_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8958 ( .Y(T8958_Y), .A(T12133_Y), .B(T6432_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8956 ( .Y(T8956_Y), .A(T8924_Y), .B(T1245_Y),     .S0(T2312_Y));
KC_MXI2_X1 T8929 ( .Y(T8929_Y), .A(T1340_Y), .B(T8972_Y),     .S0(T8926_Y));
KC_MXI2_X1 T8928 ( .Y(T8928_Y), .A(T12323_Y), .B(T6683_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8927 ( .Y(T8927_Y), .A(T12121_Y), .B(T6424_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8926 ( .Y(T8926_Y), .A(T1742_Y), .B(T6416_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8925 ( .Y(T8925_Y), .A(T616_Y), .B(T6371_Q), .S0(T7919_Y));
KC_MXI2_X1 T8924 ( .Y(T8924_Y), .A(T10210_Y), .B(T6684_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8923 ( .Y(T8923_Y), .A(T1340_Y), .B(T8972_Y),     .S0(T8915_Y));
KC_MXI2_X1 T8922 ( .Y(T8922_Y), .A(T1245_Y), .B(T8924_Y),     .S0(T8092_Y));
KC_MXI2_X1 T9499 ( .Y(T9499_Y), .A(T5732_Y), .B(T9499_B),     .S0(T16281_Y));
KC_MXI2_X1 T9492 ( .Y(T9492_Y), .A(T12323_Y), .B(T9492_B),     .S0(T5299_Y));
KC_MXI2_X1 T9491 ( .Y(T9491_Y), .A(T615_Y), .B(T9491_B), .S0(T5299_Y));
KC_MXI2_X1 T9183 ( .Y(T9183_Y), .A(T12332_Y), .B(T9183_B),     .S0(T5299_Y));
KC_MXI2_X1 T9179 ( .Y(T9179_Y), .A(T12112_Y), .B(T9179_B),     .S0(T5299_Y));
KC_MXI2_X1 T9178 ( .Y(T9178_Y), .A(T4816_Y), .B(T9207_Y),     .S0(T8987_Y));
KC_MXI2_X1 T9134 ( .Y(T9134_Y), .A(T771_Q), .B(T9134_B), .S0(T5299_Y));
KC_MXI2_X1 T9133 ( .Y(T9133_Y), .A(T4801_Y), .B(T15091_Y),     .S0(T15092_Y));
KC_MXI2_X1 T9084 ( .Y(T9084_Y), .A(T1003_Q), .B(T9084_B),     .S0(T5299_Y));
KC_MXI2_X1 T9083 ( .Y(T9083_Y), .A(T772_Q), .B(T9083_B), .S0(T5299_Y));
KC_MXI2_X1 T9082 ( .Y(T9082_Y), .A(T1603_Y), .B(T9083_Y),     .S0(T9491_Y));
KC_MXI2_X1 T9250 ( .Y(T9250_Y), .A(T619_Y), .B(T9250_B),     .S0(T16281_Y));
KC_MXI2_X1 T9249 ( .Y(T9249_Y), .A(T1742_Y), .B(T9249_B),     .S0(T5299_Y));
KC_MXI2_X1 T9248 ( .Y(T9248_Y), .A(T12125_Y), .B(T9248_B),     .S0(T5299_Y));
KC_MXI2_X1 T9238 ( .Y(T9238_Y), .A(T12113_Y), .B(T9238_B),     .S0(T16281_Y));
KC_MXI2_X1 T9237 ( .Y(T9237_Y), .A(T12120_Y), .B(T9237_B),     .S0(T5299_Y));
KC_MXI2_X1 T9236 ( .Y(T9236_Y), .A(T10210_Y), .B(T9236_B),     .S0(T5299_Y));
KC_MXI2_X1 T9217 ( .Y(T9217_Y), .A(T616_Y), .B(T9217_B),     .S0(T16281_Y));
KC_MXI2_X1 T9216 ( .Y(T9216_Y), .A(T12122_Y), .B(T9216_B),     .S0(T5299_Y));
KC_MXI2_X1 T9215 ( .Y(T9215_Y), .A(T10223_Y), .B(T9215_B),     .S0(T5299_Y));
KC_MXI2_X1 T9214 ( .Y(T9214_Y), .A(T12187_Y), .B(T9214_B),     .S0(T5299_Y));
KC_MXI2_X1 T9213 ( .Y(T9213_Y), .A(T12192_Y), .B(T9213_B),     .S0(T5299_Y));
KC_MXI2_X1 T9212 ( .Y(T9212_Y), .A(T12133_Y), .B(T9212_B),     .S0(T5299_Y));
KC_MXI2_X1 T9211 ( .Y(T9211_Y), .A(T430_Y), .B(T9211_B),     .S0(T16281_Y));
KC_MXI2_X1 T9210 ( .Y(T9210_Y), .A(T617_Y), .B(T9210_B),     .S0(T16281_Y));
KC_MXI2_X1 T9209 ( .Y(T9209_Y), .A(T12190_Y), .B(T9209_B),     .S0(T16281_Y));
KC_MXI2_X1 T9208 ( .Y(T9208_Y), .A(T618_Y), .B(T9208_B),     .S0(T16281_Y));
KC_MXI2_X1 T9207 ( .Y(T9207_Y), .A(T12121_Y), .B(T9207_B),     .S0(T16281_Y));
KC_MXI2_X1 T9206 ( .Y(T9206_Y), .A(T10283_Y), .B(T9206_B),     .S0(T16281_Y));
KC_MXI2_X1 T9205 ( .Y(T9205_Y), .A(T1281_Y), .B(T9205_B),     .S0(T16281_Y));
KC_MXI2_X1 T9204 ( .Y(T9204_Y), .A(T12188_Y), .B(T9204_B),     .S0(T16281_Y));
KC_MXI2_X1 T9203 ( .Y(T9203_Y), .A(T5418_Y), .B(T9203_B),     .S0(T16281_Y));
KC_MXI2_X1 T9202 ( .Y(T9202_Y), .A(T3926_Y), .B(T9202_B),     .S0(T16281_Y));
KC_MXI2_X1 T9201 ( .Y(T9201_Y), .A(T12166_Y), .B(T9201_B),     .S0(T16281_Y));
KC_MXI2_X1 T8574 ( .Y(T8574_Y), .A(T273_Q), .B(T265_Y), .S0(T283_Q));
KC_MXI2_X1 T8627 ( .Y(T8627_Y), .A(T155_Q), .B(T6465_Y), .S0(T153_Q));
KC_MXI2_X1 T8626 ( .Y(T8626_Y), .A(T954_Y), .B(T160_Q), .S0(T348_Y));
KC_MXI2_X1 T8647 ( .Y(T8647_Y), .A(T15388_Y), .B(T170_Q), .S0(T397_Y));
KC_MXI2_X1 T8667 ( .Y(T8667_Y), .A(T360_Q), .B(T506_Y), .S0(T5278_Q));
KC_MXI2_X1 T8702 ( .Y(T8702_Y), .A(T16331_Y), .B(T16329_Y),     .S0(T7628_Y));
KC_MXI2_X1 T8701 ( .Y(T8701_Y), .A(T918_Y), .B(T16325_Y),     .S0(T7674_Y));
KC_MXI2_X1 T8700 ( .Y(T8700_Y), .A(T16331_Y), .B(T16329_Y),     .S0(T7578_Y));
KC_MXI2_X1 T8699 ( .Y(T8699_Y), .A(T9389_Y), .B(T7832_Y),     .S0(T7567_Y));
KC_MXI2_X1 T9422 ( .Y(T9422_Y), .A(T1334_Y), .B(T1272_Y),     .S0(T7863_Y));
KC_MXI2_X1 T8870 ( .Y(T8870_Y), .A(T8949_Y), .B(T8080_Y),     .S0(T7902_Y));
KC_MXI2_X1 T8779 ( .Y(T8779_Y), .A(T9398_Y), .B(T6944_Y), .S0(T235_Q));
KC_MXI2_X1 T8964 ( .Y(T8964_Y), .A(T1354_Y), .B(T9203_Y),     .S0(T8147_Y));
KC_MXI2_X1 T8915 ( .Y(T8915_Y), .A(T12191_Y), .B(T6363_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8914 ( .Y(T8914_Y), .A(T8948_Y), .B(T8099_Y),     .S0(T16391_Y));
KC_MXI2_X1 T8913 ( .Y(T8913_Y), .A(T8077_Y), .B(T8081_Y),     .S0(T7906_Y));
KC_MXI2_X1 T8912 ( .Y(T8912_Y), .A(T1266_Y), .B(T1286_Y),     .S0(T7904_Y));
KC_MXI2_X1 T8911 ( .Y(T8911_Y), .A(T1334_Y), .B(T1272_Y),     .S0(T7858_Y));
KC_MXI2_X1 T9483 ( .Y(T9483_Y), .A(T9484_Y), .B(T16191_Y),     .S0(T654_Y));
KC_MXI2_X1 T9198 ( .Y(T9198_Y), .A(T1617_Y), .B(T9198_B),     .S0(T16281_Y));
KC_MXI2_X1 T9197 ( .Y(T9197_Y), .A(T12344_Y), .B(T9197_B),     .S0(T16281_Y));
KC_MXI2_X1 T8572 ( .Y(T8572_Y), .A(T6313_Y), .B(T440_Q), .S0(T250_Y));
KC_MXI2_X1 T8749 ( .Y(T8749_Y), .A(T512_Q), .B(T913_Y), .S0(T530_Q));
KC_MXI2_X1 T9193 ( .Y(T9193_Y), .A(T567_Q), .B(T1599_Y), .S0(T1279_Y));
KC_MXI2_X1 T9279 ( .Y(T9279_Y), .A(T276_Q), .B(T310_Y), .S0(T628_Q));
KC_MXI2_X1 T8583 ( .Y(T8583_Y), .A(T15355_Y), .B(T5195_Q),     .S0(T15349_Y));
KC_MXI2_X1 T9311 ( .Y(T9311_Y), .A(T6638_Y), .B(T680_Q), .S0(T6700_Y));
KC_MXI2_X1 T8661 ( .Y(T8661_Y), .A(T695_Q), .B(T15406_Y),     .S0(T9340_Q));
KC_MXI2_X1 T8737 ( .Y(T8737_Y), .A(T701_Q), .B(T906_Y), .S0(T717_Q));
KC_MXI2_X1 T9415 ( .Y(T9415_Y), .A(T5385_Q), .B(T5387_Q),     .S0(T9446_Y));
KC_MXI2_X1 T9411 ( .Y(T9411_Y), .A(T5387_Q), .B(T5385_Q),     .S0(T15795_Q));
KC_MXI2_X1 T9409 ( .Y(T9409_Y), .A(T1153_Q), .B(T773_Y),     .S0(T15795_Q));
KC_MXI2_X1 T9408 ( .Y(T9408_Y), .A(T16232_Q), .B(T1152_Q),     .S0(T15795_Q));
KC_MXI2_X1 T9407 ( .Y(T9407_Y), .A(T761_Q), .B(T767_Q), .S0(T9446_Y));
KC_MXI2_X1 T8853 ( .Y(T8853_Y), .A(T963_Q), .B(T759_Y), .S0(T15795_Q));
KC_MXI2_X1 T8852 ( .Y(T8852_Y), .A(T963_Q), .B(T759_Y), .S0(T15795_Q));
KC_MXI2_X1 T8851 ( .Y(T8851_Y), .A(T999_Q), .B(T4844_Y),     .S0(T15795_Q));
KC_MXI2_X1 T8803 ( .Y(T8803_Y), .A(T767_Q), .B(T761_Q), .S0(T15795_Q));
KC_MXI2_X1 T8802 ( .Y(T8802_Y), .A(T1160_Q), .B(T9459_Q),     .S0(T15795_Q));
KC_MXI2_X1 T9010 ( .Y(T9010_Y), .A(T1000_Q), .B(T995_Q), .S0(T9446_Y));
KC_MXI2_X1 T9001 ( .Y(T9001_Y), .A(T995_Q), .B(T1000_Q),     .S0(T15795_Q));
KC_MXI2_X1 T8942 ( .Y(T8942_Y), .A(T983_Q), .B(T978_Q), .S0(T9446_Y));
KC_MXI2_X1 T8939 ( .Y(T8939_Y), .A(T978_Q), .B(T983_Q), .S0(T15795_Q));
KC_MXI2_X1 T8899 ( .Y(T8899_Y), .A(T760_Q), .B(T765_Q), .S0(T9446_Y));
KC_MXI2_X1 T8898 ( .Y(T8898_Y), .A(T762_Q), .B(T768_Q), .S0(T9446_Y));
KC_MXI2_X1 T8895 ( .Y(T8895_Y), .A(T765_Q), .B(T760_Q), .S0(T15795_Q));
KC_MXI2_X1 T8894 ( .Y(T8894_Y), .A(T768_Q), .B(T762_Q), .S0(T15795_Q));
KC_MXI2_X1 T8893 ( .Y(T8893_Y), .A(T1159_Q), .B(T9458_Q),     .S0(T15795_Q));
KC_MXI2_X1 T9240 ( .Y(T9240_Y), .A(T15658_Y), .B(T781_Q),     .S0(T9464_Y));
KC_MXI2_X1 T9273 ( .Y(T9273_Y), .A(T6257_Y), .B(T825_Q), .S0(T244_Y));
KC_MXI2_X1 T9256 ( .Y(T9256_Y), .A(T377_Y), .B(T671_Q), .S0(T15387_Y));
KC_MXI2_X1 T9412 ( .Y(T9412_Y), .A(T1151_Q), .B(T985_Y),     .S0(T15795_Q));
KC_MXI2_X1 T8801 ( .Y(T8801_Y), .A(T12445_Y), .B(T7838_Y),     .S0(T926_Y));
KC_MXI2_X1 T8995 ( .Y(T8995_Y), .A(T982_Q), .B(T976_Q), .S0(T8060_Y));
KC_MXI2_X1 T9222 ( .Y(T9222_Y), .A(T2719_Y), .B(T16301_Q),     .S0(T10260_Y));
KC_MXI2_X1 T9221 ( .Y(T9221_Y), .A(T2719_Y), .B(T16301_Q),     .S0(T10262_Y));
KC_MXI2_X1 T9219 ( .Y(T9219_Y), .A(T15912_Y), .B(T5380_Q),     .S0(T10534_Y));
KC_MXI2_X1 T9186 ( .Y(T9186_Y), .A(T15912_Y), .B(T5380_Q),     .S0(T1021_Y));
KC_MXI2_X1 T9184 ( .Y(T9184_Y), .A(T15855_Y), .B(T15796_Q),     .S0(T1020_Y));
KC_MXI2_X1 T9817 ( .Y(T9817_Y), .A(T7385_Y), .B(T1071_Q),     .S0(T8026_Y));
KC_MXI2_X1 T9814 ( .Y(T9814_Y), .A(T7385_Y), .B(T1073_Q),     .S0(T8028_Y));
KC_MXI2_X1 T9813 ( .Y(T9813_Y), .A(T15722_Y), .B(T1064_Q),     .S0(T8028_Y));
KC_MXI2_X1 T9783 ( .Y(T9783_Y), .A(T15722_Y), .B(T1061_Q),     .S0(T8026_Y));
KC_MXI2_X1 T9928 ( .Y(T9928_Y), .A(T15722_Y), .B(T8834_Q),     .S0(T7978_Y));
KC_MXI2_X1 T9927 ( .Y(T9927_Y), .A(T15722_Y), .B(T1121_Q),     .S0(T8027_Y));
KC_MXI2_X1 T9916 ( .Y(T9916_Y), .A(T9919_Y), .B(T9918_Y),     .S0(T1209_Q));
KC_MXI2_X1 T9358 ( .Y(T9358_Y), .A(T7385_Y), .B(T1122_Q),     .S0(T7978_Y));
KC_MXI2_X1 T9984 ( .Y(T9984_Y), .A(T16275_Y), .B(T10942_Y),     .S0(T5376_Q));
KC_MXI2_X1 T10237 ( .Y(T10237_Y), .A(T2127_Y), .B(T15798_Q),     .S0(T1005_Q));
KC_MXI2_X1 T10236 ( .Y(T10236_Y), .A(T15882_Y), .B(T964_Q),     .S0(T1018_Y));
KC_MXI2_X1 T10235 ( .Y(T10235_Y), .A(T16474_Y), .B(T15005_Y),     .S0(T1161_Y));
KC_MXI2_X1 T10234 ( .Y(T10234_Y), .A(T15857_Y), .B(T16088_Q),     .S0(T1173_Y));
KC_MXI2_X1 T10232 ( .Y(T10232_Y), .A(T15853_Y), .B(T15844_Q),     .S0(T1178_Y));
KC_MXI2_X1 T10231 ( .Y(T10231_Y), .A(T15856_Y), .B(T15808_Q),     .S0(T1175_Y));
KC_MXI2_X1 T10230 ( .Y(T10230_Y), .A(T15854_Y), .B(T16299_Q),     .S0(T1171_Y));
KC_MXI2_X1 T10222 ( .Y(T10222_Y), .A(T15881_Y), .B(T15797_Q),     .S0(T994_Y));
KC_MXI2_X1 T10221 ( .Y(T10221_Y), .A(T15857_Y), .B(T16088_Q),     .S0(T15327_Y));
KC_MXI2_X1 T10220 ( .Y(T10220_Y), .A(T15881_Y), .B(T15797_Q),     .S0(T1017_Y));
KC_MXI2_X1 T10219 ( .Y(T10219_Y), .A(T1748_Y), .B(T15805_Q),     .S0(T1157_Q));
KC_MXI2_X1 T10216 ( .Y(T10216_Y), .A(T1748_Y), .B(T15805_Q),     .S0(T1177_Y));
KC_MXI2_X1 T10215 ( .Y(T10215_Y), .A(T15853_Y), .B(T15844_Q),     .S0(T5384_Q));
KC_MXI2_X1 T10214 ( .Y(T10214_Y), .A(T2751_Y), .B(T15807_Q),     .S0(T1251_Y));
KC_MXI2_X1 T10213 ( .Y(T10213_Y), .A(T2751_Y), .B(T15807_Q),     .S0(T1146_Y));
KC_MXI2_X1 T10212 ( .Y(T10212_Y), .A(T15856_Y), .B(T15808_Q),     .S0(T1172_Y));
KC_MXI2_X1 T10208 ( .Y(T10208_Y), .A(T15858_Y), .B(T15809_Q),     .S0(T1269_Y));
KC_MXI2_X1 T9220 ( .Y(T9220_Y), .A(T16474_Y), .B(T15005_Y),     .S0(T1019_Y));
KC_MXI2_X1 T9185 ( .Y(T9185_Y), .A(T15882_Y), .B(T964_Q),     .S0(T1014_Y));
KC_MXI2_X1 T10286 ( .Y(T10286_Y), .A(T10245_Y), .B(T15804_Q),     .S0(T1267_Y));
KC_MXI2_X1 T10153 ( .Y(T10153_Y), .A(T15529_Y), .B(T13121_Y),     .S0(T1250_Q));
KC_MXI2_X1 T10141 ( .Y(T10141_Y), .A(T1365_Y), .B(T13125_Y),     .S0(T1265_Q));
KC_MXI2_X1 T10137 ( .Y(T10137_Y), .A(T1362_Y), .B(T10936_Y),     .S0(T1264_Q));
KC_MXI2_X1 T10136 ( .Y(T10136_Y), .A(T1366_Y), .B(T10934_Y),     .S0(T1271_Q));
KC_MXI2_X1 T10124 ( .Y(T10124_Y), .A(T10245_Y), .B(T15804_Q),     .S0(T4862_Q));
KC_MXI2_X1 T10218 ( .Y(T10218_Y), .A(T5382_Y), .B(T13056_Q),     .S0(T1275_Y));
KC_MXI2_X1 T10217 ( .Y(T10217_Y), .A(T15895_Y), .B(T15803_Q),     .S0(T16506_Y));
KC_MXI2_X1 T10123 ( .Y(T10123_Y), .A(T15527_Y), .B(T4825_Y),     .S0(T10285_Y));
KC_MXI2_X1 T9785 ( .Y(T9785_Y), .A(T809_Y), .B(T1661_Q), .S0(T1660_Q));
KC_MXI2_X1 T10531 ( .Y(T10531_Y), .A(T16372_Y), .B(T1717_Q),     .S0(T8880_Q));
KC_MXI2_X1 T10530 ( .Y(T10530_Y), .A(T1192_Y), .B(T1707_Q),     .S0(T1719_Q));
KC_MXI2_X1 T10529 ( .Y(T10529_Y), .A(T16374_Y), .B(T8877_Q),     .S0(T10530_Y));
KC_MXI2_X1 T9977 ( .Y(T9977_Y), .A(T1148_Y), .B(T16433_Q),     .S0(T5364_Q));
KC_MXI2_X1 T9976 ( .Y(T9976_Y), .A(T1148_Y), .B(T16433_Q),     .S0(T2012_Q));
KC_MXI2_X1 T10086 ( .Y(T10086_Y), .A(T1519_Y), .B(T1735_Q),     .S0(T5362_Q));
KC_MXI2_X1 T10070 ( .Y(T10070_Y), .A(T16373_Y), .B(T1691_Q),     .S0(T16413_Q));
KC_MXI2_X1 T10068 ( .Y(T10068_Y), .A(T16372_Y), .B(T1717_Q),     .S0(T5391_Q));
KC_MXI2_X1 T10067 ( .Y(T10067_Y), .A(T16373_Y), .B(T1691_Q),     .S0(T1736_Q));
KC_MXI2_X1 T10066 ( .Y(T10066_Y), .A(T1192_Y), .B(T1707_Q),     .S0(T2002_Q));
KC_MXI2_X1 T8253 ( .Y(T8253_Y), .A(T1766_Y), .B(T8251_Y),     .S0(T11530_Y));
KC_MXI2_X1 T10521 ( .Y(T10521_Y), .A(T2015_Q), .B(T16378_Y),     .S0(T5434_Q));
KC_MXI2_X1 T10515 ( .Y(T10515_Y), .A(T2023_Q), .B(T15478_Y),     .S0(T4971_Q));
KC_MXI2_X1 T9966 ( .Y(T9966_Y), .A(T2016_Q), .B(T1116_Y),     .S0(T2115_Q));
KC_MXI2_X1 T9958 ( .Y(T9958_Y), .A(T2024_Y), .B(T11259_Y),     .S0(T1162_Y));
KC_MXI2_X1 T9941 ( .Y(T9941_Y), .A(T9958_Y), .B(T2020_Y),     .S0(T9940_Y));
KC_MXI2_X1 T9940 ( .Y(T9940_Y), .A(T1998_Y), .B(T2020_Y),     .S0(T2024_Y));
KC_MXI2_X1 T10120 ( .Y(T10120_Y), .A(T2053_Q), .B(T1517_Y),     .S0(T4969_Q));
KC_MXI2_X1 T10113 ( .Y(T10113_Y), .A(T5397_Q), .B(T16269_Y),     .S0(T2692_Q));
KC_MXI2_X1 T10112 ( .Y(T10112_Y), .A(T2002_Q), .B(T15511_Y),     .S0(T5432_Q));
KC_MXI2_X1 T10111 ( .Y(T10111_Y), .A(T2012_Q), .B(T1532_Y),     .S0(T5438_Q));
KC_MXI2_X1 T10110 ( .Y(T10110_Y), .A(T5391_Q), .B(T1533_Y),     .S0(T5442_Q));
KC_MXI2_X1 T10109 ( .Y(T10109_Y), .A(T1736_Q), .B(T15512_Y),     .S0(T5429_Q));
KC_MXI2_X1 T10108 ( .Y(T10108_Y), .A(T1735_Q), .B(T1519_Y),     .S0(T2095_Q));
KC_MXI2_X1 T10107 ( .Y(T10107_Y), .A(T1533_Y), .B(T5391_Q),     .S0(T5390_Q));
KC_MXI2_X1 T10106 ( .Y(T10106_Y), .A(T15511_Y), .B(T2002_Q),     .S0(T2053_Q));
KC_MXI2_X1 T10092 ( .Y(T10092_Y), .A(T16269_Y), .B(T5397_Q),     .S0(T10082_Y));
KC_MXI2_X1 T10088 ( .Y(T10088_Y), .A(T4425_Y), .B(T2627_Q),     .S0(T16411_Y));
KC_MXI2_X1 T10082 ( .Y(T10082_Y), .A(T1532_Y), .B(T2012_Q),     .S0(T1736_Q));
KC_MXI2_X1 T10063 ( .Y(T10063_Y), .A(T16269_Y), .B(T5397_Q),     .S0(T5364_Q));
KC_MXI2_X1 T8199 ( .Y(T8199_Y), .A(T6097_Co), .B(T2121_Y),     .S0(T2100_Y));
KC_MXI2_X1 T8497 ( .Y(T8497_Y), .A(T11436_Y), .B(T2152_Q),     .S0(T8316_Y));
KC_MXI2_X1 T8240 ( .Y(T8240_Y), .A(T5927_Y), .B(T15138_Q),     .S0(T15005_Y));
KC_MXI2_X1 T8296 ( .Y(T8296_Y), .A(T5991_Y), .B(T2275_Q),     .S0(T16076_Y));
KC_MXI2_X1 T8282 ( .Y(T8282_Y), .A(T6028_Y), .B(T2316_Q),     .S0(T15796_Q));
KC_MXI2_X1 T8341 ( .Y(T8341_Y), .A(T4968_Y), .B(T16082_Q),     .S0(T15797_Q));
KC_MXI2_X1 T8340 ( .Y(T8340_Y), .A(T2239_Y), .B(T2237_Q),     .S0(T16235_Y));
KC_MXI2_X1 T8328 ( .Y(T8328_Y), .A(T2247_Y), .B(T2314_Q),     .S0(T15844_Q));
KC_MXI2_X1 T8327 ( .Y(T8327_Y), .A(T2240_Y), .B(T4964_Q),     .S0(T16301_Q));
KC_MXI2_X1 T8319 ( .Y(T8319_Y), .A(T2246_Y), .B(T5486_Q),     .S0(T15807_Q));
KC_MXI2_X1 T8310 ( .Y(T8310_Y), .A(T2250_Y), .B(T2313_Q),     .S0(T15808_Q));
KC_MXI2_X1 T8309 ( .Y(T8309_Y), .A(T1788_Y), .B(T2311_Q),     .S0(T15809_Q));
KC_MXI2_X1 T8374 ( .Y(T8374_Y), .A(T16082_Q), .B(T4968_Y),     .S0(T8352_Q));
KC_MXI2_X1 T8363 ( .Y(T8363_Y), .A(T16041_Y), .B(T2278_Q),     .S0(T2264_Y));
KC_MXI2_X1 T8353 ( .Y(T8353_Y), .A(T2279_Y), .B(T6419_Q),     .S0(T16299_Q));
KC_MXI2_X1 T8347 ( .Y(T8347_Y), .A(T2245_Y), .B(T5494_Q),     .S0(T15805_Q));
KC_MXI2_X1 T8402 ( .Y(T8402_Y), .A(T2279_Y), .B(T6419_Q),     .S0(T10627_Y));
KC_MXI2_X1 T8400 ( .Y(T8400_Y), .A(T2247_Y), .B(T2314_Q),     .S0(T10597_Y));
KC_MXI2_X1 T8388 ( .Y(T8388_Y), .A(T2240_Y), .B(T4964_Q),     .S0(T10626_Y));
KC_MXI2_X1 T8414 ( .Y(T8414_Y), .A(T5527_Q), .B(T1833_Q),     .S0(T2353_Q));
KC_MXI2_X1 T8413 ( .Y(T8413_Y), .A(T2364_Q), .B(T1832_Q),     .S0(T2353_Q));
KC_MXI2_X1 T8412 ( .Y(T8412_Y), .A(T8411_Y), .B(T8404_Y),     .S0(T1830_Q));
KC_MXI2_X1 T8411 ( .Y(T8411_Y), .A(T8413_Y), .B(T8414_Y),     .S0(T5526_Q));
KC_MXI2_X1 T8404 ( .Y(T8404_Y), .A(T8427_Y), .B(T8428_Y),     .S0(T5526_Q));
KC_MXI2_X1 T8428 ( .Y(T8428_Y), .A(T1857_Q), .B(T2388_Q),     .S0(T2353_Q));
KC_MXI2_X1 T8427 ( .Y(T8427_Y), .A(T5529_Q), .B(T1856_Q),     .S0(T2353_Q));
KC_MXI2_X1 T9652 ( .Y(T9652_Y), .A(T13769_Q), .B(T418_Y),     .S0(T12559_Y));
KC_MXI2_X1 T9638 ( .Y(T9638_Y), .A(T14766_Q), .B(T404_Y),     .S0(T3018_Y));
KC_MXI2_X1 T8524 ( .Y(T8524_Y), .A(T14928_Q), .B(T411_Y),     .S0(T2446_Y));
KC_MXI2_X1 T9774 ( .Y(T9774_Y), .A(T633_Y), .B(T2466_Y),     .S0(T10475_Y));
KC_MXI2_X1 T9877 ( .Y(T9877_Y), .A(T859_Y), .B(T14032_Q),     .S0(T3099_Y));
KC_MXI2_X1 T9838 ( .Y(T9838_Y), .A(T9743_Y), .B(T16404_Y),     .S0(T9877_Y));
KC_MXI2_X1 T9948 ( .Y(T9948_Y), .A(T1141_Y), .B(T2591_Q),     .S0(T2592_Q));
KC_MXI2_X1 T9938 ( .Y(T9938_Y), .A(T14884_Q), .B(T16405_Y),     .S0(T2568_Y));
KC_MXI2_X1 T10118 ( .Y(T10118_Y), .A(T14367_Q), .B(T1546_Y),     .S0(T2556_Y));
KC_MXI2_X1 T10089 ( .Y(T10089_Y), .A(T1499_Y), .B(T10103_Y),     .S0(T2610_Y));
KC_MXI2_X1 T10269 ( .Y(T10269_Y), .A(T10271_Y), .B(T10244_Y),     .S0(T14954_Q));
KC_MXI2_X1 T8441 ( .Y(T8441_Y), .A(T14954_Q), .B(T5766_Y),     .S0(T11342_Y));
KC_MXI2_X1 T8496 ( .Y(T8496_Y), .A(T15805_Q), .B(T1748_Y),     .S0(T5462_Q));
KC_MXI2_X1 T8495 ( .Y(T8495_Y), .A(T15005_Y), .B(T16474_Y),     .S0(T12980_Q));
KC_MXI2_X1 T8234 ( .Y(T8234_Y), .A(T2127_Y), .B(T15798_Q),     .S0(T13104_Q));
KC_MXI2_X1 T8233 ( .Y(T8233_Y), .A(T15804_Q), .B(T10245_Y),     .S0(T13119_Q));
KC_MXI2_X1 T8232 ( .Y(T8232_Y), .A(T16299_Q), .B(T15854_Y),     .S0(T13096_Q));
KC_MXI2_X1 T8227 ( .Y(T8227_Y), .A(T16088_Q), .B(T15857_Y),     .S0(T3970_Q));
KC_MXI2_X1 T8226 ( .Y(T8226_Y), .A(T964_Q), .B(T15882_Y),     .S0(T13103_Q));
KC_MXI2_X1 T8225 ( .Y(T8225_Y), .A(T16301_Q), .B(T2719_Y),     .S0(T13316_Q));
KC_MXI2_X1 T8218 ( .Y(T8218_Y), .A(T15808_Q), .B(T15856_Y),     .S0(T13298_Q));
KC_MXI2_X1 T8217 ( .Y(T8217_Y), .A(T15809_Q), .B(T15858_Y),     .S0(T13299_Q));
KC_MXI2_X1 T8216 ( .Y(T8216_Y), .A(T15803_Q), .B(T15895_Y),     .S0(T3257_Q));
KC_MXI2_X1 T8211 ( .Y(T8211_Y), .A(T15566_Y), .B(T2163_Y),     .S0(T13106_Y));
KC_MXI2_X1 T8209 ( .Y(T8209_Y), .A(T15796_Q), .B(T15855_Y),     .S0(T5451_Q));
KC_MXI2_X1 T8207 ( .Y(T8207_Y), .A(T15844_Q), .B(T15853_Y),     .S0(T13297_Q));
KC_MXI2_X1 T8248 ( .Y(T8248_Y), .A(T15797_Q), .B(T15881_Y),     .S0(T3971_Q));
KC_MXI2_X1 T8339 ( .Y(T8339_Y), .A(T15912_Y), .B(T5380_Q),     .S0(T2345_Q));
KC_MXI2_X1 T8338 ( .Y(T8338_Y), .A(T2811_Y), .B(T13139_Y),     .S0(T2782_Y));
KC_MXI2_X1 T8335 ( .Y(T8335_Y), .A(T11651_Y), .B(T10954_Y),     .S0(T3294_Y));
KC_MXI2_X1 T8315 ( .Y(T8315_Y), .A(T16017_Y), .B(T8352_Q),     .S0(T16088_Q));
KC_MXI2_X1 T8308 ( .Y(T8308_Y), .A(T6055_Y), .B(T2843_Q),     .S0(T9162_Y));
KC_MXI2_X1 T8509 ( .Y(T8509_Y), .A(T4748_Y), .B(T16101_Y),     .S0(T16088_Q));
KC_MXI2_X1 T8351 ( .Y(T8351_Y), .A(T5497_Q), .B(T2280_Y),     .S0(T15804_Q));
KC_MXI2_X1 T8387 ( .Y(T8387_Y), .A(T6183_Y), .B(T2873_Y),     .S0(T11699_Y));
KC_MXI2_X1 T8422 ( .Y(T8422_Y), .A(T12105_Y), .B(T16131_Y),     .S0(T4999_Y));
KC_MXI2_X1 T8408 ( .Y(T8408_Y), .A(T12103_Y), .B(T16130_Y),     .S0(T2898_Y));
KC_MXI2_X1 T8407 ( .Y(T8407_Y), .A(T6222_Y), .B(T12106_Y),     .S0(T11771_Y));
KC_MXI2_X1 T8403 ( .Y(T8403_Y), .A(T12107_Y), .B(T6225_Y),     .S0(T11770_Y));
KC_MXI2_X1 T8152 ( .Y(T8152_Y), .A(T5536_Q), .B(T6509_Y),     .S0(T2932_Y));
KC_MXI2_X1 T9666 ( .Y(T9666_Y), .A(T13767_Q), .B(T15403_Y),     .S0(T12556_Y));
KC_MXI2_X1 T9663 ( .Y(T9663_Y), .A(T13781_Q), .B(T483_Y),     .S0(T3017_Y));
KC_MXI2_X1 T8523 ( .Y(T8523_Y), .A(T14931_Q), .B(T6761_Y),     .S0(T3015_Y));
KC_MXI2_X1 T9837 ( .Y(T9837_Y), .A(T14082_Q), .B(T872_Y),     .S0(T5288_Y));
KC_MXI2_X1 T8224 ( .Y(T8224_Y), .A(T11460_Y), .B(T3269_Y),     .S0(T6163_Y));
KC_MXI2_X1 T8208 ( .Y(T8208_Y), .A(T2753_Y), .B(T2730_Y),     .S0(T10201_Y));
KC_MXI2_X1 T8266 ( .Y(T8266_Y), .A(T6230_S), .B(T12210_Y),     .S0(T6230_Co));
KC_MXI2_X1 T8322 ( .Y(T8322_Y), .A(T3340_Y), .B(T3353_Y),     .S0(T3346_Y));
KC_MXI2_X1 T8361 ( .Y(T8361_Y), .A(T2841_Q), .B(T15802_Q),     .S0(T11646_Y));
KC_MXI2_X1 T8431 ( .Y(T8431_Y), .A(T15640_Y), .B(T4164_Q),     .S0(T11813_Y));
KC_MXI2_X1 T8440 ( .Y(T8440_Y), .A(T15546_Y), .B(T5760_Y),     .S0(T15835_Y));
KC_MXI2_X1 T8179 ( .Y(T8179_Y), .A(T11345_Y), .B(T3821_Y),     .S0(T4465_Q));
KC_MXI2_X1 T8188 ( .Y(T8188_Y), .A(T12167_Y), .B(T12181_Y),     .S0(T16153_Y));
KC_MXI2_X1 T8229 ( .Y(T8229_Y), .A(T3861_Y), .B(T12807_Y),     .S0(T3884_Q));
KC_MXI2_X1 T8222 ( .Y(T8222_Y), .A(T10926_Y), .B(T10633_Y),     .S0(T3889_Q));
KC_MXI2_X1 T8213 ( .Y(T8213_Y), .A(T14551_Q), .B(T5852_Y),     .S0(T11433_Y));
KC_MXI2_X1 T8256 ( .Y(T8256_Y), .A(T3916_Y), .B(T13115_Y),     .S0(T3936_Q));
KC_MXI2_X1 T8255 ( .Y(T8255_Y), .A(T3905_Y), .B(T5892_Y),     .S0(T12204_Y));
KC_MXI2_X1 T8237 ( .Y(T8237_Y), .A(T15971_Y), .B(T4968_Y),     .S0(T10937_Y));
KC_MXI2_X1 T8477 ( .Y(T8477_Y), .A(T5956_Y), .B(T12243_Y),     .S0(T11614_Y));
KC_MXI2_X1 T8289 ( .Y(T8289_Y), .A(T5972_Y), .B(T3970_Q),     .S0(T3971_Q));
KC_MXI2_X1 T8505 ( .Y(T8505_Y), .A(T4748_Y), .B(T12035_Y),     .S0(T11717_Y));
KC_MXI2_X1 T8504 ( .Y(T8504_Y), .A(T6077_Y), .B(T8507_Y),     .S0(T5055_Y));
KC_MXI2_X1 T8372 ( .Y(T8372_Y), .A(T5466_Y), .B(T6077_Y),     .S0(T15797_Q));
KC_MXI2_X1 T8371 ( .Y(T8371_Y), .A(T5525_Q), .B(T6048_Y),     .S0(T5528_Q));
KC_MXI2_X1 T8360 ( .Y(T8360_Y), .A(T6555_Q), .B(T16035_Y),     .S0(T5532_Q));
KC_MXI2_X1 T8359 ( .Y(T8359_Y), .A(T4046_Y), .B(T16108_Y),     .S0(T15005_Y));
KC_MXI2_X1 T8357 ( .Y(T8357_Y), .A(T15760_Q), .B(T6044_Y),     .S0(T4171_Q));
KC_MXI2_X1 T8356 ( .Y(T8356_Y), .A(T6526_Q), .B(T5070_Y),     .S0(T4178_Q));
KC_MXI2_X1 T8399 ( .Y(T8399_Y), .A(T6170_Y), .B(T12288_Y),     .S0(T4067_Y));
KC_MXI2_X1 T8392 ( .Y(T8392_Y), .A(T4716_Y), .B(T5504_Y),     .S0(T12281_Y));
KC_MXI2_X1 T8391 ( .Y(T8391_Y), .A(T5510_Y), .B(T6137_Y), .S0(T964_Q));
KC_MXI2_X1 T8514 ( .Y(T8514_Y), .A(T4147_Q), .B(T6175_Y),     .S0(T4163_Q));
KC_MXI2_X1 T8513 ( .Y(T8513_Y), .A(T6156_Y), .B(T11794_Y),     .S0(T12966_Y));
KC_MXI2_X1 T8512 ( .Y(T8512_Y), .A(T5530_Q), .B(T6034_Y),     .S0(T4164_Q));
KC_MXI2_X1 T8421 ( .Y(T8421_Y), .A(T6587_Y), .B(T11793_Y),     .S0(T5111_Y));
KC_MXI2_X1 T8164 ( .Y(T8164_Y), .A(T6079_Y), .B(T12866_Y),     .S0(T3437_Y));
KC_MXI2_X1 T8430 ( .Y(T8430_Y), .A(T6517_Y), .B(T4168_Q),     .S0(T11001_Y));
KC_MXI2_X1 T8429 ( .Y(T8429_Y), .A(T6524_Y), .B(T4169_Q),     .S0(T11830_Y));
KC_MXI2_X1 T8425 ( .Y(T8425_Y), .A(T4171_Q), .B(T6527_Y),     .S0(T5533_Y));
KC_MXI2_X1 T8184 ( .Y(T8184_Y), .A(T14523_Q), .B(T15557_Y),     .S0(T14943_Q));
KC_MXI2_X1 T8202 ( .Y(T8202_Y), .A(T3831_Y), .B(T4394_Y),     .S0(T5553_Y));
KC_MXI2_X1 T8442 ( .Y(T8442_Y), .A(T14548_Q), .B(T14551_Q),     .S0(T4463_Y));
KC_MXI2_X1 T8501 ( .Y(T8501_Y), .A(T5499_Q), .B(T6075_Y),     .S0(T4773_Y));
KC_MXI2_X1 T8500 ( .Y(T8500_Y), .A(T4669_Q), .B(T16111_Y),     .S0(T4775_Y));
KC_MXI2_X1 T8499 ( .Y(T8499_Y), .A(T5498_Q), .B(T6076_Y),     .S0(T4764_Y));
KC_MXI2_X1 T8462 ( .Y(T8462_Y), .A(T6103_Y), .B(T16460_Q),     .S0(T4629_Q));
KC_MXI2_X1 T8461 ( .Y(T8461_Y), .A(T6103_Y), .B(T16460_Q),     .S0(T5162_Q));
KC_MXI2_X1 T8460 ( .Y(T8460_Y), .A(T6103_Y), .B(T16460_Q),     .S0(T5488_Q));
KC_MXI2_X1 T8366 ( .Y(T8366_Y), .A(T6029_Y), .B(T4661_Y),     .S0(T4668_Y));
KC_MXI2_X1 T8344 ( .Y(T8344_Y), .A(T16460_Q), .B(T6103_Y),     .S0(T4627_Q));
KC_MXI2_X1 T8379 ( .Y(T8379_Y), .A(T6104_Y), .B(T4735_Y),     .S0(T4703_Y));
KC_MXI2_X1 T8406 ( .Y(T8406_Y), .A(T6420_S), .B(T11758_Y),     .S0(T6187_Y));
KC_MXI2_X1 T9496 ( .Y(T9496_Y), .A(T9471_Q), .B(T9496_B),     .S0(T5299_Y));
KC_MXI2_X1 T9495 ( .Y(T9495_Y), .A(T5416_Q), .B(T9495_B),     .S0(T5299_Y));
KC_MXI2_X1 T9494 ( .Y(T9494_Y), .A(T9470_Q), .B(T9494_B),     .S0(T5299_Y));
KC_MXI2_X1 T9493 ( .Y(T9493_Y), .A(T12331_Y), .B(T9493_B),     .S0(T5299_Y));
KC_MXI2_X1 T9451 ( .Y(T9451_Y), .A(T9084_Y), .B(T16283_Y),     .S0(T9236_Y));
KC_MXI2_X1 T9484 ( .Y(T9484_Y), .A(T769_Q), .B(T9484_B),     .S0(T16281_Y));
KC_MXI2_X1 T9377 ( .Y(T9377_Y), .A(T9375_Y), .B(T7824_Y),     .S0(T7688_Y));
KC_MXI2_X1 T9376 ( .Y(T9376_Y), .A(T9384_Y), .B(T7822_Y),     .S0(T7569_Y));
KC_MXI2_X1 T9445 ( .Y(T9445_Y), .A(T9457_Q), .B(T997_Q), .S0(T9446_Y));
KC_MXI2_X1 T9357 ( .Y(T9357_Y), .A(T7385_Y), .B(T1078_Q),     .S0(T8027_Y));
KC_MXI2_X1 T10287 ( .Y(T10287_Y), .A(T15895_Y), .B(T15803_Q),     .S0(T1155_Y));
KC_MXI2_X1 T10532 ( .Y(T10532_Y), .A(T16374_Y), .B(T8877_Q),     .S0(T1735_Q));
KC_MXI2_X1 T16291 ( .Y(T16291_Y), .A(T5390_Q), .B(T15519_Y),     .S0(T4970_Q));
KC_MXI2_X1 T10522 ( .Y(T10522_Y), .A(T16269_Y), .B(T5397_Q),     .S0(T10520_Y));
KC_MXI2_X1 T8473 ( .Y(T8473_Y), .A(T16041_Y), .B(T2278_Q),     .S0(T964_Q));
KC_MXI2_X1 T8471 ( .Y(T8471_Y), .A(T6040_Y), .B(T5481_Q),     .S0(T16073_Y));
KC_MXI2_X1 T8470 ( .Y(T8470_Y), .A(T16042_Y), .B(T5571_Q),     .S0(T15798_Q));
KC_MXI2_X1 T10540 ( .Y(T10540_Y), .A(T13063_Q), .B(T13291_Q),     .S0(T2669_Q));
KC_MXI2_X1 T8484 ( .Y(T8484_Y), .A(T6383_Y), .B(T3977_Y),     .S0(T3294_Y));
KC_MXI2_X1 T8472 ( .Y(T8472_Y), .A(T5008_Y), .B(T2854_Y),     .S0(T2815_Q));
KC_MXI2_X1 T8482 ( .Y(T8482_Y), .A(T3391_Y), .B(T10955_Y),     .S0(T3294_Y));
KC_MXI2_X1 T8506 ( .Y(T8506_Y), .A(T5135_Y), .B(T6157_Y),     .S0(T5380_Q));
KC_MXI2_X1 T8165 ( .Y(T8165_Y), .A(T3996_Y), .B(T6525_Y),     .S0(T12318_Y));
KC_MXI2_X1 T8459 ( .Y(T8459_Y), .A(T6103_Y), .B(T16460_Q),     .S0(T4630_Q));
KC_MXI2_X1 T8458 ( .Y(T8458_Y), .A(T6103_Y), .B(T16460_Q),     .S0(T4628_Q));
KC_MXI2_X1 T8457 ( .Y(T8457_Y), .A(T16460_Q), .B(T6103_Y),     .S0(T4626_Q));
KC_MXI2_X1 T8456 ( .Y(T8456_Y), .A(T6103_Y), .B(T16460_Q),     .S0(T5573_Q));
KC_MXI2_X1 T9667 ( .Y(T9667_Y), .A(T13770_Q), .B(T477_Y),     .S0(T12567_Y));
KC_MXI2_X1 T9516 ( .Y(T9516_Y), .A(T4799_Q), .B(T6233_Y), .S0(T173_Q));
KC_MXI2_X1 T8525 ( .Y(T8525_Y), .A(T15683_Y), .B(T2467_Y),     .S0(T8524_Y));
KC_MXI2_X1 T9836 ( .Y(T9836_Y), .A(T9743_Y), .B(T16404_Y),     .S0(T9837_Y));
KC_MXI2_X1 T9915 ( .Y(T9915_Y), .A(T1209_Q), .B(T1060_Y),     .S0(T1208_Q));
KC_MXI2_X1 T9410 ( .Y(T9410_Y), .A(T1156_Q), .B(T996_Q),     .S0(T15795_Q));
KC_MXI2_X1 T8854 ( .Y(T8854_Y), .A(T1158_Q), .B(T766_Y),     .S0(T15795_Q));
KC_MXI2_X1 T8957 ( .Y(T8957_Y), .A(T10283_Y), .B(T6417_Q),     .S0(T7919_Y));
KC_MXI2_X1 T8935 ( .Y(T8935_Y), .A(T1346_Y), .B(T1458_Y), .S0(T980_Q));
KC_MXI2_X1 T10233 ( .Y(T10233_Y), .A(T15854_Y), .B(T16299_Q),     .S0(T1176_Y));
KC_MXI2_X1 T10227 ( .Y(T10227_Y), .A(T13059_Q), .B(T5381_Y),     .S0(T1505_Y));
KC_MXI2_X1 T10209 ( .Y(T10209_Y), .A(T15858_Y), .B(T15809_Q),     .S0(T1154_Q));
KC_MXI2_X1 T9218 ( .Y(T9218_Y), .A(T12191_Y), .B(T9218_B),     .S0(T16281_Y));
KC_MXI2_X1 T8265 ( .Y(T8265_Y), .A(T5939_Y), .B(T13104_Q),     .S0(T13096_Q));
KC_MXI2_X1 T8251 ( .Y(T8251_Y), .A(T1733_Y), .B(T15815_Q),     .S0(T1775_Q));
KC_MXI2_X1 T8274 ( .Y(T8274_Y), .A(T16301_Q), .B(T2719_Y),     .S0(T5568_Q));
KC_MXI2_X1 T8343 ( .Y(T8343_Y), .A(T1786_Y), .B(T2315_Q),     .S0(T15803_Q));
KC_MXI2_X1 T8354 ( .Y(T8354_Y), .A(T16042_Y), .B(T5571_Q),     .S0(T11652_Y));
KC_MXI2_X1 T8405 ( .Y(T8405_Y), .A(T6207_Y), .B(T11762_Y),     .S0(T12856_Y));
KC_MXI2_X1 T9497 ( .Y(T9497_Y), .A(T15525_Y), .B(T9496_Y),     .S0(T5415_Y));
KC_NOR2_X2 T9255 ( .Y(T9255_Y), .A(T5220_Q), .B(T54_Q));
KC_NOR2_X2 T9254 ( .Y(T9254_Y), .A(T5220_Q), .B(T5606_Y));
KC_NOR2_X2 T9253 ( .Y(T9253_Y), .A(T15169_Y), .B(T5633_Y));
KC_NOR2_X2 T9251 ( .Y(T9251_Y), .A(T83_Q), .B(T5624_Y));
KC_NOR2_X2 T8549 ( .Y(T8549_Y), .A(T81_Q), .B(T9253_Y));
KC_NOR2_X2 T9252 ( .Y(T9252_Y), .A(T5624_Y), .B(T87_Y));
KC_NOR2_X2 T8548 ( .Y(T8548_Y), .A(T5185_Q), .B(T83_Q));
KC_NOR2_X2 T8564 ( .Y(T8564_Y), .A(T15324_Y), .B(T5634_Y));
KC_NOR2_X2 T8559 ( .Y(T8559_Y), .A(T103_Q), .B(T114_Q));
KC_NOR2_X2 T8555 ( .Y(T8555_Y), .A(T5202_Q), .B(T106_Q));
KC_NOR2_X2 T8547 ( .Y(T8547_Y), .A(T16006_Y), .B(T15320_Y));
KC_NOR2_X2 T8546 ( .Y(T8546_Y), .A(T5630_Y), .B(T12369_Y));
KC_NOR2_X2 T8545 ( .Y(T8545_Y), .A(T103_Q), .B(T15319_Y));
KC_NOR2_X2 T8543 ( .Y(T8543_Y), .A(T107_Q), .B(T5596_Y));
KC_NOR2_X2 T8537 ( .Y(T8537_Y), .A(T8536_Y), .B(T5631_Y));
KC_NOR2_X2 T33 ( .Y(T33_Y), .A(T1201_Y), .B(T16310_Y));
KC_NOR2_X2 T8558 ( .Y(T8558_Y), .A(T15316_Y), .B(T16479_Y));
KC_NOR2_X2 T8557 ( .Y(T8557_Y), .A(T8556_Y), .B(T8538_Y));
KC_NOR2_X2 T8556 ( .Y(T8556_Y), .A(T106_Q), .B(T5603_Y));
KC_NOR2_X2 T8553 ( .Y(T8553_Y), .A(T106_Q), .B(T5604_Y));
KC_NOR2_X2 T9296 ( .Y(T9296_Y), .A(T123_Y), .B(T12475_Y));
KC_NOR2_X2 T8563 ( .Y(T8563_Y), .A(T12384_Y), .B(T15841_Y));
KC_NOR2_X2 T8601 ( .Y(T8601_Y), .A(T133_Q), .B(T6321_Y));
KC_NOR2_X2 T8600 ( .Y(T8600_Y), .A(T8576_Y), .B(T12384_Y));
KC_NOR2_X2 T8599 ( .Y(T8599_Y), .A(T8598_Y), .B(T6971_Y));
KC_NOR2_X2 T8598 ( .Y(T8598_Y), .A(T236_Y), .B(T6321_Y));
KC_NOR2_X2 T8580 ( .Y(T8580_Y), .A(T136_Q), .B(T6317_Y));
KC_NOR2_X2 T8579 ( .Y(T8579_Y), .A(T5222_Q), .B(T150_Q));
KC_NOR2_X2 T8578 ( .Y(T8578_Y), .A(T6317_Y), .B(T260_Y));
KC_NOR2_X2 T8577 ( .Y(T8577_Y), .A(T15358_Y), .B(T257_Y));
KC_NOR2_X2 T8576 ( .Y(T8576_Y), .A(T8581_Y), .B(T9289_Y));
KC_NOR2_X2 T8608 ( .Y(T8608_Y), .A(T7833_Y), .B(T12383_Y));
KC_NOR2_X2 T8745 ( .Y(T8745_Y), .A(T16006_Y), .B(T646_Y));
KC_NOR2_X2 T8744 ( .Y(T8744_Y), .A(T7671_Y), .B(T12608_Y));
KC_NOR2_X2 T9026 ( .Y(T9026_Y), .A(T9079_Y), .B(T16287_Y));
KC_NOR2_X2 T9180 ( .Y(T9180_Y), .A(T15100_Y), .B(T15118_Y));
KC_NOR2_X2 T9136 ( .Y(T9136_Y), .A(T4800_Y), .B(T9181_Y));
KC_NOR2_X2 T9135 ( .Y(T9135_Y), .A(T15150_Y), .B(T15100_Y));
KC_NOR2_X2 T9087 ( .Y(T9087_Y), .A(T4818_Y), .B(T15100_Y));
KC_NOR2_X2 T9085 ( .Y(T9085_Y), .A(T4800_Y), .B(T9091_Y));
KC_NOR2_X2 T8589 ( .Y(T8589_Y), .A(T284_Q), .B(T264_Y));
KC_NOR2_X2 T8588 ( .Y(T8588_Y), .A(T278_Q), .B(T251_Y));
KC_NOR2_X2 T8575 ( .Y(T8575_Y), .A(T1487_Y), .B(T8589_Y));
KC_NOR2_X2 T8639 ( .Y(T8639_Y), .A(T5243_Q), .B(T15373_Y));
KC_NOR2_X2 T8614 ( .Y(T8614_Y), .A(T294_Q), .B(T331_Y));
KC_NOR2_X2 T8613 ( .Y(T8613_Y), .A(T6354_Y), .B(T8614_Y));
KC_NOR2_X2 T8609 ( .Y(T8609_Y), .A(T6378_Y), .B(T8639_Y));
KC_NOR2_X2 T8675 ( .Y(T8675_Y), .A(T569_Y), .B(T5281_Q));
KC_NOR2_X2 T8740 ( .Y(T8740_Y), .A(T742_Y), .B(T15429_Y));
KC_NOR2_X2 T8697 ( .Y(T8697_Y), .A(T15429_Y), .B(T9111_Y));
KC_NOR2_X2 T9425 ( .Y(T9425_Y), .A(T8950_Y), .B(T8080_Y));
KC_NOR2_X2 T9424 ( .Y(T9424_Y), .A(T9489_Y), .B(T967_Y));
KC_NOR2_X2 T9423 ( .Y(T9423_Y), .A(T1272_Y), .B(T8082_Y));
KC_NOR2_X2 T9421 ( .Y(T9421_Y), .A(T9019_Y), .B(T967_Y));
KC_NOR2_X2 T9385 ( .Y(T9385_Y), .A(T7628_Y), .B(T7816_Y));
KC_NOR2_X2 T9384 ( .Y(T9384_Y), .A(T382_Y), .B(T7825_Y));
KC_NOR2_X2 T9383 ( .Y(T9383_Y), .A(T9381_Y), .B(T7822_Y));
KC_NOR2_X2 T9375 ( .Y(T9375_Y), .A(T15429_Y), .B(T7816_Y));
KC_NOR2_X2 T8873 ( .Y(T8873_Y), .A(T7862_Y), .B(T16418_Y));
KC_NOR2_X2 T8872 ( .Y(T8872_Y), .A(T8949_Y), .B(T8080_Y));
KC_NOR2_X2 T8867 ( .Y(T8867_Y), .A(T968_Y), .B(T967_Y));
KC_NOR2_X2 T8866 ( .Y(T8866_Y), .A(T9488_Y), .B(T967_Y));
KC_NOR2_X2 T8865 ( .Y(T8865_Y), .A(T371_Y), .B(T13241_Q));
KC_NOR2_X2 T8838 ( .Y(T8838_Y), .A(T235_Q), .B(T5354_Q));
KC_NOR2_X2 T8811 ( .Y(T8811_Y), .A(T968_Y), .B(T15429_Y));
KC_NOR2_X2 T8784 ( .Y(T8784_Y), .A(T8782_Y), .B(T15452_Y));
KC_NOR2_X2 T8783 ( .Y(T8783_Y), .A(T7831_Y), .B(T8747_Y));
KC_NOR2_X2 T8782 ( .Y(T8782_Y), .A(T235_Q), .B(T921_Y));
KC_NOR2_X2 T8781 ( .Y(T8781_Y), .A(T7833_Y), .B(T8747_Y));
KC_NOR2_X2 T8780 ( .Y(T8780_Y), .A(T9384_Y), .B(T7822_Y));
KC_NOR2_X2 T8776 ( .Y(T8776_Y), .A(T382_Y), .B(T16514_Y));
KC_NOR2_X2 T8775 ( .Y(T8775_Y), .A(T16514_Y), .B(T15429_Y));
KC_NOR2_X2 T9027 ( .Y(T9027_Y), .A(T9092_Y), .B(T9078_Y));
KC_NOR2_X2 T9021 ( .Y(T9021_Y), .A(T9158_Y), .B(T9078_Y));
KC_NOR2_X2 T8965 ( .Y(T8965_Y), .A(T7858_Y), .B(T8101_Y));
KC_NOR2_X2 T8962 ( .Y(T8962_Y), .A(T16513_Y), .B(T15429_Y));
KC_NOR2_X2 T8950 ( .Y(T8950_Y), .A(T371_Y), .B(T8101_Y));
KC_NOR2_X2 T8949 ( .Y(T8949_Y), .A(T371_Y), .B(T8100_Y));
KC_NOR2_X2 T8948 ( .Y(T8948_Y), .A(T15429_Y), .B(T8101_Y));
KC_NOR2_X2 T8916 ( .Y(T8916_Y), .A(T1272_Y), .B(T8948_Y));
KC_NOR2_X2 T9171 ( .Y(T9171_Y), .A(T9174_Y), .B(T9182_Y));
KC_NOR2_X2 T9170 ( .Y(T9170_Y), .A(T9174_Y), .B(T9156_Y));
KC_NOR2_X2 T9169 ( .Y(T9169_Y), .A(T9156_Y), .B(T9014_Y));
KC_NOR2_X2 T9168 ( .Y(T9168_Y), .A(T9182_Y), .B(T9014_Y));
KC_NOR2_X2 T9165 ( .Y(T9165_Y), .A(T9127_Y), .B(T9125_Y));
KC_NOR2_X2 T9150 ( .Y(T9150_Y), .A(T9121_Y), .B(T9124_Y));
KC_NOR2_X2 T9147 ( .Y(T9147_Y), .A(T9128_Y), .B(T15524_Y));
KC_NOR2_X2 T9146 ( .Y(T9146_Y), .A(T9127_Y), .B(T15524_Y));
KC_NOR2_X2 T9122 ( .Y(T9122_Y), .A(T9127_Y), .B(T15523_Y));
KC_NOR2_X2 T9121 ( .Y(T9121_Y), .A(T15092_Y), .B(T9126_Y));
KC_NOR2_X2 T9120 ( .Y(T9120_Y), .A(T15092_Y), .B(T4801_Y));
KC_NOR2_X2 T9119 ( .Y(T9119_Y), .A(T4801_Y), .B(T2392_Y));
KC_NOR2_X2 T9118 ( .Y(T9118_Y), .A(T2392_Y), .B(T15091_Y));
KC_NOR2_X2 T9117 ( .Y(T9117_Y), .A(T15093_Y), .B(T15109_Y));
KC_NOR2_X2 T9108 ( .Y(T9108_Y), .A(T9128_Y), .B(T9125_Y));
KC_NOR2_X2 T9106 ( .Y(T9106_Y), .A(T9128_Y), .B(T15523_Y));
KC_NOR2_X2 T9105 ( .Y(T9105_Y), .A(T9129_Y), .B(T15523_Y));
KC_NOR2_X2 T9103 ( .Y(T9103_Y), .A(T9129_Y), .B(T9125_Y));
KC_NOR2_X2 T9086 ( .Y(T9086_Y), .A(T11302_Y), .B(T9073_Y));
KC_NOR2_X2 T9070 ( .Y(T9070_Y), .A(T9077_Y), .B(T9125_Y));
KC_NOR2_X2 T9069 ( .Y(T9069_Y), .A(T2390_Y), .B(T15109_Y));
KC_NOR2_X2 T9063 ( .Y(T9063_Y), .A(T9077_Y), .B(T15523_Y));
KC_NOR2_X2 T9199 ( .Y(T9199_Y), .A(T4917_Y), .B(T5228_Y));
KC_NOR2_X2 T9295 ( .Y(T9295_Y), .A(T6347_Y), .B(T9294_Y));
KC_NOR2_X2 T9294 ( .Y(T9294_Y), .A(T272_Q), .B(T217_Y));
KC_NOR2_X2 T9284 ( .Y(T9284_Y), .A(T273_Q), .B(T285_Y));
KC_NOR2_X2 T8594 ( .Y(T8594_Y), .A(T283_Q), .B(T15357_Y));
KC_NOR2_X2 T8587 ( .Y(T8587_Y), .A(T511_Y), .B(T8594_Y));
KC_NOR2_X2 T9265 ( .Y(T9265_Y), .A(T1498_Y), .B(T9284_Y));
KC_NOR2_X2 T9257 ( .Y(T9257_Y), .A(T6376_Y), .B(T8623_Y));
KC_NOR2_X2 T8623 ( .Y(T8623_Y), .A(T274_Q), .B(T342_Y));
KC_NOR2_X2 T8652 ( .Y(T8652_Y), .A(T7268_Y), .B(T7255_Y));
KC_NOR2_X2 T8644 ( .Y(T8644_Y), .A(T9512_Y), .B(T7289_Y));
KC_NOR2_X2 T9345 ( .Y(T9345_Y), .A(T7604_Y), .B(T7452_Y));
KC_NOR2_X2 T8680 ( .Y(T8680_Y), .A(T7625_Y), .B(T7386_Y));
KC_NOR2_X2 T8673 ( .Y(T8673_Y), .A(T6397_Y), .B(T535_Y));
KC_NOR2_X2 T8672 ( .Y(T8672_Y), .A(T7624_Y), .B(T7429_Y));
KC_NOR2_X2 T8668 ( .Y(T8668_Y), .A(T7396_Y), .B(T9326_Y));
KC_NOR2_X2 T8662 ( .Y(T8662_Y), .A(T499_Y), .B(T699_Q));
KC_NOR2_X2 T8753 ( .Y(T8753_Y), .A(T8086_Y), .B(T794_Y));
KC_NOR2_X2 T8752 ( .Y(T8752_Y), .A(T9016_Y), .B(T794_Y));
KC_NOR2_X2 T8742 ( .Y(T8742_Y), .A(T742_Y), .B(T794_Y));
KC_NOR2_X2 T8741 ( .Y(T8741_Y), .A(T382_Y), .B(T9111_Y));
KC_NOR2_X2 T8698 ( .Y(T8698_Y), .A(T9178_Y), .B(T794_Y));
KC_NOR2_X2 T8868 ( .Y(T8868_Y), .A(T371_Y), .B(T9110_Y));
KC_NOR2_X2 T8864 ( .Y(T8864_Y), .A(T15841_Y), .B(T8067_Y));
KC_NOR2_X2 T8863 ( .Y(T8863_Y), .A(T8946_Y), .B(T69_Y));
KC_NOR2_X2 T8810 ( .Y(T8810_Y), .A(T7697_Y), .B(T7844_Y));
KC_NOR2_X2 T8777 ( .Y(T8777_Y), .A(T382_Y), .B(T13241_Q));
KC_NOR2_X2 T9013 ( .Y(T9013_Y), .A(T9028_Y), .B(T745_Y));
KC_NOR2_X2 T8981 ( .Y(T8981_Y), .A(T5378_Q), .B(T5377_Q));
KC_NOR2_X2 T8980 ( .Y(T8980_Y), .A(T750_Q), .B(T8116_Y));
KC_NOR2_X2 T8979 ( .Y(T8979_Y), .A(T8119_Y), .B(T1200_Y));
KC_NOR2_X2 T8963 ( .Y(T8963_Y), .A(T371_Y), .B(T16513_Y));
KC_NOR2_X2 T9107 ( .Y(T9107_Y), .A(T1841_Y), .B(T9113_Y));
KC_NOR2_X2 T9062 ( .Y(T9062_Y), .A(T1594_Y), .B(T9060_Y));
KC_NOR2_X2 T9061 ( .Y(T9061_Y), .A(T605_Q), .B(T1593_Y));
KC_NOR2_X2 T9060 ( .Y(T9060_Y), .A(T1593_Y), .B(T598_Y));
KC_NOR2_X2 T9243 ( .Y(T9243_Y), .A(T4842_Y), .B(T15538_Y));
KC_NOR2_X2 T9194 ( .Y(T9194_Y), .A(T4842_Y), .B(T15540_Y));
KC_NOR2_X2 T9292 ( .Y(T9292_Y), .A(T5196_Q), .B(T15352_Y));
KC_NOR2_X2 T8562 ( .Y(T8562_Y), .A(T12881_Y), .B(T12375_Y));
KC_NOR2_X2 T8593 ( .Y(T8593_Y), .A(T443_Q), .B(T237_Y));
KC_NOR2_X2 T8592 ( .Y(T8592_Y), .A(T12474_Y), .B(T12388_Y));
KC_NOR2_X2 T8584 ( .Y(T8584_Y), .A(T12478_Y), .B(T12386_Y));
KC_NOR2_X2 T8570 ( .Y(T8570_Y), .A(T626_Q), .B(T246_Y));
KC_NOR2_X2 T8565 ( .Y(T8565_Y), .A(T628_Q), .B(T15351_Y));
KC_NOR2_X2 T9264 ( .Y(T9264_Y), .A(T276_Q), .B(T6304_Y));
KC_NOR2_X2 T8617 ( .Y(T8617_Y), .A(T435_Q), .B(T6331_Y));
KC_NOR2_X2 T8616 ( .Y(T8616_Y), .A(T12495_Y), .B(T6330_Y));
KC_NOR2_X2 T8612 ( .Y(T8612_Y), .A(T5198_Q), .B(T324_Y));
KC_NOR2_X2 T8604 ( .Y(T8604_Y), .A(T12880_Y), .B(T6258_Y));
KC_NOR2_X2 T8650 ( .Y(T8650_Y), .A(T673_Y), .B(T13232_Y));
KC_NOR2_X2 T9334 ( .Y(T9334_Y), .A(T7685_Y), .B(T7645_Y));
KC_NOR2_X2 T8735 ( .Y(T8735_Y), .A(T7646_Y), .B(T900_Y));
KC_NOR2_X2 T8734 ( .Y(T8734_Y), .A(T8832_Y), .B(T7563_Y));
KC_NOR2_X2 T8733 ( .Y(T8733_Y), .A(T8832_Y), .B(T7644_Y));
KC_NOR2_X2 T9416 ( .Y(T9416_Y), .A(T8120_Y), .B(T941_Y));
KC_NOR2_X2 T8860 ( .Y(T8860_Y), .A(T7892_Y), .B(T720_Y));
KC_NOR2_X2 T8859 ( .Y(T8859_Y), .A(T15842_Y), .B(T720_Y));
KC_NOR2_X2 T8855 ( .Y(T8855_Y), .A(T15842_Y), .B(T9446_Y));
KC_NOR2_X2 T8805 ( .Y(T8805_Y), .A(T8859_Y), .B(T8860_Y));
KC_NOR2_X2 T8769 ( .Y(T8769_Y), .A(T7645_Y), .B(T900_Y));
KC_NOR2_X2 T8767 ( .Y(T8767_Y), .A(T900_Y), .B(T7801_Y));
KC_NOR2_X2 T8766 ( .Y(T8766_Y), .A(T7563_Y), .B(T900_Y));
KC_NOR2_X2 T9011 ( .Y(T9011_Y), .A(T16006_Y), .B(T16278_Y));
KC_NOR2_X2 T8978 ( .Y(T8978_Y), .A(T16311_Y), .B(T1323_Y));
KC_NOR2_X2 T8977 ( .Y(T8977_Y), .A(T556_Q), .B(T8130_Y));
KC_NOR2_X2 T8975 ( .Y(T8975_Y), .A(T13241_Q), .B(T9014_Y));
KC_NOR2_X2 T8944 ( .Y(T8944_Y), .A(T12456_Y), .B(T1255_Y));
KC_NOR2_X2 T8943 ( .Y(T8943_Y), .A(T8941_Y), .B(T8034_Y));
KC_NOR2_X2 T8902 ( .Y(T8902_Y), .A(T12456_Y), .B(T12368_Y));
KC_NOR2_X2 T8901 ( .Y(T8901_Y), .A(T8902_Y), .B(T11267_Y));
KC_NOR2_X2 T9439 ( .Y(T9439_Y), .A(T10941_Y), .B(T9437_Y));
KC_NOR2_X2 T8569 ( .Y(T8569_Y), .A(T12476_Y), .B(T12380_Y));
KC_NOR2_X2 T8630 ( .Y(T8630_Y), .A(T11085_Y), .B(T16510_Y));
KC_NOR2_X2 T8611 ( .Y(T8611_Y), .A(T12497_Y), .B(T12391_Y));
KC_NOR2_X2 T9501 ( .Y(T9501_Y), .A(T7592_Y), .B(T6630_Y));
KC_NOR2_X2 T9500 ( .Y(T9500_Y), .A(T7592_Y), .B(T6700_Y));
KC_NOR2_X2 T8640 ( .Y(T8640_Y), .A(T829_Q), .B(T380_Y));
KC_NOR2_X2 T6826 ( .Y(T6826_Y), .A(T15408_Y), .B(T9360_Y));
KC_NOR2_X2 T9313 ( .Y(T9313_Y), .A(T7685_Y), .B(T7644_Y));
KC_NOR2_X2 T9303 ( .Y(T9303_Y), .A(T15408_Y), .B(T8758_Y));
KC_NOR2_X2 T9301 ( .Y(T9301_Y), .A(T15408_Y), .B(T8762_Y));
KC_NOR2_X2 T8670 ( .Y(T8670_Y), .A(T7839_Y), .B(T553_Y));
KC_NOR2_X2 T8656 ( .Y(T8656_Y), .A(T15408_Y), .B(T1039_Y));
KC_NOR2_X2 T8748 ( .Y(T8748_Y), .A(T7839_Y), .B(T10942_Y));
KC_NOR2_X2 T8727 ( .Y(T8727_Y), .A(T15454_Y), .B(T7614_Y));
KC_NOR2_X2 T8725 ( .Y(T8725_Y), .A(T886_Y), .B(T652_Y));
KC_NOR2_X2 T8718 ( .Y(T8718_Y), .A(T7592_Y), .B(T730_Y));
KC_NOR2_X2 T8716 ( .Y(T8716_Y), .A(T7592_Y), .B(T7614_Y));
KC_NOR2_X2 T8715 ( .Y(T8715_Y), .A(T9359_Y), .B(T15408_Y));
KC_NOR2_X2 T8707 ( .Y(T8707_Y), .A(T15408_Y), .B(T9362_Y));
KC_NOR2_X2 T8682 ( .Y(T8682_Y), .A(T744_Y), .B(T7557_Y));
KC_NOR2_X2 T9367 ( .Y(T9367_Y), .A(T16159_Y), .B(T4872_Y));
KC_NOR2_X2 T9366 ( .Y(T9366_Y), .A(T9367_Y), .B(T764_Y));
KC_NOR2_X2 T8847 ( .Y(T8847_Y), .A(T950_Y), .B(T8936_Y));
KC_NOR2_X2 T8846 ( .Y(T8846_Y), .A(T992_Q), .B(T981_Q));
KC_NOR2_X2 T8845 ( .Y(T8845_Y), .A(T992_Q), .B(T15457_Y));
KC_NOR2_X2 T8831 ( .Y(T8831_Y), .A(T16275_Y), .B(T10880_Y));
KC_NOR2_X2 T8829 ( .Y(T8829_Y), .A(T16275_Y), .B(T16274_Y));
KC_NOR2_X2 T8828 ( .Y(T8828_Y), .A(T16159_Y), .B(T15999_Y));
KC_NOR2_X2 T8827 ( .Y(T8827_Y), .A(T16159_Y), .B(T10941_Y));
KC_NOR2_X2 T8804 ( .Y(T8804_Y), .A(T16509_Y), .B(T8801_Y));
KC_NOR2_X2 T8797 ( .Y(T8797_Y), .A(T9406_Y), .B(T8799_Y));
KC_NOR2_X2 T8796 ( .Y(T8796_Y), .A(T15458_Y), .B(T949_Q));
KC_NOR2_X2 T8795 ( .Y(T8795_Y), .A(T939_Q), .B(T949_Q));
KC_NOR2_X2 T8794 ( .Y(T8794_Y), .A(T1133_Q), .B(T8798_Y));
KC_NOR2_X2 T8792 ( .Y(T8792_Y), .A(T8797_Y), .B(T16006_Y));
KC_NOR2_X2 T8791 ( .Y(T8791_Y), .A(T947_Y), .B(T7881_Y));
KC_NOR2_X2 T8790 ( .Y(T8790_Y), .A(T7841_Y), .B(T7881_Y));
KC_NOR2_X2 T8771 ( .Y(T8771_Y), .A(T758_Y), .B(T7848_Y));
KC_NOR2_X2 T8770 ( .Y(T8770_Y), .A(T8946_Y), .B(T908_Y));
KC_NOR2_X2 T8768 ( .Y(T8768_Y), .A(T1247_Q), .B(T1249_Q));
KC_NOR2_X2 T8765 ( .Y(T8765_Y), .A(T1249_Q), .B(T903_Y));
KC_NOR2_X2 T8763 ( .Y(T8763_Y), .A(T758_Y), .B(T12449_Y));
KC_NOR2_X2 T8762 ( .Y(T8762_Y), .A(T10941_Y), .B(T7802_Y));
KC_NOR2_X2 T8761 ( .Y(T8761_Y), .A(T8760_Y), .B(T8759_Y));
KC_NOR2_X2 T8760 ( .Y(T8760_Y), .A(T786_Y), .B(T764_Y));
KC_NOR2_X2 T8759 ( .Y(T8759_Y), .A(T8827_Y), .B(T764_Y));
KC_NOR2_X2 T8758 ( .Y(T8758_Y), .A(T4872_Y), .B(T7802_Y));
KC_NOR2_X2 T8757 ( .Y(T8757_Y), .A(T4872_Y), .B(T783_Y));
KC_NOR2_X2 T8756 ( .Y(T8756_Y), .A(T8938_Y), .B(T10941_Y));
KC_NOR2_X2 T8997 ( .Y(T8997_Y), .A(T4847_Y), .B(T9438_Y));
KC_NOR2_X2 T8936 ( .Y(T8936_Y), .A(T941_Y), .B(T9402_Y));
KC_NOR2_X2 T8889 ( .Y(T8889_Y), .A(T8031_Y), .B(T12884_Y));
KC_NOR2_X2 T9440 ( .Y(T9440_Y), .A(T4872_Y), .B(T9437_Y));
KC_NOR2_X2 T9032 ( .Y(T9032_Y), .A(T4847_Y), .B(T10301_Y));
KC_NOR2_X2 T6825 ( .Y(T6825_Y), .A(T7839_Y), .B(T6822_Y));
KC_NOR2_X2 T9723 ( .Y(T9723_Y), .A(T15775_Y), .B(T7549_Y));
KC_NOR2_X2 T9302 ( .Y(T9302_Y), .A(T8717_Y), .B(T7592_Y));
KC_NOR2_X2 T9819 ( .Y(T9819_Y), .A(T15841_Y), .B(T9817_Y));
KC_NOR2_X2 T9818 ( .Y(T9818_Y), .A(T15841_Y), .B(T9813_Y));
KC_NOR2_X2 T9815 ( .Y(T9815_Y), .A(T15841_Y), .B(T9814_Y));
KC_NOR2_X2 T8726 ( .Y(T8726_Y), .A(T5561_Q), .B(T5297_Q));
KC_NOR2_X2 T8717 ( .Y(T8717_Y), .A(T16091_Y), .B(T7612_Y));
KC_NOR2_X2 T8686 ( .Y(T8686_Y), .A(T15841_Y), .B(T9783_Y));
KC_NOR2_X2 T8685 ( .Y(T8685_Y), .A(T15841_Y), .B(T9357_Y));
KC_NOR2_X2 T8684 ( .Y(T8684_Y), .A(T5359_Q), .B(T5360_Q));
KC_NOR2_X2 T8683 ( .Y(T8683_Y), .A(T15792_Y), .B(T7554_Y));
KC_NOR2_X2 T10651 ( .Y(T10651_Y), .A(T16422_Q), .B(T1007_Y));
KC_NOR2_X2 T9919 ( .Y(T9919_Y), .A(T1095_Q), .B(T1100_Q));
KC_NOR2_X2 T9900 ( .Y(T9900_Y), .A(T8849_Y), .B(T7976_Y));
KC_NOR2_X2 T9899 ( .Y(T9899_Y), .A(T9402_Y), .B(T540_Y));
KC_NOR2_X2 T9898 ( .Y(T9898_Y), .A(T9402_Y), .B(T1042_Y));
KC_NOR2_X2 T9897 ( .Y(T9897_Y), .A(T9402_Y), .B(T378_Y));
KC_NOR2_X2 T9896 ( .Y(T9896_Y), .A(T1062_Y), .B(T9402_Y));
KC_NOR2_X2 T9891 ( .Y(T9891_Y), .A(T1481_Y), .B(T1131_Q));
KC_NOR2_X2 T9890 ( .Y(T9890_Y), .A(T15841_Y), .B(T11245_Y));
KC_NOR2_X2 T9368 ( .Y(T9368_Y), .A(T15841_Y), .B(T9358_Y));
KC_NOR2_X2 T8830 ( .Y(T8830_Y), .A(T15841_Y), .B(T9928_Y));
KC_NOR2_X2 T10049 ( .Y(T10049_Y), .A(T1133_Q), .B(T1130_Q));
KC_NOR2_X2 T10023 ( .Y(T10023_Y), .A(T5376_Q), .B(T10045_Y));
KC_NOR2_X2 T9988 ( .Y(T9988_Y), .A(T10008_Y), .B(T1341_Y));
KC_NOR2_X2 T8974 ( .Y(T8974_Y), .A(T140_Y), .B(T10004_Y));
KC_NOR2_X2 T8891 ( .Y(T8891_Y), .A(T951_Y), .B(T7879_Y));
KC_NOR2_X2 T8890 ( .Y(T8890_Y), .A(T7879_Y), .B(T11894_Y));
KC_NOR2_X2 T10162 ( .Y(T10162_Y), .A(T16420_Y), .B(T12724_Y));
KC_NOR2_X2 T10160 ( .Y(T10160_Y), .A(T1133_Q), .B(T10007_Y));
KC_NOR2_X2 T9031 ( .Y(T9031_Y), .A(T4847_Y), .B(T10303_Y));
KC_NOR2_X2 T9926 ( .Y(T9926_Y), .A(T9898_Y), .B(T1085_Y));
KC_NOR2_X2 T9917 ( .Y(T9917_Y), .A(T5334_Q), .B(T1210_Q));
KC_NOR2_X2 T10040 ( .Y(T10040_Y), .A(T1249_Q), .B(T10046_Y));
KC_NOR2_X2 T10024 ( .Y(T10024_Y), .A(T1249_Q), .B(T1125_Y));
KC_NOR2_X2 T10006 ( .Y(T10006_Y), .A(T1222_Q), .B(T5375_Q));
KC_NOR2_X2 T10005 ( .Y(T10005_Y), .A(T7949_Y), .B(T1248_Y));
KC_NOR2_X2 T10004 ( .Y(T10004_Y), .A(T10159_Y), .B(T10302_Y));
KC_NOR2_X2 T10003 ( .Y(T10003_Y), .A(T7949_Y), .B(T10002_Y));
KC_NOR2_X2 T10002 ( .Y(T10002_Y), .A(T7951_Y), .B(T10315_Y));
KC_NOR2_X2 T9998 ( .Y(T9998_Y), .A(T11914_Y), .B(T10302_Y));
KC_NOR2_X2 T9981 ( .Y(T9981_Y), .A(T7949_Y), .B(T10737_Y));
KC_NOR2_X2 T10284 ( .Y(T10284_Y), .A(T13053_Q), .B(T4865_Y));
KC_NOR2_X2 T10163 ( .Y(T10163_Y), .A(T12446_Y), .B(T16005_Y));
KC_NOR2_X2 T10161 ( .Y(T10161_Y), .A(T4868_Y), .B(T10158_Y));
KC_NOR2_X2 T10156 ( .Y(T10156_Y), .A(T16275_Y), .B(T4868_Y));
KC_NOR2_X2 T10155 ( .Y(T10155_Y), .A(T1365_Y), .B(T4902_Y));
KC_NOR2_X2 T10154 ( .Y(T10154_Y), .A(T4847_Y), .B(T4838_Y));
KC_NOR2_X2 T10139 ( .Y(T10139_Y), .A(T1362_Y), .B(T1366_Y));
KC_NOR2_X2 T10130 ( .Y(T10130_Y), .A(T2717_Y), .B(T4831_Y));
KC_NOR2_X2 T16171 ( .Y(T16171_Y), .A(T1505_Y), .B(T13059_Q));
KC_NOR2_X2 T9586 ( .Y(T9586_Y), .A(T7182_Y), .B(T9581_Y));
KC_NOR2_X2 T9585 ( .Y(T9585_Y), .A(T356_Y), .B(T9581_Y));
KC_NOR2_X2 T9579 ( .Y(T9579_Y), .A(T356_Y), .B(T9582_Y));
KC_NOR2_X2 T9578 ( .Y(T9578_Y), .A(T15378_Y), .B(T9633_Y));
KC_NOR2_X2 T9577 ( .Y(T9577_Y), .A(T15378_Y), .B(T9631_Y));
KC_NOR2_X2 T9576 ( .Y(T9576_Y), .A(T15378_Y), .B(T9632_Y));
KC_NOR2_X2 T9575 ( .Y(T9575_Y), .A(T356_Y), .B(T10403_Y));
KC_NOR2_X2 T9574 ( .Y(T9574_Y), .A(T7182_Y), .B(T10403_Y));
KC_NOR2_X2 T9573 ( .Y(T9573_Y), .A(T7182_Y), .B(T9582_Y));
KC_NOR2_X2 T10423 ( .Y(T10423_Y), .A(T5674_Y), .B(T10426_Y));
KC_NOR2_X2 T10422 ( .Y(T10422_Y), .A(T7339_Y), .B(T10372_Y));
KC_NOR2_X2 T10421 ( .Y(T10421_Y), .A(T6748_Y), .B(T10424_Y));
KC_NOR2_X2 T10420 ( .Y(T10420_Y), .A(T5674_Y), .B(T10427_Y));
KC_NOR2_X2 T10419 ( .Y(T10419_Y), .A(T15677_Y), .B(T10427_Y));
KC_NOR2_X2 T10418 ( .Y(T10418_Y), .A(T15677_Y), .B(T10428_Y));
KC_NOR2_X2 T10206 ( .Y(T10206_Y), .A(T1361_Q), .B(T16081_Q));
KC_NOR2_X2 T10388 ( .Y(T10388_Y), .A(T3728_Y), .B(T3070_Y));
KC_NOR2_X2 T9539 ( .Y(T9539_Y), .A(T3728_Y), .B(T3070_Y));
KC_NOR2_X2 T9719 ( .Y(T9719_Y), .A(T3728_Y), .B(T3070_Y));
KC_NOR2_X2 T10013 ( .Y(T10013_Y), .A(T3728_Y), .B(T3070_Y));
KC_NOR2_X2 T10362 ( .Y(T10362_Y), .A(T6791_Y), .B(T10356_Y));
KC_NOR2_X2 T10347 ( .Y(T10347_Y), .A(T5650_Y), .B(T10410_Y));
KC_NOR2_X2 T10346 ( .Y(T10346_Y), .A(T6789_Y), .B(T10410_Y));
KC_NOR2_X2 T9712 ( .Y(T9712_Y), .A(T5663_Y), .B(T10356_Y));
KC_NOR2_X2 T9706 ( .Y(T9706_Y), .A(T6789_Y), .B(T10411_Y));
KC_NOR2_X2 T9704 ( .Y(T9704_Y), .A(T5650_Y), .B(T10411_Y));
KC_NOR2_X2 T9809 ( .Y(T9809_Y), .A(T3728_Y), .B(T3070_Y));
KC_NOR2_X2 T9781 ( .Y(T9781_Y), .A(T4919_Y), .B(T4920_Y));
KC_NOR2_X2 T8862 ( .Y(T8862_Y), .A(T8002_Y), .B(T9924_Y));
KC_NOR2_X2 T10306 ( .Y(T10306_Y), .A(T1479_Y), .B(T9894_Y));
KC_NOR2_X2 T9902 ( .Y(T9902_Y), .A(T8004_Y), .B(T9921_Y));
KC_NOR2_X2 T9893 ( .Y(T9893_Y), .A(T1054_Y), .B(T9921_Y));
KC_NOR2_X2 T9892 ( .Y(T9892_Y), .A(T1054_Y), .B(T10319_Y));
KC_NOR2_X2 T9883 ( .Y(T9883_Y), .A(T8002_Y), .B(T9894_Y));
KC_NOR2_X2 T10033 ( .Y(T10033_Y), .A(T1479_Y), .B(T9922_Y));
KC_NOR2_X2 T10009 ( .Y(T10009_Y), .A(T8002_Y), .B(T9922_Y));
KC_NOR2_X2 T10397 ( .Y(T10397_Y), .A(T6462_Y), .B(T9612_Y));
KC_NOR2_X2 T9580 ( .Y(T9580_Y), .A(T6462_Y), .B(T9611_Y));
KC_NOR2_X2 T10408 ( .Y(T10408_Y), .A(T6768_Y), .B(T6751_Y));
KC_NOR2_X2 T10407 ( .Y(T10407_Y), .A(T6768_Y), .B(T15693_Y));
KC_NOR2_X2 T10406 ( .Y(T10406_Y), .A(T6768_Y), .B(T6752_Y));
KC_NOR2_X2 T9686 ( .Y(T9686_Y), .A(T6768_Y), .B(T458_Y));
KC_NOR2_X2 T9657 ( .Y(T9657_Y), .A(T6768_Y), .B(T461_Y));
KC_NOR2_X2 T9604 ( .Y(T9604_Y), .A(T6768_Y), .B(T494_Y));
KC_NOR2_X2 T8535 ( .Y(T8535_Y), .A(T6768_Y), .B(T6753_Y));
KC_NOR2_X2 T8534 ( .Y(T8534_Y), .A(T6768_Y), .B(T15675_Y));
KC_NOR2_X2 T10094 ( .Y(T10094_Y), .A(T10070_Y), .B(T15073_Y));
KC_NOR2_X2 T10223 ( .Y(T10223_Y), .A(T15904_Y), .B(T1805_Y));
KC_NOR2_X2 T10210 ( .Y(T10210_Y), .A(T15904_Y), .B(T4968_Y));
KC_NOR2_X2 T5910 ( .Y(T5910_Y), .A(T12815_Y), .B(T15974_Y));
KC_NOR2_X2 T5904 ( .Y(T5904_Y), .A(T5899_Y), .B(T1770_Y));
KC_NOR2_X2 T5899 ( .Y(T5899_Y), .A(T1768_Y), .B(T2175_Y));
KC_NOR2_X2 T11532 ( .Y(T11532_Y), .A(T1762_Y), .B(T1772_Y));
KC_NOR2_X2 T11531 ( .Y(T11531_Y), .A(T1762_Y), .B(T2175_Y));
KC_NOR2_X2 T11502 ( .Y(T11502_Y), .A(T1768_Y), .B(T5460_Y));
KC_NOR2_X2 T11494 ( .Y(T11494_Y), .A(T1768_Y), .B(T1772_Y));
KC_NOR2_X2 T11493 ( .Y(T11493_Y), .A(T11532_Y), .B(T11494_Y));
KC_NOR2_X2 T11482 ( .Y(T11482_Y), .A(T1767_Y), .B(T1773_Y));
KC_NOR2_X2 T11047 ( .Y(T11047_Y), .A(T6519_Y), .B(T11828_Y));
KC_NOR2_X2 T11757 ( .Y(T11757_Y), .A(T6519_Y), .B(T11756_Y));
KC_NOR2_X2 T11756 ( .Y(T11756_Y), .A(T11766_Y), .B(T2338_Y));
KC_NOR2_X2 T11755 ( .Y(T11755_Y), .A(T6199_Y), .B(T2326_Y));
KC_NOR2_X2 T11754 ( .Y(T11754_Y), .A(T6201_Y), .B(T2326_Y));
KC_NOR2_X2 T11753 ( .Y(T11753_Y), .A(T2338_Y), .B(T2326_Y));
KC_NOR2_X2 T11752 ( .Y(T11752_Y), .A(T6520_Y), .B(T11756_Y));
KC_NOR2_X2 T11751 ( .Y(T11751_Y), .A(T6522_Y), .B(T11756_Y));
KC_NOR2_X2 T11046 ( .Y(T11046_Y), .A(T6518_Y), .B(T11756_Y));
KC_NOR2_X2 T11045 ( .Y(T11045_Y), .A(T6522_Y), .B(T11828_Y));
KC_NOR2_X2 T11044 ( .Y(T11044_Y), .A(T6518_Y), .B(T11828_Y));
KC_NOR2_X2 T11845 ( .Y(T11845_Y), .A(T8434_Y), .B(T6494_Y));
KC_NOR2_X2 T11828 ( .Y(T11828_Y), .A(T11766_Y), .B(T2960_Y));
KC_NOR2_X2 T9681 ( .Y(T9681_Y), .A(T15682_Y), .B(T409_Y));
KC_NOR2_X2 T9680 ( .Y(T9680_Y), .A(T15682_Y), .B(T490_Y));
KC_NOR2_X2 T9679 ( .Y(T9679_Y), .A(T6768_Y), .B(T485_Y));
KC_NOR2_X2 T9678 ( .Y(T9678_Y), .A(T15682_Y), .B(T491_Y));
KC_NOR2_X2 T9677 ( .Y(T9677_Y), .A(T15682_Y), .B(T15399_Y));
KC_NOR2_X2 T9646 ( .Y(T9646_Y), .A(T6768_Y), .B(T451_Y));
KC_NOR2_X2 T9642 ( .Y(T9642_Y), .A(T2449_Y), .B(T2448_Y));
KC_NOR2_X2 T8532 ( .Y(T8532_Y), .A(T6768_Y), .B(T15692_Y));
KC_NOR2_X2 T8531 ( .Y(T8531_Y), .A(T6768_Y), .B(T6777_Y));
KC_NOR2_X2 T8530 ( .Y(T8530_Y), .A(T6768_Y), .B(T6756_Y));
KC_NOR2_X2 T8527 ( .Y(T8527_Y), .A(T6768_Y), .B(T6757_Y));
KC_NOR2_X2 T9880 ( .Y(T9880_Y), .A(T15474_Y), .B(T4973_Y));
KC_NOR2_X2 T9843 ( .Y(T9843_Y), .A(T16406_Y), .B(T2025_Y));
KC_NOR2_X2 T10524 ( .Y(T10524_Y), .A(T10526_Y), .B(T10519_Y));
KC_NOR2_X2 T10523 ( .Y(T10523_Y), .A(T2023_Q), .B(T2008_Q));
KC_NOR2_X2 T10516 ( .Y(T10516_Y), .A(T2016_Q), .B(T16366_Y));
KC_NOR2_X2 T9970 ( .Y(T9970_Y), .A(T10100_Y), .B(T1496_Y));
KC_NOR2_X2 T9969 ( .Y(T9969_Y), .A(T2005_Q), .B(T9973_Y));
KC_NOR2_X2 T9968 ( .Y(T9968_Y), .A(T2018_Y), .B(T2040_Y));
KC_NOR2_X2 T9950 ( .Y(T9950_Y), .A(T2016_Q), .B(T1985_Y));
KC_NOR2_X2 T9949 ( .Y(T9949_Y), .A(T1116_Y), .B(T1990_Y));
KC_NOR2_X2 T10093 ( .Y(T10093_Y), .A(T10106_Y), .B(T15089_Y));
KC_NOR2_X2 T10078 ( .Y(T10078_Y), .A(T2550_Y), .B(T16411_Y));
KC_NOR2_X2 T10064 ( .Y(T10064_Y), .A(T2034_Y), .B(T5369_Y));
KC_NOR2_X2 T10184 ( .Y(T10184_Y), .A(T13131_Y), .B(T16266_Y));
KC_NOR2_X2 T11432 ( .Y(T11432_Y), .A(T15916_Y), .B(T4942_Y));
KC_NOR2_X2 T11474 ( .Y(T11474_Y), .A(T5058_Y), .B(T2165_Y));
KC_NOR2_X2 T11473 ( .Y(T11473_Y), .A(T5058_Y), .B(T2722_Y));
KC_NOR2_X2 T11450 ( .Y(T11450_Y), .A(T5455_Q), .B(T2151_Q));
KC_NOR2_X2 T11437 ( .Y(T11437_Y), .A(T5058_Y), .B(T2145_Y));
KC_NOR2_X2 T11436 ( .Y(T11436_Y), .A(T15882_Y), .B(T15943_Y));
KC_NOR2_X2 T11530 ( .Y(T11530_Y), .A(T5460_Y), .B(T1762_Y));
KC_NOR2_X2 T11517 ( .Y(T11517_Y), .A(T2800_Y), .B(T8238_Y));
KC_NOR2_X2 T11501 ( .Y(T11501_Y), .A(T5983_Y), .B(T8238_Y));
KC_NOR2_X2 T11500 ( .Y(T11500_Y), .A(T11025_Y), .B(T2168_Y));
KC_NOR2_X2 T11492 ( .Y(T11492_Y), .A(T15590_Y), .B(T8238_Y));
KC_NOR2_X2 T11586 ( .Y(T11586_Y), .A(T2800_Y), .B(T6511_Y));
KC_NOR2_X2 T11551 ( .Y(T11551_Y), .A(T5058_Y), .B(T6511_Y));
KC_NOR2_X2 T11622 ( .Y(T11622_Y), .A(T2854_Y), .B(T12219_Y));
KC_NOR2_X2 T11613 ( .Y(T11613_Y), .A(T2854_Y), .B(T2217_Y));
KC_NOR2_X2 T10626 ( .Y(T10626_Y), .A(T2345_Q), .B(T2261_Y));
KC_NOR2_X2 T10612 ( .Y(T10612_Y), .A(T2315_Q), .B(T2293_Y));
KC_NOR2_X2 T10597 ( .Y(T10597_Y), .A(T2316_Q), .B(T2298_Y));
KC_NOR2_X2 T10573 ( .Y(T10573_Y), .A(T16270_Y), .B(T12103_Y));
KC_NOR2_X2 T11776 ( .Y(T11776_Y), .A(T6559_Y), .B(T3483_Y));
KC_NOR2_X2 T11775 ( .Y(T11775_Y), .A(T2344_Y), .B(T3483_Y));
KC_NOR2_X2 T11774 ( .Y(T11774_Y), .A(T12105_Y), .B(T6229_Y));
KC_NOR2_X2 T11773 ( .Y(T11773_Y), .A(T4926_Y), .B(T3483_Y));
KC_NOR2_X2 T11750 ( .Y(T11750_Y), .A(T2838_Y), .B(T8172_Y));
KC_NOR2_X2 T10562 ( .Y(T10562_Y), .A(T15713_Y), .B(T2343_Y));
KC_NOR2_X2 T10558 ( .Y(T10558_Y), .A(T15712_Y), .B(T6101_Y));
KC_NOR2_X2 T11826 ( .Y(T11826_Y), .A(T6543_Y), .B(T291_Y));
KC_NOR2_X2 T8155 ( .Y(T8155_Y), .A(T12879_Y), .B(T6605_Y));
KC_NOR2_X2 T10438 ( .Y(T10438_Y), .A(T15682_Y), .B(T6457_Y));
KC_NOR2_X2 T9671 ( .Y(T9671_Y), .A(T15682_Y), .B(T444_Y));
KC_NOR2_X2 T9670 ( .Y(T9670_Y), .A(T15682_Y), .B(T477_Y));
KC_NOR2_X2 T9656 ( .Y(T9656_Y), .A(T15682_Y), .B(T437_Y));
KC_NOR2_X2 T9653 ( .Y(T9653_Y), .A(T15682_Y), .B(T418_Y));
KC_NOR2_X2 T9645 ( .Y(T9645_Y), .A(T15682_Y), .B(T6758_Y));
KC_NOR2_X2 T9641 ( .Y(T9641_Y), .A(T15682_Y), .B(T6458_Y));
KC_NOR2_X2 T9640 ( .Y(T9640_Y), .A(T15682_Y), .B(T406_Y));
KC_NOR2_X2 T9639 ( .Y(T9639_Y), .A(T15682_Y), .B(T404_Y));
KC_NOR2_X2 T10493 ( .Y(T10493_Y), .A(T10941_Y), .B(T2068_Y));
KC_NOR2_X2 T9780 ( .Y(T9780_Y), .A(T16275_Y), .B(T2632_Y));
KC_NOR2_X2 T9779 ( .Y(T9779_Y), .A(T4872_Y), .B(T16267_Y));
KC_NOR2_X2 T9772 ( .Y(T9772_Y), .A(T15422_Y), .B(T15691_Y));
KC_NOR2_X2 T9754 ( .Y(T9754_Y), .A(T6768_Y), .B(T6770_Y));
KC_NOR2_X2 T9753 ( .Y(T9753_Y), .A(T6768_Y), .B(T6775_Y));
KC_NOR2_X2 T9748 ( .Y(T9748_Y), .A(T611_Y), .B(T15419_Y));
KC_NOR2_X2 T9747 ( .Y(T9747_Y), .A(T4872_Y), .B(T2068_Y));
KC_NOR2_X2 T9746 ( .Y(T9746_Y), .A(T611_Y), .B(T2454_Y));
KC_NOR2_X2 T9745 ( .Y(T9745_Y), .A(T15419_Y), .B(T634_Y));
KC_NOR2_X2 T9744 ( .Y(T9744_Y), .A(T610_Y), .B(T2478_Y));
KC_NOR2_X2 T9743 ( .Y(T9743_Y), .A(T15442_Y), .B(T2466_Y));
KC_NOR2_X2 T16165 ( .Y(T16165_Y), .A(T2861_Y), .B(T2505_Y));
KC_NOR2_X2 T9874 ( .Y(T9874_Y), .A(T10941_Y), .B(T16267_Y));
KC_NOR2_X2 T9854 ( .Y(T9854_Y), .A(T10942_Y), .B(T2632_Y));
KC_NOR2_X2 T10518 ( .Y(T10518_Y), .A(T2584_Q), .B(T2570_Q));
KC_NOR2_X2 T10517 ( .Y(T10517_Y), .A(T2575_Q), .B(T2571_Q));
KC_NOR2_X2 T9957 ( .Y(T9957_Y), .A(T10239_Y), .B(T1114_Y));
KC_NOR2_X2 T9946 ( .Y(T9946_Y), .A(T1114_Y), .B(T2549_Y));
KC_NOR2_X2 T16294 ( .Y(T16294_Y), .A(T15518_Y), .B(T10064_Y));
KC_NOR2_X2 T10103 ( .Y(T10103_Y), .A(T10100_Y), .B(T10090_Y));
KC_NOR2_X2 T10102 ( .Y(T10102_Y), .A(T10101_Y), .B(T10104_Y));
KC_NOR2_X2 T10101 ( .Y(T10101_Y), .A(T9967_Y), .B(T1499_Y));
KC_NOR2_X2 T10100 ( .Y(T10100_Y), .A(T2844_Q), .B(T2597_Y));
KC_NOR2_X2 T10091 ( .Y(T10091_Y), .A(T2550_Y), .B(T10058_Y));
KC_NOR2_X2 T10090 ( .Y(T10090_Y), .A(T1509_Y), .B(T2598_Y));
KC_NOR2_X2 T10061 ( .Y(T10061_Y), .A(T2623_Y), .B(T15501_Y));
KC_NOR2_X2 T10060 ( .Y(T10060_Y), .A(T16411_Y), .B(T15503_Y));
KC_NOR2_X2 T10059 ( .Y(T10059_Y), .A(T2611_Y), .B(T15518_Y));
KC_NOR2_X2 T10058 ( .Y(T10058_Y), .A(T10517_Y), .B(T12090_Y));
KC_NOR2_X2 T10057 ( .Y(T10057_Y), .A(T2842_Q), .B(T2631_Q));
KC_NOR2_X2 T10203 ( .Y(T10203_Y), .A(T16236_Y), .B(T2643_Y));
KC_NOR2_X2 T10195 ( .Y(T10195_Y), .A(T4898_Y), .B(T15535_Y));
KC_NOR2_X2 T10188 ( .Y(T10188_Y), .A(T2064_Y), .B(T2066_Y));
KC_NOR2_X2 T10180 ( .Y(T10180_Y), .A(T15533_Y), .B(T1546_Y));
KC_NOR2_X2 T16160 ( .Y(T16160_Y), .A(T2661_Y), .B(T2652_Y));
KC_NOR2_X2 T10279 ( .Y(T10279_Y), .A(T10274_Y), .B(T10275_Y));
KC_NOR2_X2 T10278 ( .Y(T10278_Y), .A(T5754_Y), .B(T5018_Q));
KC_NOR2_X2 T10277 ( .Y(T10277_Y), .A(T5018_Q), .B(T5576_Q));
KC_NOR2_X2 T10276 ( .Y(T10276_Y), .A(T11960_Y), .B(T10273_Y));
KC_NOR2_X2 T10275 ( .Y(T10275_Y), .A(T2661_Y), .B(T2655_Y));
KC_NOR2_X2 T10274 ( .Y(T10274_Y), .A(T2653_Y), .B(T2664_Y));
KC_NOR2_X2 T10273 ( .Y(T10273_Y), .A(T2655_Y), .B(T2664_Y));
KC_NOR2_X2 T10272 ( .Y(T10272_Y), .A(T10275_Y), .B(T10270_Y));
KC_NOR2_X2 T10271 ( .Y(T10271_Y), .A(T2662_Y), .B(T2655_Y));
KC_NOR2_X2 T10270 ( .Y(T10270_Y), .A(T2652_Y), .B(T2662_Y));
KC_NOR2_X2 T10252 ( .Y(T10252_Y), .A(T2653_Y), .B(T2663_Y));
KC_NOR2_X2 T10251 ( .Y(T10251_Y), .A(T5717_Y), .B(T2652_Y));
KC_NOR2_X2 T10250 ( .Y(T10250_Y), .A(T15827_Y), .B(T2665_Y));
KC_NOR2_X2 T10249 ( .Y(T10249_Y), .A(T2652_Y), .B(T2663_Y));
KC_NOR2_X2 T10244 ( .Y(T10244_Y), .A(T2653_Y), .B(T2662_Y));
KC_NOR2_X2 T10243 ( .Y(T10243_Y), .A(T2661_Y), .B(T2653_Y));
KC_NOR2_X2 T10242 ( .Y(T10242_Y), .A(T2652_Y), .B(T2664_Y));
KC_NOR2_X2 T10241 ( .Y(T10241_Y), .A(T2652_Y), .B(T2663_Y));
KC_NOR2_X2 T15849 ( .Y(T15849_Y), .A(T14525_Q), .B(T2681_Y));
KC_NOR2_X2 T11964 ( .Y(T11964_Y), .A(T2664_Y), .B(T10281_Y));
KC_NOR2_X2 T11963 ( .Y(T11963_Y), .A(T5766_Y), .B(T2675_Y));
KC_NOR2_X2 T11362 ( .Y(T11362_Y), .A(T14537_Q), .B(T2788_Y));
KC_NOR2_X2 T11343 ( .Y(T11343_Y), .A(T14536_Q), .B(T14535_Q));
KC_NOR2_X2 T11342 ( .Y(T11342_Y), .A(T14533_Q), .B(T5786_Y));
KC_NOR2_X2 T11341 ( .Y(T11341_Y), .A(T14954_Q), .B(T2677_Y));
KC_NOR2_X2 T11321 ( .Y(T11321_Y), .A(T14527_Q), .B(T2698_Y));
KC_NOR2_X2 T11431 ( .Y(T11431_Y), .A(T16082_Q), .B(T11414_Y));
KC_NOR2_X2 T11414 ( .Y(T11414_Y), .A(T10887_Y), .B(T2701_Y));
KC_NOR2_X2 T11397 ( .Y(T11397_Y), .A(T12163_Y), .B(T6095_Y));
KC_NOR2_X2 T11472 ( .Y(T11472_Y), .A(T2778_Y), .B(T10245_Y));
KC_NOR2_X2 T11464 ( .Y(T11464_Y), .A(T5380_Q), .B(T2719_Y));
KC_NOR2_X2 T11463 ( .Y(T11463_Y), .A(T2778_Y), .B(T15882_Y));
KC_NOR2_X2 T11449 ( .Y(T11449_Y), .A(T15853_Y), .B(T15796_Q));
KC_NOR2_X2 T11448 ( .Y(T11448_Y), .A(T2729_Y), .B(T2732_Y));
KC_NOR2_X2 T10643 ( .Y(T10643_Y), .A(T2777_Y), .B(T16474_Y));
KC_NOR2_X2 T10641 ( .Y(T10641_Y), .A(T10949_Y), .B(T16474_Y));
KC_NOR2_X2 T10640 ( .Y(T10640_Y), .A(T10949_Y), .B(T2719_Y));
KC_NOR2_X2 T11527 ( .Y(T11527_Y), .A(T2777_Y), .B(T15882_Y));
KC_NOR2_X2 T11499 ( .Y(T11499_Y), .A(T5070_Y), .B(T3354_Y));
KC_NOR2_X2 T11498 ( .Y(T11498_Y), .A(T2777_Y), .B(T10245_Y));
KC_NOR2_X2 T11491 ( .Y(T11491_Y), .A(T2778_Y), .B(T2751_Y));
KC_NOR2_X2 T11490 ( .Y(T11490_Y), .A(T2778_Y), .B(T16474_Y));
KC_NOR2_X2 T11489 ( .Y(T11489_Y), .A(T10949_Y), .B(T15855_Y));
KC_NOR2_X2 T11488 ( .Y(T11488_Y), .A(T3311_Y), .B(T2763_Y));
KC_NOR2_X2 T11480 ( .Y(T11480_Y), .A(T16035_Y), .B(T3355_Y));
KC_NOR2_X2 T11479 ( .Y(T11479_Y), .A(T2778_Y), .B(T15858_Y));
KC_NOR2_X2 T11593 ( .Y(T11593_Y), .A(T13140_Q), .B(T13141_Q));
KC_NOR2_X2 T11582 ( .Y(T11582_Y), .A(T10949_Y), .B(T15881_Y));
KC_NOR2_X2 T11581 ( .Y(T11581_Y), .A(T2777_Y), .B(T15912_Y));
KC_NOR2_X2 T11580 ( .Y(T11580_Y), .A(T10949_Y), .B(T15912_Y));
KC_NOR2_X2 T11567 ( .Y(T11567_Y), .A(T2777_Y), .B(T15855_Y));
KC_NOR2_X2 T11566 ( .Y(T11566_Y), .A(T2778_Y), .B(T15856_Y));
KC_NOR2_X2 T11565 ( .Y(T11565_Y), .A(T10949_Y), .B(T15856_Y));
KC_NOR2_X2 T11564 ( .Y(T11564_Y), .A(T2778_Y), .B(T15881_Y));
KC_NOR2_X2 T11563 ( .Y(T11563_Y), .A(T10949_Y), .B(T10245_Y));
KC_NOR2_X2 T11562 ( .Y(T11562_Y), .A(T2777_Y), .B(T15856_Y));
KC_NOR2_X2 T11548 ( .Y(T11548_Y), .A(T2778_Y), .B(T15855_Y));
KC_NOR2_X2 T11547 ( .Y(T11547_Y), .A(T2793_Q), .B(T2794_Q));
KC_NOR2_X2 T11620 ( .Y(T11620_Y), .A(T2803_Y), .B(T6511_Y));
KC_NOR2_X2 T11604 ( .Y(T11604_Y), .A(T6555_Q), .B(T3355_Y));
KC_NOR2_X2 T12047 ( .Y(T12047_Y), .A(T16148_Y), .B(T6182_Y));
KC_NOR2_X2 T12046 ( .Y(T12046_Y), .A(T10966_Y), .B(T3415_Y));
KC_NOR2_X2 T11679 ( .Y(T11679_Y), .A(T2854_Y), .B(T6399_Y));
KC_NOR2_X2 T11666 ( .Y(T11666_Y), .A(T2630_Y), .B(T3412_Q));
KC_NOR2_X2 T11651 ( .Y(T11651_Y), .A(T2841_Q), .B(T11660_Y));
KC_NOR2_X2 T11650 ( .Y(T11650_Y), .A(T8351_Y), .B(T3388_Y));
KC_NOR2_X2 T11633 ( .Y(T11633_Y), .A(T12297_Y), .B(T3402_Y));
KC_NOR2_X2 T11632 ( .Y(T11632_Y), .A(T3423_Y), .B(T5999_Y));
KC_NOR2_X2 T11731 ( .Y(T11731_Y), .A(T2822_Y), .B(T2868_Y));
KC_NOR2_X2 T11730 ( .Y(T11730_Y), .A(T8352_Q), .B(T16082_Q));
KC_NOR2_X2 T11729 ( .Y(T11729_Y), .A(T12317_Y), .B(T3530_Y));
KC_NOR2_X2 T11728 ( .Y(T11728_Y), .A(T2838_Y), .B(T11729_Y));
KC_NOR2_X2 T11727 ( .Y(T11727_Y), .A(T2854_Y), .B(T12064_Y));
KC_NOR2_X2 T10623 ( .Y(T10623_Y), .A(T2906_Y), .B(T11743_Y));
KC_NOR2_X2 T10622 ( .Y(T10622_Y), .A(T6139_Y), .B(T12048_Y));
KC_NOR2_X2 T10607 ( .Y(T10607_Y), .A(T5523_Y), .B(T4015_Y));
KC_NOR2_X2 T10595 ( .Y(T10595_Y), .A(T16132_Y), .B(T2890_Y));
KC_NOR2_X2 T10594 ( .Y(T10594_Y), .A(T2879_Y), .B(T2890_Y));
KC_NOR2_X2 T10593 ( .Y(T10593_Y), .A(T2838_Y), .B(T6208_Y));
KC_NOR2_X2 T10592 ( .Y(T10592_Y), .A(T2865_Y), .B(T3514_Y));
KC_NOR2_X2 T10589 ( .Y(T10589_Y), .A(T12038_Y), .B(T5523_Y));
KC_NOR2_X2 T10572 ( .Y(T10572_Y), .A(T2877_Y), .B(T12060_Y));
KC_NOR2_X2 T10569 ( .Y(T10569_Y), .A(T12064_Y), .B(T3426_Y));
KC_NOR2_X2 T11810 ( .Y(T11810_Y), .A(T12105_Y), .B(T4999_Y));
KC_NOR2_X2 T11809 ( .Y(T11809_Y), .A(T2910_Y), .B(T2917_Y));
KC_NOR2_X2 T11808 ( .Y(T11808_Y), .A(T5515_Y), .B(T6573_Y));
KC_NOR2_X2 T11771 ( .Y(T11771_Y), .A(T12103_Y), .B(T2898_Y));
KC_NOR2_X2 T11770 ( .Y(T11770_Y), .A(T11771_Y), .B(T6222_Y));
KC_NOR2_X2 T11769 ( .Y(T11769_Y), .A(T2918_Y), .B(T6190_Y));
KC_NOR2_X2 T11747 ( .Y(T11747_Y), .A(T15633_Y), .B(T16130_Y));
KC_NOR2_X2 T11746 ( .Y(T11746_Y), .A(T2948_Y), .B(T4054_Y));
KC_NOR2_X2 T11745 ( .Y(T11745_Y), .A(T2938_Y), .B(T10881_Y));
KC_NOR2_X2 T11744 ( .Y(T11744_Y), .A(T2936_Y), .B(T4096_Y));
KC_NOR2_X2 T11743 ( .Y(T11743_Y), .A(T2918_Y), .B(T6192_Y));
KC_NOR2_X2 T11742 ( .Y(T11742_Y), .A(T2952_Q), .B(T2911_Y));
KC_NOR2_X2 T11741 ( .Y(T11741_Y), .A(T2911_Y), .B(T6195_Y));
KC_NOR2_X2 T11739 ( .Y(T11739_Y), .A(T10977_Y), .B(T6192_Y));
KC_NOR2_X2 T11043 ( .Y(T11043_Y), .A(T2941_Y), .B(T4055_Y));
KC_NOR2_X2 T11042 ( .Y(T11042_Y), .A(T6531_Y), .B(T4055_Y));
KC_NOR2_X2 T11041 ( .Y(T11041_Y), .A(T2948_Y), .B(T290_Y));
KC_NOR2_X2 T11037 ( .Y(T11037_Y), .A(T4096_Y), .B(T2938_Y));
KC_NOR2_X2 T10555 ( .Y(T10555_Y), .A(T6578_Y), .B(T6222_Y));
KC_NOR2_X2 T10554 ( .Y(T10554_Y), .A(T10561_Y), .B(T6582_Y));
KC_NOR2_X2 T10553 ( .Y(T10553_Y), .A(T10547_Y), .B(T3514_Y));
KC_NOR2_X2 T10552 ( .Y(T10552_Y), .A(T6582_Y), .B(T10559_Y));
KC_NOR2_X2 T11846 ( .Y(T11846_Y), .A(T2943_Q), .B(T2944_Q));
KC_NOR2_X2 T11844 ( .Y(T11844_Y), .A(T6516_Y), .B(T6491_Y));
KC_NOR2_X2 T11837 ( .Y(T11837_Y), .A(T6509_Y), .B(T2934_Y));
KC_NOR2_X2 T11836 ( .Y(T11836_Y), .A(T11002_Y), .B(T11005_Y));
KC_NOR2_X2 T11823 ( .Y(T11823_Y), .A(T15643_Y), .B(T2959_Y));
KC_NOR2_X2 T11822 ( .Y(T11822_Y), .A(T5540_Y), .B(T6537_Y));
KC_NOR2_X2 T10436 ( .Y(T10436_Y), .A(T3014_Y), .B(T9651_Y));
KC_NOR2_X2 T9669 ( .Y(T9669_Y), .A(T2448_Y), .B(T3020_Y));
KC_NOR2_X2 T9668 ( .Y(T9668_Y), .A(T15422_Y), .B(T483_Y));
KC_NOR2_X2 T9664 ( .Y(T9664_Y), .A(T475_Y), .B(T9651_Y));
KC_NOR2_X2 T9655 ( .Y(T9655_Y), .A(T5080_Y), .B(T2448_Y));
KC_NOR2_X2 T9654 ( .Y(T9654_Y), .A(T15422_Y), .B(T15403_Y));
KC_NOR2_X2 T9636 ( .Y(T9636_Y), .A(T3014_Y), .B(T9649_Y));
KC_NOR2_X2 T8526 ( .Y(T8526_Y), .A(T15422_Y), .B(T6761_Y));
KC_NOR2_X2 T631 ( .Y(T631_Y), .A(T602_Y), .B(T9736_Y));
KC_NOR2_X2 T9768 ( .Y(T9768_Y), .A(T3051_Y), .B(T9736_Y));
KC_NOR2_X2 T9767 ( .Y(T9767_Y), .A(T3621_Y), .B(T9769_Y));
KC_NOR2_X2 T9765 ( .Y(T9765_Y), .A(T602_Y), .B(T9737_Y));
KC_NOR2_X2 T9739 ( .Y(T9739_Y), .A(T15032_Y), .B(T16265_Y));
KC_NOR2_X2 T9732 ( .Y(T9732_Y), .A(T3051_Y), .B(T9738_Y));
KC_NOR2_X2 T9731 ( .Y(T9731_Y), .A(T602_Y), .B(T9738_Y));
KC_NOR2_X2 T9730 ( .Y(T9730_Y), .A(T3051_Y), .B(T9737_Y));
KC_NOR2_X2 T9878 ( .Y(T9878_Y), .A(T5026_Y), .B(T16405_Y));
KC_NOR2_X2 T9839 ( .Y(T9839_Y), .A(T5026_Y), .B(T872_Y));
KC_NOR2_X2 T16442 ( .Y(T16442_Y), .A(T16403_Y), .B(T10505_Y));
KC_NOR2_X2 T9937 ( .Y(T9937_Y), .A(T3712_Y), .B(T10506_Y));
KC_NOR2_X2 T10268 ( .Y(T10268_Y), .A(T14950_Q), .B(T5077_Y));
KC_NOR2_X2 T10267 ( .Y(T10267_Y), .A(T5748_Y), .B(T6014_Y));
KC_NOR2_X2 T10266 ( .Y(T10266_Y), .A(T14515_Q), .B(T14516_Q));
KC_NOR2_X2 T10265 ( .Y(T10265_Y), .A(T14520_Q), .B(T10268_Y));
KC_NOR2_X2 T11988 ( .Y(T11988_Y), .A(T11977_Y), .B(T11370_Y));
KC_NOR2_X2 T11987 ( .Y(T11987_Y), .A(T3840_Y), .B(T5816_Y));
KC_NOR2_X2 T11959 ( .Y(T11959_Y), .A(T16160_Y), .B(T2660_Y));
KC_NOR2_X2 T11358 ( .Y(T11358_Y), .A(T15007_Y), .B(T3202_Y));
KC_NOR2_X2 T11357 ( .Y(T11357_Y), .A(T14526_Q), .B(T5784_Y));
KC_NOR2_X2 T11356 ( .Y(T11356_Y), .A(T13079_Q), .B(T4381_Q));
KC_NOR2_X2 T11355 ( .Y(T11355_Y), .A(T13067_Q), .B(T13079_Q));
KC_NOR2_X2 T11337 ( .Y(T11337_Y), .A(T11355_Y), .B(T5774_Y));
KC_NOR2_X2 T11325 ( .Y(T11325_Y), .A(T3840_Y), .B(T3816_Y));
KC_NOR2_X2 T11320 ( .Y(T11320_Y), .A(T5428_Q), .B(T3213_Q));
KC_NOR2_X2 T11413 ( .Y(T11413_Y), .A(T14546_Q), .B(T11412_Y));
KC_NOR2_X2 T11412 ( .Y(T11412_Y), .A(T14544_Q), .B(T15010_Y));
KC_NOR2_X2 T11411 ( .Y(T11411_Y), .A(T3855_Y), .B(T6109_Y));
KC_NOR2_X2 T11460 ( .Y(T11460_Y), .A(T3253_Y), .B(T11459_Y));
KC_NOR2_X2 T11459 ( .Y(T11459_Y), .A(T3269_Y), .B(T3253_Y));
KC_NOR2_X2 T11458 ( .Y(T11458_Y), .A(T2777_Y), .B(T2751_Y));
KC_NOR2_X2 T11457 ( .Y(T11457_Y), .A(T2777_Y), .B(T2719_Y));
KC_NOR2_X2 T11456 ( .Y(T11456_Y), .A(T2778_Y), .B(T15857_Y));
KC_NOR2_X2 T11455 ( .Y(T11455_Y), .A(T2778_Y), .B(T15854_Y));
KC_NOR2_X2 T10642 ( .Y(T10642_Y), .A(T10949_Y), .B(T15854_Y));
KC_NOR2_X2 T10639 ( .Y(T10639_Y), .A(T2777_Y), .B(T15854_Y));
KC_NOR2_X2 T10638 ( .Y(T10638_Y), .A(T2777_Y), .B(T15857_Y));
KC_NOR2_X2 T10637 ( .Y(T10637_Y), .A(T10949_Y), .B(T2751_Y));
KC_NOR2_X2 T11526 ( .Y(T11526_Y), .A(T5022_Y), .B(T5939_Y));
KC_NOR2_X2 T11525 ( .Y(T11525_Y), .A(T10949_Y), .B(T15857_Y));
KC_NOR2_X2 T11515 ( .Y(T11515_Y), .A(T2777_Y), .B(T2127_Y));
KC_NOR2_X2 T11497 ( .Y(T11497_Y), .A(T2778_Y), .B(T2719_Y));
KC_NOR2_X2 T11487 ( .Y(T11487_Y), .A(T3314_Y), .B(T3292_Y));
KC_NOR2_X2 T11477 ( .Y(T11477_Y), .A(T2778_Y), .B(T15853_Y));
KC_NOR2_X2 T15984 ( .Y(T15984_Y), .A(T10949_Y), .B(T1748_Y));
KC_NOR2_X2 T15981 ( .Y(T15981_Y), .A(T2777_Y), .B(T15881_Y));
KC_NOR2_X2 T11592 ( .Y(T11592_Y), .A(T12826_Y), .B(T3320_Y));
KC_NOR2_X2 T11579 ( .Y(T11579_Y), .A(T2778_Y), .B(T1748_Y));
KC_NOR2_X2 T11578 ( .Y(T11578_Y), .A(T2777_Y), .B(T1748_Y));
KC_NOR2_X2 T11561 ( .Y(T11561_Y), .A(T10949_Y), .B(T15895_Y));
KC_NOR2_X2 T11560 ( .Y(T11560_Y), .A(T2778_Y), .B(T2127_Y));
KC_NOR2_X2 T11559 ( .Y(T11559_Y), .A(T10949_Y), .B(T2127_Y));
KC_NOR2_X2 T11558 ( .Y(T11558_Y), .A(T10949_Y), .B(T15858_Y));
KC_NOR2_X2 T11545 ( .Y(T11545_Y), .A(T2778_Y), .B(T15912_Y));
KC_NOR2_X2 T11603 ( .Y(T11603_Y), .A(T16035_Y), .B(T5070_Y));
KC_NOR2_X2 T11597 ( .Y(T11597_Y), .A(T5896_Y), .B(T6046_Y));
KC_NOR2_X2 T6049 ( .Y(T6049_Y), .A(T16039_Y), .B(T11628_Y));
KC_NOR2_X2 T12044 ( .Y(T12044_Y), .A(T16103_Y), .B(T16149_Y));
KC_NOR2_X2 T12043 ( .Y(T12043_Y), .A(T16039_Y), .B(T12322_Y));
KC_NOR2_X2 T12004 ( .Y(T12004_Y), .A(T16036_Y), .B(T4036_Y));
KC_NOR2_X2 T12003 ( .Y(T12003_Y), .A(T5525_Q), .B(T16031_Y));
KC_NOR2_X2 T12002 ( .Y(T12002_Y), .A(T3359_Y), .B(T16139_Y));
KC_NOR2_X2 T11677 ( .Y(T11677_Y), .A(T6083_Y), .B(T4021_Y));
KC_NOR2_X2 T11676 ( .Y(T11676_Y), .A(T15616_Y), .B(T10584_Y));
KC_NOR2_X2 T11675 ( .Y(T11675_Y), .A(T6560_Y), .B(T16103_Y));
KC_NOR2_X2 T11674 ( .Y(T11674_Y), .A(T6086_Y), .B(T3378_Y));
KC_NOR2_X2 T11664 ( .Y(T11664_Y), .A(T3383_Y), .B(T3468_Y));
KC_NOR2_X2 T11663 ( .Y(T11663_Y), .A(T5522_Y), .B(T10964_Y));
KC_NOR2_X2 T11662 ( .Y(T11662_Y), .A(T2841_Q), .B(T6087_Y));
KC_NOR2_X2 T11661 ( .Y(T11661_Y), .A(T3394_Y), .B(T4031_Y));
KC_NOR2_X2 T11660 ( .Y(T11660_Y), .A(T11818_Y), .B(T16102_Y));
KC_NOR2_X2 T11658 ( .Y(T11658_Y), .A(T4024_Y), .B(T3389_Y));
KC_NOR2_X2 T11647 ( .Y(T11647_Y), .A(T3355_Y), .B(T4034_Y));
KC_NOR2_X2 T11646 ( .Y(T11646_Y), .A(T3362_Y), .B(T3394_Y));
KC_NOR2_X2 T11645 ( .Y(T11645_Y), .A(T11639_Y), .B(T11642_Y));
KC_NOR2_X2 T11644 ( .Y(T11644_Y), .A(T10962_Y), .B(T4034_Y));
KC_NOR2_X2 T11643 ( .Y(T11643_Y), .A(T4035_Y), .B(T3393_Y));
KC_NOR2_X2 T11642 ( .Y(T11642_Y), .A(T4034_Y), .B(T3400_Y));
KC_NOR2_X2 T11641 ( .Y(T11641_Y), .A(T16035_Y), .B(T3394_Y));
KC_NOR2_X2 T11639 ( .Y(T11639_Y), .A(T10963_Y), .B(T4033_Y));
KC_NOR2_X2 T11631 ( .Y(T11631_Y), .A(T2848_Y), .B(T3411_Y));
KC_NOR2_X2 T11630 ( .Y(T11630_Y), .A(T16036_Y), .B(T15760_Q));
KC_NOR2_X2 T8502 ( .Y(T8502_Y), .A(T2865_Y), .B(T6179_Y));
KC_NOR2_X2 T11725 ( .Y(T11725_Y), .A(T3429_Y), .B(T2879_Y));
KC_NOR2_X2 T11724 ( .Y(T11724_Y), .A(T2865_Y), .B(T4104_Y));
KC_NOR2_X2 T10624 ( .Y(T10624_Y), .A(T6067_Y), .B(T3445_Y));
KC_NOR2_X2 T10620 ( .Y(T10620_Y), .A(T3429_Y), .B(T4015_Y));
KC_NOR2_X2 T10619 ( .Y(T10619_Y), .A(T10620_Y), .B(T11716_Y));
KC_NOR2_X2 T10608 ( .Y(T10608_Y), .A(T15621_Y), .B(T16104_Y));
KC_NOR2_X2 T10606 ( .Y(T10606_Y), .A(T3394_Y), .B(T11027_Y));
KC_NOR2_X2 T10590 ( .Y(T10590_Y), .A(T3515_Y), .B(T2910_Y));
KC_NOR2_X2 T10587 ( .Y(T10587_Y), .A(T6119_Y), .B(T3439_Y));
KC_NOR2_X2 T10585 ( .Y(T10585_Y), .A(T15636_Y), .B(T4083_Y));
KC_NOR2_X2 T10584 ( .Y(T10584_Y), .A(T15636_Y), .B(T16141_Y));
KC_NOR2_X2 T10581 ( .Y(T10581_Y), .A(T2865_Y), .B(T6119_Y));
KC_NOR2_X2 T10571 ( .Y(T10571_Y), .A(T6106_Y), .B(T6039_Y));
KC_NOR2_X2 T10570 ( .Y(T10570_Y), .A(T4051_Q), .B(T6145_Y));
KC_NOR2_X2 T10568 ( .Y(T10568_Y), .A(T10606_Y), .B(T3443_Y));
KC_NOR2_X2 T11804 ( .Y(T11804_Y), .A(T12322_Y), .B(T6080_Y));
KC_NOR2_X2 T11803 ( .Y(T11803_Y), .A(T2906_Y), .B(T11801_Y));
KC_NOR2_X2 T11802 ( .Y(T11802_Y), .A(T15234_Y), .B(T12464_Y));
KC_NOR2_X2 T11801 ( .Y(T11801_Y), .A(T5522_Y), .B(T3473_Y));
KC_NOR2_X2 T11782 ( .Y(T11782_Y), .A(T6236_Y), .B(T3427_Y));
KC_NOR2_X2 T11765 ( .Y(T11765_Y), .A(T16050_Y), .B(T6215_Y));
KC_NOR2_X2 T11764 ( .Y(T11764_Y), .A(T4178_Q), .B(T6209_Y));
KC_NOR2_X2 T10550 ( .Y(T10550_Y), .A(T16135_Y), .B(T2800_Y));
KC_NOR2_X2 T10545 ( .Y(T10545_Y), .A(T16138_Y), .B(T8361_Y));
KC_NOR2_X2 T11843 ( .Y(T11843_Y), .A(T3522_Q), .B(T6489_Y));
KC_NOR2_X2 T11835 ( .Y(T11835_Y), .A(T3520_Q), .B(T3522_Q));
KC_NOR2_X2 T11834 ( .Y(T11834_Y), .A(T3521_Q), .B(T6510_Y));
KC_NOR2_X2 T11833 ( .Y(T11833_Y), .A(T6512_Y), .B(T3506_Y));
KC_NOR2_X2 T11832 ( .Y(T11832_Y), .A(T6510_Y), .B(T3525_Q));
KC_NOR2_X2 T11818 ( .Y(T11818_Y), .A(T11007_Y), .B(T3511_Y));
KC_NOR2_X2 T11817 ( .Y(T11817_Y), .A(T2865_Y), .B(T10985_Y));
KC_NOR2_X2 T11816 ( .Y(T11816_Y), .A(T11007_Y), .B(T3508_Y));
KC_NOR2_X2 T8150 ( .Y(T8150_Y), .A(T3519_Q), .B(T3523_Q));
KC_NOR2_X2 T6482 ( .Y(T6482_Y), .A(T3608_Y), .B(T8521_Y));
KC_NOR2_X2 T9665 ( .Y(T9665_Y), .A(T15402_Y), .B(T8521_Y));
KC_NOR2_X2 T9637 ( .Y(T9637_Y), .A(T3608_Y), .B(T8520_Y));
KC_NOR2_X2 T9635 ( .Y(T9635_Y), .A(T15402_Y), .B(T8520_Y));
KC_NOR2_X2 T9764 ( .Y(T9764_Y), .A(T3621_Y), .B(T9771_Y));
KC_NOR2_X2 T9763 ( .Y(T9763_Y), .A(T607_Y), .B(T9771_Y));
KC_NOR2_X2 T9729 ( .Y(T9729_Y), .A(T607_Y), .B(T9770_Y));
KC_NOR2_X2 T9868 ( .Y(T9868_Y), .A(T3666_Y), .B(T9830_Y));
KC_NOR2_X2 T9867 ( .Y(T9867_Y), .A(T879_Y), .B(T9870_Y));
KC_NOR2_X2 T9866 ( .Y(T9866_Y), .A(T879_Y), .B(T9827_Y));
KC_NOR2_X2 T9865 ( .Y(T9865_Y), .A(T3666_Y), .B(T9827_Y));
KC_NOR2_X2 T9864 ( .Y(T9864_Y), .A(T879_Y), .B(T9830_Y));
KC_NOR2_X2 T9863 ( .Y(T9863_Y), .A(T3666_Y), .B(T9870_Y));
KC_NOR2_X2 T9862 ( .Y(T9862_Y), .A(T3667_Y), .B(T9833_Y));
KC_NOR2_X2 T9825 ( .Y(T9825_Y), .A(T3667_Y), .B(T9829_Y));
KC_NOR2_X2 T9824 ( .Y(T9824_Y), .A(T3667_Y), .B(T9828_Y));
KC_NOR2_X2 T9823 ( .Y(T9823_Y), .A(T856_Y), .B(T9828_Y));
KC_NOR2_X2 T9822 ( .Y(T9822_Y), .A(T856_Y), .B(T9833_Y));
KC_NOR2_X2 T9936 ( .Y(T9936_Y), .A(T3712_Y), .B(T10500_Y));
KC_NOR2_X2 T9932 ( .Y(T9932_Y), .A(T16403_Y), .B(T10500_Y));
KC_NOR2_X2 T11983 ( .Y(T11983_Y), .A(T4486_Y), .B(T3836_Y));
KC_NOR2_X2 T11982 ( .Y(T11982_Y), .A(T15908_Y), .B(T5800_Y));
KC_NOR2_X2 T11981 ( .Y(T11981_Y), .A(T145_Q), .B(T15907_Y));
KC_NOR2_X2 T11353 ( .Y(T11353_Y), .A(T5838_Y), .B(T3794_Y));
KC_NOR2_X2 T11352 ( .Y(T11352_Y), .A(T5780_Y), .B(T3797_Y));
KC_NOR2_X2 T11336 ( .Y(T11336_Y), .A(T16153_Y), .B(T5770_Y));
KC_NOR2_X2 T11335 ( .Y(T11335_Y), .A(T3840_Y), .B(T4436_Y));
KC_NOR2_X2 T11318 ( .Y(T11318_Y), .A(T144_Q), .B(T15907_Y));
KC_NOR2_X2 T11317 ( .Y(T11317_Y), .A(T5780_Y), .B(T5816_Y));
KC_NOR2_X2 T15897 ( .Y(T15897_Y), .A(T144_Q), .B(T4486_Y));
KC_NOR2_X2 T15888 ( .Y(T15888_Y), .A(T5802_Y), .B(T144_Q));
KC_NOR2_X2 T11428 ( .Y(T11428_Y), .A(T4487_Q), .B(T16154_Y));
KC_NOR2_X2 T11427 ( .Y(T11427_Y), .A(T4465_Q), .B(T4487_Q));
KC_NOR2_X2 T11426 ( .Y(T11426_Y), .A(T5815_Y), .B(T5788_Y));
KC_NOR2_X2 T11410 ( .Y(T11410_Y), .A(T15908_Y), .B(T16153_Y));
KC_NOR2_X2 T11409 ( .Y(T11409_Y), .A(T14494_Q), .B(T14495_Q));
KC_NOR2_X2 T11408 ( .Y(T11408_Y), .A(T15908_Y), .B(T16154_Y));
KC_NOR2_X2 T11394 ( .Y(T11394_Y), .A(T5788_Y), .B(T5801_Y));
KC_NOR2_X2 T11393 ( .Y(T11393_Y), .A(T16154_Y), .B(T5789_Y));
KC_NOR2_X2 T11381 ( .Y(T11381_Y), .A(T5789_Y), .B(T3856_Y));
KC_NOR2_X2 T11380 ( .Y(T11380_Y), .A(T5838_Y), .B(T5816_Y));
KC_NOR2_X2 T11379 ( .Y(T11379_Y), .A(T16154_Y), .B(T3849_Y));
KC_NOR2_X2 T11378 ( .Y(T11378_Y), .A(T144_Q), .B(T145_Q));
KC_NOR2_X2 T11377 ( .Y(T11377_Y), .A(T4486_Y), .B(T5803_Y));
KC_NOR2_X2 T11376 ( .Y(T11376_Y), .A(T144_Q), .B(T4487_Q));
KC_NOR2_X2 T11375 ( .Y(T11375_Y), .A(T145_Q), .B(T11969_Y));
KC_NOR2_X2 T11367 ( .Y(T11367_Y), .A(T145_Q), .B(T4487_Q));
KC_NOR2_X2 T15932 ( .Y(T15932_Y), .A(T3885_Q), .B(T5454_Y));
KC_NOR2_X2 T11444 ( .Y(T11444_Y), .A(T10923_Y), .B(T5859_Y));
KC_NOR2_X2 T10635 ( .Y(T10635_Y), .A(T3890_Q), .B(T10943_Y));
KC_NOR2_X2 T10634 ( .Y(T10634_Y), .A(T3873_Q), .B(T10943_Y));
KC_NOR2_X2 T10633 ( .Y(T10633_Y), .A(T10635_Y), .B(T10634_Y));
KC_NOR2_X2 T10632 ( .Y(T10632_Y), .A(T12208_Y), .B(T4523_Y));
KC_NOR2_X2 T11524 ( .Y(T11524_Y), .A(T5981_Y), .B(T11519_Y));
KC_NOR2_X2 T11523 ( .Y(T11523_Y), .A(T6219_Y), .B(T11519_Y));
KC_NOR2_X2 T11522 ( .Y(T11522_Y), .A(T5981_Y), .B(T11587_Y));
KC_NOR2_X2 T11505 ( .Y(T11505_Y), .A(T5457_Y), .B(T5981_Y));
KC_NOR2_X2 T11496 ( .Y(T11496_Y), .A(T15955_Y), .B(T11509_Y));
KC_NOR2_X2 T11495 ( .Y(T11495_Y), .A(T15955_Y), .B(T13124_Y));
KC_NOR2_X2 T11484 ( .Y(T11484_Y), .A(T3912_Y), .B(T5120_Y));
KC_NOR2_X2 T11483 ( .Y(T11483_Y), .A(T5120_Y), .B(T3912_Y));
KC_NOR2_X2 T11476 ( .Y(T11476_Y), .A(T3964_Q), .B(T3968_Q));
KC_NOR2_X2 T11590 ( .Y(T11590_Y), .A(T11555_Y), .B(T3946_Y));
KC_NOR2_X2 T11577 ( .Y(T11577_Y), .A(T3964_Q), .B(T3947_Y));
KC_NOR2_X2 T11576 ( .Y(T11576_Y), .A(T5973_Y), .B(T3947_Y));
KC_NOR2_X2 T11575 ( .Y(T11575_Y), .A(T8289_Y), .B(T15159_Y));
KC_NOR2_X2 T11574 ( .Y(T11574_Y), .A(T3964_Q), .B(T11576_Y));
KC_NOR2_X2 T11556 ( .Y(T11556_Y), .A(T3974_Q), .B(T3944_Y));
KC_NOR2_X2 T11543 ( .Y(T11543_Y), .A(T3974_Q), .B(T5984_Y));
KC_NOR2_X2 T11618 ( .Y(T11618_Y), .A(T4596_Y), .B(T3976_Y));
KC_NOR2_X2 T11617 ( .Y(T11617_Y), .A(T11618_Y), .B(T4589_Y));
KC_NOR2_X2 T11616 ( .Y(T11616_Y), .A(T15609_Y), .B(T3976_Y));
KC_NOR2_X2 T11615 ( .Y(T11615_Y), .A(T4606_Q), .B(T5158_Q));
KC_NOR2_X2 T11614 ( .Y(T11614_Y), .A(T11618_Y), .B(T3988_Y));
KC_NOR2_X2 T12038 ( .Y(T12038_Y), .A(T4748_Y), .B(T6077_Y));
KC_NOR2_X2 T11671 ( .Y(T11671_Y), .A(T5530_Q), .B(T6079_Y));
KC_NOR2_X2 T11659 ( .Y(T11659_Y), .A(T16035_Y), .B(T6048_Y));
KC_NOR2_X2 T11656 ( .Y(T11656_Y), .A(T5525_Q), .B(T4049_Y));
KC_NOR2_X2 T11638 ( .Y(T11638_Y), .A(T6175_Y), .B(T15760_Q));
KC_NOR2_X2 T11636 ( .Y(T11636_Y), .A(T15601_Y), .B(T13130_Q));
KC_NOR2_X2 T11626 ( .Y(T11626_Y), .A(T5530_Q), .B(T4176_Q));
KC_NOR2_X2 T11715 ( .Y(T11715_Y), .A(T4016_Y), .B(T16108_Y));
KC_NOR2_X2 T11714 ( .Y(T11714_Y), .A(T11657_Y), .B(T5056_Y));
KC_NOR2_X2 T11713 ( .Y(T11713_Y), .A(T5568_Q), .B(T15619_Y));
KC_NOR2_X2 T11712 ( .Y(T11712_Y), .A(T5135_Y), .B(T4060_Y));
KC_NOR2_X2 T11711 ( .Y(T11711_Y), .A(T10624_Y), .B(T3406_Y));
KC_NOR2_X2 T11710 ( .Y(T11710_Y), .A(T4106_Y), .B(T16051_Y));
KC_NOR2_X2 T11709 ( .Y(T11709_Y), .A(T11636_Y), .B(T2849_Y));
KC_NOR2_X2 T10618 ( .Y(T10618_Y), .A(T4071_Y), .B(T12281_Y));
KC_NOR2_X2 T10617 ( .Y(T10617_Y), .A(T5568_Q), .B(T5135_Y));
KC_NOR2_X2 T10616 ( .Y(T10616_Y), .A(T10617_Y), .B(T4068_Y));
KC_NOR2_X2 T10615 ( .Y(T10615_Y), .A(T6155_Y), .B(T6106_Y));
KC_NOR2_X2 T10605 ( .Y(T10605_Y), .A(T6046_Y), .B(T5056_Y));
KC_NOR2_X2 T10604 ( .Y(T10604_Y), .A(T6157_Y), .B(T4060_Y));
KC_NOR2_X2 T10602 ( .Y(T10602_Y), .A(T4095_Y), .B(T10616_Y));
KC_NOR2_X2 T10586 ( .Y(T10586_Y), .A(T10617_Y), .B(T3515_Y));
KC_NOR2_X2 T10582 ( .Y(T10582_Y), .A(T6112_Y), .B(T6098_Y));
KC_NOR2_X2 T10579 ( .Y(T10579_Y), .A(T8385_Y), .B(T10577_Y));
KC_NOR2_X2 T10578 ( .Y(T10578_Y), .A(T4087_Y), .B(T3459_Y));
KC_NOR2_X2 T10577 ( .Y(T10577_Y), .A(T4083_Y), .B(T6107_Y));
KC_NOR2_X2 T10567 ( .Y(T10567_Y), .A(T6610_S), .B(T4093_Y));
KC_NOR2_X2 T10566 ( .Y(T10566_Y), .A(T4083_Y), .B(T4073_Y));
KC_NOR2_X2 T10565 ( .Y(T10565_Y), .A(T8385_Y), .B(T4102_Y));
KC_NOR2_X2 T10564 ( .Y(T10564_Y), .A(T11715_Y), .B(T6157_Y));
KC_NOR2_X2 T11796 ( .Y(T11796_Y), .A(T11795_Y), .B(T11804_Y));
KC_NOR2_X2 T11795 ( .Y(T11795_Y), .A(T6119_Y), .B(T10580_Y));
KC_NOR2_X2 T11781 ( .Y(T11781_Y), .A(T5051_Y), .B(T3427_Y));
KC_NOR2_X2 T11736 ( .Y(T11736_Y), .A(T4171_Q), .B(T4169_Q));
KC_NOR2_X2 T10543 ( .Y(T10543_Y), .A(T6155_Y), .B(T4091_Y));
KC_NOR2_X2 T11842 ( .Y(T11842_Y), .A(T9163_Y), .B(T2708_Y));
KC_NOR2_X2 T11830 ( .Y(T11830_Y), .A(T4168_Q), .B(T11001_Y));
KC_NOR2_X2 T11814 ( .Y(T11814_Y), .A(T8424_Y), .B(T4148_Y));
KC_NOR2_X2 T11813 ( .Y(T11813_Y), .A(T4163_Q), .B(T4119_Y));
KC_NOR2_X2 T9858 ( .Y(T9858_Y), .A(T12785_Y), .B(T422_Y));
KC_NOR2_X2 T10115 ( .Y(T10115_Y), .A(T3728_Y), .B(T3070_Y));
KC_NOR2_X2 T10246 ( .Y(T10246_Y), .A(T4376_Q), .B(T3185_Y));
KC_NOR2_X2 T11975 ( .Y(T11975_Y), .A(T13305_Y), .B(T11974_Y));
KC_NOR2_X2 T11349 ( .Y(T11349_Y), .A(T14942_Q), .B(T15907_Y));
KC_NOR2_X2 T11348 ( .Y(T11348_Y), .A(T11347_Y), .B(T5838_Y));
KC_NOR2_X2 T11347 ( .Y(T11347_Y), .A(T5777_Y), .B(T11349_Y));
KC_NOR2_X2 T11322 ( .Y(T11322_Y), .A(T3794_Y), .B(T4394_Y));
KC_NOR2_X2 T11313 ( .Y(T11313_Y), .A(T5830_Y), .B(T11310_Y));
KC_NOR2_X2 T11312 ( .Y(T11312_Y), .A(T4487_Q), .B(T4448_Y));
KC_NOR2_X2 T11422 ( .Y(T11422_Y), .A(T3850_Y), .B(T4445_Y));
KC_NOR2_X2 T11421 ( .Y(T11421_Y), .A(T145_Q), .B(T16153_Y));
KC_NOR2_X2 T11402 ( .Y(T11402_Y), .A(T16153_Y), .B(T4486_Y));
KC_NOR2_X2 T11401 ( .Y(T11401_Y), .A(T4457_Y), .B(T4439_Y));
KC_NOR2_X2 T11389 ( .Y(T11389_Y), .A(T3825_Y), .B(T4439_Y));
KC_NOR2_X2 T11372 ( .Y(T11372_Y), .A(T5802_Y), .B(T4448_Y));
KC_NOR2_X2 T11371 ( .Y(T11371_Y), .A(T4457_Y), .B(T3856_Y));
KC_NOR2_X2 T11370 ( .Y(T11370_Y), .A(T5800_Y), .B(T4394_Y));
KC_NOR2_X2 T11365 ( .Y(T11365_Y), .A(T5815_Y), .B(T5787_Y));
KC_NOR2_X2 T11466 ( .Y(T11466_Y), .A(T15572_Y), .B(T5873_Y));
KC_NOR2_X2 T11454 ( .Y(T11454_Y), .A(T4483_Y), .B(T15570_Y));
KC_NOR2_X2 T11453 ( .Y(T11453_Y), .A(T10924_Y), .B(T5862_Y));
KC_NOR2_X2 T11452 ( .Y(T11452_Y), .A(T2757_Y), .B(T12354_Y));
KC_NOR2_X2 T11451 ( .Y(T11451_Y), .A(T4474_Y), .B(T5141_Y));
KC_NOR2_X2 T11442 ( .Y(T11442_Y), .A(T14550_Q), .B(T14548_Q));
KC_NOR2_X2 T11433 ( .Y(T11433_Y), .A(T14547_Q), .B(T10922_Y));
KC_NOR2_X2 T10629 ( .Y(T10629_Y), .A(T5932_Y), .B(T15935_Y));
KC_NOR2_X2 T10628 ( .Y(T10628_Y), .A(T15935_Y), .B(T4472_Y));
KC_NOR2_X2 T11521 ( .Y(T11521_Y), .A(T4493_Q), .B(T4601_Y));
KC_NOR2_X2 T11520 ( .Y(T11520_Y), .A(T4489_Y), .B(T5929_Y));
KC_NOR2_X2 T11519 ( .Y(T11519_Y), .A(T4506_Y), .B(T4472_Y));
KC_NOR2_X2 T11508 ( .Y(T11508_Y), .A(T4527_Q), .B(T5139_Y));
KC_NOR2_X2 T11507 ( .Y(T11507_Y), .A(T4527_Q), .B(T4526_Q));
KC_NOR2_X2 T11506 ( .Y(T11506_Y), .A(T5914_Y), .B(T4560_Y));
KC_NOR2_X2 T11475 ( .Y(T11475_Y), .A(T4528_Q), .B(T15706_Y));
KC_NOR2_X2 T12015 ( .Y(T12015_Y), .A(T5157_Y), .B(T4545_Y));
KC_NOR2_X2 T12014 ( .Y(T12014_Y), .A(T4576_Q), .B(T5952_Y));
KC_NOR2_X2 T11589 ( .Y(T11589_Y), .A(T2757_Y), .B(T12232_Y));
KC_NOR2_X2 T11588 ( .Y(T11588_Y), .A(T5914_Y), .B(T5149_Y));
KC_NOR2_X2 T11587 ( .Y(T11587_Y), .A(T4551_Y), .B(T5914_Y));
KC_NOR2_X2 T11573 ( .Y(T11573_Y), .A(T4570_Y), .B(T15988_Y));
KC_NOR2_X2 T11572 ( .Y(T11572_Y), .A(T4570_Y), .B(T15988_Y));
KC_NOR2_X2 T11570 ( .Y(T11570_Y), .A(T12015_Y), .B(T4550_Y));
KC_NOR2_X2 T11555 ( .Y(T11555_Y), .A(T4577_Y), .B(T4561_Y));
KC_NOR2_X2 T11554 ( .Y(T11554_Y), .A(T11536_Y), .B(T11553_Y));
KC_NOR2_X2 T11542 ( .Y(T11542_Y), .A(T4572_Q), .B(T11020_Y));
KC_NOR2_X2 T11541 ( .Y(T11541_Y), .A(T4576_Q), .B(T5947_Y));
KC_NOR2_X2 T11540 ( .Y(T11540_Y), .A(T15584_Y), .B(T4572_Q));
KC_NOR2_X2 T11539 ( .Y(T11539_Y), .A(T4556_Y), .B(T4547_Y));
KC_NOR2_X2 T11538 ( .Y(T11538_Y), .A(T4578_Q), .B(T4576_Q));
KC_NOR2_X2 T11537 ( .Y(T11537_Y), .A(T4578_Q), .B(T5954_Y));
KC_NOR2_X2 T11536 ( .Y(T11536_Y), .A(T5953_Y), .B(T4547_Y));
KC_NOR2_X2 T11535 ( .Y(T11535_Y), .A(T4546_Y), .B(T4556_Y));
KC_NOR2_X2 T11534 ( .Y(T11534_Y), .A(T11535_Y), .B(T5955_Y));
KC_NOR2_X2 T11533 ( .Y(T11533_Y), .A(T5953_Y), .B(T4546_Y));
KC_NOR2_X2 T11608 ( .Y(T11608_Y), .A(T4608_Q), .B(T4607_Q));
KC_NOR2_X2 T11607 ( .Y(T11607_Y), .A(T5159_Q), .B(T10957_Y));
KC_NOR2_X2 T11624 ( .Y(T11624_Y), .A(T4638_Y), .B(T16045_Y));
KC_NOR2_X2 T11707 ( .Y(T11707_Y), .A(T6169_Y), .B(T4694_Y));
KC_NOR2_X2 T11706 ( .Y(T11706_Y), .A(T4713_Q), .B(T4717_Q));
KC_NOR2_X2 T11705 ( .Y(T11705_Y), .A(T10601_Y), .B(T4739_Y));
KC_NOR2_X2 T10614 ( .Y(T10614_Y), .A(T16146_Y), .B(T10989_Y));
KC_NOR2_X2 T10613 ( .Y(T10613_Y), .A(T15757_Y), .B(T4711_Y));
KC_NOR2_X2 T10601 ( .Y(T10601_Y), .A(T4720_Q), .B(T4722_Q));
KC_NOR2_X2 T10600 ( .Y(T10600_Y), .A(T4719_Q), .B(T15757_Y));
KC_NOR2_X2 T10599 ( .Y(T10599_Y), .A(T4701_Y), .B(T4695_Y));
KC_NOR2_X2 T10598 ( .Y(T10598_Y), .A(T16146_Y), .B(T10981_Y));
KC_NOR2_X2 T10575 ( .Y(T10575_Y), .A(T6102_Y), .B(T6126_Y));
KC_NOR2_X2 T10574 ( .Y(T10574_Y), .A(T4720_Q), .B(T10575_Y));
KC_NOR2_X2 T11788 ( .Y(T11788_Y), .A(T4750_Q), .B(T4718_Q));
KC_NOR2_X2 T11787 ( .Y(T11787_Y), .A(T16145_Y), .B(T6244_Y));
KC_NOR2_X2 T11786 ( .Y(T11786_Y), .A(T16460_Q), .B(T11787_Y));
KC_NOR2_X2 T11779 ( .Y(T11779_Y), .A(T4758_Q), .B(T4731_Y));
KC_NOR2_X2 T11778 ( .Y(T11778_Y), .A(T4757_Q), .B(T4731_Y));
KC_NOR2_X2 T11777 ( .Y(T11777_Y), .A(T6234_Y), .B(T11786_Y));
KC_NOR2_X2 T10541 ( .Y(T10541_Y), .A(T4738_Y), .B(T10576_Y));
KC_NOR2_X2 T9394 ( .Y(T9394_Y), .A(T15195_Y), .B(T9393_Y));
KC_NOR2_X2 T9393 ( .Y(T9393_Y), .A(T15656_Y), .B(T7833_Y));
KC_NOR2_X2 T9392 ( .Y(T9392_Y), .A(T7582_Y), .B(T7696_Y));
KC_NOR2_X2 T9391 ( .Y(T9391_Y), .A(T7696_Y), .B(T7698_Y));
KC_NOR2_X2 T9356 ( .Y(T9356_Y), .A(T15841_Y), .B(T650_Y));
KC_NOR2_X2 T9485 ( .Y(T9485_Y), .A(T9174_Y), .B(T9125_Y));
KC_NOR2_X2 T9449 ( .Y(T9449_Y), .A(T9157_Y), .B(T9014_Y));
KC_NOR2_X2 T9448 ( .Y(T9448_Y), .A(T9126_Y), .B(T16287_Y));
KC_NOR2_X2 T9447 ( .Y(T9447_Y), .A(T16285_Y), .B(T9014_Y));
KC_NOR2_X2 T9382 ( .Y(T9382_Y), .A(T7676_Y), .B(T7582_Y));
KC_NOR2_X2 T9381 ( .Y(T9381_Y), .A(T382_Y), .B(T7816_Y));
KC_NOR2_X2 T9380 ( .Y(T9380_Y), .A(T16329_Y), .B(T9387_Y));
KC_NOR2_X2 T9379 ( .Y(T9379_Y), .A(T16329_Y), .B(T9375_Y));
KC_NOR2_X2 T9476 ( .Y(T9476_Y), .A(T4842_Y), .B(T9478_Y));
KC_NOR2_X2 T9475 ( .Y(T9475_Y), .A(T9166_Y), .B(T16185_Y));
KC_NOR2_X2 T9343 ( .Y(T9343_Y), .A(T6662_Y), .B(T5305_Q));
KC_NOR2_X2 T9258 ( .Y(T9258_Y), .A(T9513_Y), .B(T7067_Y));
KC_NOR2_X2 T9371 ( .Y(T9371_Y), .A(T7644_Y), .B(T900_Y));
KC_NOR2_X2 T9342 ( .Y(T9342_Y), .A(T8832_Y), .B(T7646_Y));
KC_NOR2_X2 T9341 ( .Y(T9341_Y), .A(T8832_Y), .B(T7645_Y));
KC_NOR2_X2 T9432 ( .Y(T9432_Y), .A(T10880_Y), .B(T9987_Y));
KC_NOR2_X2 T9365 ( .Y(T9365_Y), .A(T4872_Y), .B(T8938_Y));
KC_NOR2_X2 T9363 ( .Y(T9363_Y), .A(T8760_Y), .B(T9366_Y));
KC_NOR2_X2 T9362 ( .Y(T9362_Y), .A(T9369_Y), .B(T7868_Y));
KC_NOR2_X2 T9361 ( .Y(T9361_Y), .A(T8770_Y), .B(T8763_Y));
KC_NOR2_X2 T9360 ( .Y(T9360_Y), .A(T15654_Y), .B(T9369_Y));
KC_NOR2_X2 T9359 ( .Y(T9359_Y), .A(T9369_Y), .B(T7867_Y));
KC_NOR2_X2 T9300 ( .Y(T9300_Y), .A(T7592_Y), .B(T6699_Y));
KC_NOR2_X2 T9299 ( .Y(T9299_Y), .A(T8683_Y), .B(T7592_Y));
KC_NOR2_X2 T9298 ( .Y(T9298_Y), .A(T7592_Y), .B(T6625_Y));
KC_NOR2_X2 T10299 ( .Y(T10299_Y), .A(T11913_Y), .B(T13050_Y));
KC_NOR2_X2 T10298 ( .Y(T10298_Y), .A(T16274_Y), .B(T4872_Y));
KC_NOR2_X2 T9364 ( .Y(T9364_Y), .A(T15841_Y), .B(T9927_Y));
KC_NOR2_X2 T10327 ( .Y(T10327_Y), .A(T9896_Y), .B(T1085_Y));
KC_NOR2_X2 T10326 ( .Y(T10326_Y), .A(T9897_Y), .B(T1085_Y));
KC_NOR2_X2 T10296 ( .Y(T10296_Y), .A(T10880_Y), .B(T10143_Y));
KC_NOR2_X2 T10295 ( .Y(T10295_Y), .A(T10941_Y), .B(T10143_Y));
KC_NOR2_X2 T10294 ( .Y(T10294_Y), .A(T13121_Y), .B(T10143_Y));
KC_NOR2_X2 T10293 ( .Y(T10293_Y), .A(T4902_Y), .B(T1362_Y));
KC_NOR2_X2 T10368 ( .Y(T10368_Y), .A(T15677_Y), .B(T10426_Y));
KC_NOR2_X2 T10367 ( .Y(T10367_Y), .A(T7339_Y), .B(T10425_Y));
KC_NOR2_X2 T10366 ( .Y(T10366_Y), .A(T5674_Y), .B(T10428_Y));
KC_NOR2_X2 T10361 ( .Y(T10361_Y), .A(T6791_Y), .B(T10414_Y));
KC_NOR2_X2 T10360 ( .Y(T10360_Y), .A(T5663_Y), .B(T10414_Y));
KC_NOR2_X2 T10359 ( .Y(T10359_Y), .A(T6791_Y), .B(T10415_Y));
KC_NOR2_X2 T10358 ( .Y(T10358_Y), .A(T5663_Y), .B(T10415_Y));
KC_NOR2_X2 T10283 ( .Y(T10283_Y), .A(T15904_Y), .B(T16017_Y));
KC_NOR2_X2 T12052 ( .Y(T12052_Y), .A(T5494_Q), .B(T2259_Y));
KC_NOR2_X2 T12030 ( .Y(T12030_Y), .A(T16489_Y), .B(T5908_Y));
KC_NOR2_X2 T12022 ( .Y(T12022_Y), .A(T2854_Y), .B(T12350_Y));
KC_NOR2_X2 T10557 ( .Y(T10557_Y), .A(T12102_Y), .B(T15712_Y));
KC_NOR2_X2 T10526 ( .Y(T10526_Y), .A(T2054_Q), .B(T16366_Y));
KC_NOR2_X2 T10525 ( .Y(T10525_Y), .A(T2060_Y), .B(T9974_Y));
KC_NOR2_X2 T10478 ( .Y(T10478_Y), .A(T6768_Y), .B(T6778_Y));
KC_NOR2_X2 T10477 ( .Y(T10477_Y), .A(T6768_Y), .B(T6782_Y));
KC_NOR2_X2 T10442 ( .Y(T10442_Y), .A(T6768_Y), .B(T407_Y));
KC_NOR2_X2 T16261 ( .Y(T16261_Y), .A(T15533_Y), .B(T1544_Y));
KC_NOR2_X2 T10256 ( .Y(T10256_Y), .A(T10941_Y), .B(T2633_Y));
KC_NOR2_X2 T12049 ( .Y(T12049_Y), .A(T13320_Y), .B(T13321_Y));
KC_NOR2_X2 T12048 ( .Y(T12048_Y), .A(T6145_Y), .B(T5002_Y));
KC_NOR2_X2 T12029 ( .Y(T12029_Y), .A(T10949_Y), .B(T15882_Y));
KC_NOR2_X2 T12028 ( .Y(T12028_Y), .A(T16489_Y), .B(T11025_Y));
KC_NOR2_X2 T12009 ( .Y(T12009_Y), .A(T6067_Y), .B(T11640_Y));
KC_NOR2_X2 T12008 ( .Y(T12008_Y), .A(T12001_Y), .B(T11640_Y));
KC_NOR2_X2 T12007 ( .Y(T12007_Y), .A(T11640_Y), .B(T12006_Y));
KC_NOR2_X2 T11962 ( .Y(T11962_Y), .A(T10270_Y), .B(T12335_Y));
KC_NOR2_X2 T11961 ( .Y(T11961_Y), .A(T5421_Q), .B(T2661_Y));
KC_NOR2_X2 T11960 ( .Y(T11960_Y), .A(T2661_Y), .B(T10281_Y));
KC_NOR2_X2 T11038 ( .Y(T11038_Y), .A(T1_Y), .B(T6545_Y));
KC_NOR2_X2 T10551 ( .Y(T10551_Y), .A(T2893_Y), .B(T8281_Y));
KC_NOR2_X2 T10546 ( .Y(T10546_Y), .A(T15233_Y), .B(T2866_Y));
KC_NOR2_X2 T12045 ( .Y(T12045_Y), .A(T3362_Y), .B(T3429_Y));
KC_NOR2_X2 T12027 ( .Y(T12027_Y), .A(T2777_Y), .B(T15895_Y));
KC_NOR2_X2 T12001 ( .Y(T12001_Y), .A(T10584_Y), .B(T8345_Y));
KC_NOR2_X2 T12000 ( .Y(T12000_Y), .A(T6048_Y), .B(T5896_Y));
KC_NOR2_X2 T11991 ( .Y(T11991_Y), .A(T5428_Q), .B(T3201_Y));
KC_NOR2_X2 T11990 ( .Y(T11990_Y), .A(T5040_Y), .B(T3210_Y));
KC_NOR2_X2 T11989 ( .Y(T11989_Y), .A(T3210_Y), .B(T15562_Y));
KC_NOR2_X2 T10549 ( .Y(T10549_Y), .A(T6145_Y), .B(T2888_Y));
KC_NOR2_X2 T10548 ( .Y(T10548_Y), .A(T2848_Y), .B(T10544_Y));
KC_NOR2_X2 T10547 ( .Y(T10547_Y), .A(T15621_Y), .B(T6138_Y));
KC_NOR2_X2 T10544 ( .Y(T10544_Y), .A(T16138_Y), .B(T3447_Y));
KC_NOR2_X2 T10507 ( .Y(T10507_Y), .A(T5026_Y), .B(T859_Y));
KC_NOR2_X2 T10502 ( .Y(T10502_Y), .A(T3069_Y), .B(T9834_Y));
KC_NOR2_X2 T10501 ( .Y(T10501_Y), .A(T3069_Y), .B(T9831_Y));
KC_NOR2_X2 T10437 ( .Y(T10437_Y), .A(T3014_Y), .B(T9650_Y));
KC_NOR2_X2 T12039 ( .Y(T12039_Y), .A(T12038_Y), .B(T16106_Y));
KC_NOR2_X2 T12026 ( .Y(T12026_Y), .A(T3964_Q), .B(T15971_Y));
KC_NOR2_X2 T11985 ( .Y(T11985_Y), .A(T3856_Y), .B(T5803_Y));
KC_NOR2_X2 T11984 ( .Y(T11984_Y), .A(T5842_Y), .B(T3827_Y));
KC_NOR2_X2 T11969 ( .Y(T11969_Y), .A(T5838_Y), .B(T15907_Y));
KC_NOR2_X2 T11968 ( .Y(T11968_Y), .A(T3828_Y), .B(T3849_Y));
KC_NOR2_X2 T10542 ( .Y(T10542_Y), .A(T3368_Y), .B(T4093_Y));
KC_NOR2_X2 T10504 ( .Y(T10504_Y), .A(T16402_Y), .B(T9832_Y));
KC_NOR2_X2 T10503 ( .Y(T10503_Y), .A(T16402_Y), .B(T9831_Y));
KC_NOR2_X2 T12034 ( .Y(T12034_Y), .A(T8498_Y), .B(T4736_Y));
KC_NOR2_X2 T12033 ( .Y(T12033_Y), .A(T4696_Y), .B(T5146_Y));
KC_NOR2_X2 T12032 ( .Y(T12032_Y), .A(T10601_Y), .B(T4736_Y));
KC_NOR2_X2 T12031 ( .Y(T12031_Y), .A(T8498_Y), .B(T4739_Y));
KC_NOR2_X2 T12024 ( .Y(T12024_Y), .A(T15967_Y), .B(T5155_Y));
KC_NOR2_X2 T12023 ( .Y(T12023_Y), .A(T4528_Q), .B(T4519_Y));
KC_NOR2_X2 T12016 ( .Y(T12016_Y), .A(T4573_Q), .B(T4579_Q));
KC_NOR2_X2 T11977 ( .Y(T11977_Y), .A(T15869_Y), .B(T5778_Y));
KC_NOR2_X2 T10630 ( .Y(T10630_Y), .A(T13315_Y), .B(T8494_Y));
KC_NOR2_X2 T10431 ( .Y(T10431_Y), .A(T12785_Y), .B(T422_Y));
KC_NOR2_X2 T8544 ( .Y(T8544_Y), .A(T5619_Y), .B(T5617_Y));
KC_NOR2_X2 T9274 ( .Y(T9274_Y), .A(T822_Q), .B(T6290_Y));
KC_NOR2_X2 T8602 ( .Y(T8602_Y), .A(T5192_Q), .B(T6933_Y));
KC_NOR2_X2 T8586 ( .Y(T8586_Y), .A(T6353_Y), .B(T8588_Y));
KC_NOR2_X2 T6483 ( .Y(T6483_Y), .A(T3608_Y), .B(T10470_Y));
KC_NOR2_X2 T9672 ( .Y(T9672_Y), .A(T15682_Y), .B(T15400_Y));
KC_NOR2_X2 T9502 ( .Y(T9502_Y), .A(T9723_Y), .B(T7592_Y));
KC_NOR2_X2 T9766 ( .Y(T9766_Y), .A(T607_Y), .B(T9769_Y));
KC_NOR2_X2 T9728 ( .Y(T9728_Y), .A(T3621_Y), .B(T9770_Y));
KC_NOR2_X2 T9707 ( .Y(T9707_Y), .A(T6789_Y), .B(T10413_Y));
KC_NOR2_X2 T9705 ( .Y(T9705_Y), .A(T5650_Y), .B(T10413_Y));
KC_NOR2_X2 T9312 ( .Y(T9312_Y), .A(T7563_Y), .B(T7685_Y));
KC_NOR2_X2 T9786 ( .Y(T9786_Y), .A(T803_Y), .B(T9781_Y));
KC_NOR2_X2 T8825 ( .Y(T8825_Y), .A(T5344_Y), .B(T5344_Y));
KC_NOR2_X2 T8812 ( .Y(T8812_Y), .A(T15429_Y), .B(T9110_Y));
KC_NOR2_X2 T8793 ( .Y(T8793_Y), .A(T15841_Y), .B(T11244_Y));
KC_NOR2_X2 T10079 ( .Y(T10079_Y), .A(T12091_Y), .B(T5325_Y));
KC_NOR2_X2 T9028 ( .Y(T9028_Y), .A(T16289_Y), .B(T1430_Y));
KC_NOR2_X2 T8900 ( .Y(T8900_Y), .A(T9416_Y), .B(T1199_Y));
KC_NOR2_X2 T9137 ( .Y(T9137_Y), .A(T15091_Y), .B(T15092_Y));
KC_NOR2_X2 T9104 ( .Y(T9104_Y), .A(T9129_Y), .B(T15524_Y));
KC_NOR2_X2 T9064 ( .Y(T9064_Y), .A(T9077_Y), .B(T15524_Y));
KC_NOR2_X2 T11438 ( .Y(T11438_Y), .A(T5058_Y), .B(T2140_Y));
KC_NOR2_X2 T11516 ( .Y(T11516_Y), .A(T2777_Y), .B(T15853_Y));
KC_NOR2_X2 T12013 ( .Y(T12013_Y), .A(T4558_Y), .B(T8477_Y));
KC_NOR2_X2 T11571 ( .Y(T11571_Y), .A(T11535_Y), .B(T12015_Y));
KC_NOR2_X2 T11546 ( .Y(T11546_Y), .A(T3331_Y), .B(T5570_Y));
KC_NOR2_X2 T12042 ( .Y(T12042_Y), .A(T12876_Y), .B(T10966_Y));
KC_NOR2_X2 T11996 ( .Y(T11996_Y), .A(T4176_Q), .B(T4179_Q));
KC_NOR2_X2 T11657 ( .Y(T11657_Y), .A(T11643_Y), .B(T11637_Y));
KC_NOR2_X2 T11652 ( .Y(T11652_Y), .A(T5486_Q), .B(T4912_Y));
KC_NOR2_X2 T11637 ( .Y(T11637_Y), .A(T4031_Y), .B(T3400_Y));
KC_NOR2_X2 T11627 ( .Y(T11627_Y), .A(T4176_Q), .B(T3374_Y));
KC_NOR2_X2 T10583 ( .Y(T10583_Y), .A(T4070_Y), .B(T3389_Y));
KC_NOR2_X2 T11772 ( .Y(T11772_Y), .A(T6565_Y), .B(T3483_Y));
KC_NOR2_X2 T11766 ( .Y(T11766_Y), .A(T12064_Y), .B(T3486_Y));
KC_NOR2_X2 T10627 ( .Y(T10627_Y), .A(T2313_Q), .B(T2310_Y));
KC_NOR2_X2 T11831 ( .Y(T11831_Y), .A(T3506_Y), .B(T11004_Y));
KC_NOR2_X2 T11825 ( .Y(T11825_Y), .A(T6520_Y), .B(T11828_Y));
KC_NOR2_X2 T11815 ( .Y(T11815_Y), .A(T6530_Y), .B(T11000_Y));
KC_NOR2_X2 T11976 ( .Y(T11976_Y), .A(T11402_Y), .B(T11981_Y));
KC_NOR2_X2 T11970 ( .Y(T11970_Y), .A(T15881_Y), .B(T15943_Y));
KC_NOR2_X2 T10474 ( .Y(T10474_Y), .A(T6768_Y), .B(T15686_Y));
KC_NOR2_X2 T10472 ( .Y(T10472_Y), .A(T15682_Y), .B(T411_Y));
KC_NOR2_X2 T10300 ( .Y(T10300_Y), .A(T10942_Y), .B(T10143_Y));
KC_NOR2_X2 T9452 ( .Y(T9452_Y), .A(T9093_Y), .B(T16287_Y));
KC_AOI31_X2 T8536 ( .B2(T8559_Y), .B0(T5203_Q), .Y(T8536_Y),     .A(T15317_Y), .B1(T8543_Y));
KC_AOI31_X2 T8552 ( .B2(T15314_Y), .B0(T120_Y), .Y(T8552_Y),     .A(T12470_Y), .B1(T5600_Y));
KC_AOI31_X2 T8551 ( .B2(T126_Y), .B0(T120_Y), .Y(T8551_Y),     .A(T12470_Y), .B1(T15312_Y));
KC_AOI31_X2 T8597 ( .B2(T8591_Y), .B0(T133_Q), .Y(T8597_Y),     .A(T8608_Y), .B1(T5222_Q));
KC_AOI31_X2 T8596 ( .B2(T15358_Y), .B0(T150_Q), .Y(T8596_Y),     .A(T8602_Y), .B1(T8601_Y));
KC_AOI31_X2 T8595 ( .B2(T6944_Y), .B0(T8599_Y), .Y(T8595_Y),     .A(T12475_Y), .B1(T350_Y));
KC_AOI31_X2 T8590 ( .B2(T236_Y), .B0(T255_Y), .Y(T8590_Y), .A(T6945_Y),     .B1(T8577_Y));
KC_AOI31_X2 T8567 ( .B2(T9286_Y), .B0(T6968_Y), .Y(T8567_Y),     .A(T12475_Y), .B1(T15353_Y));
KC_AOI31_X2 T8755 ( .B2(T230_Y), .B0(T8705_Y), .Y(T8755_Y),     .A(T12608_Y), .B1(T9391_Y));
KC_AOI31_X2 T8706 ( .B2(T16176_Y), .B0(T9391_Y), .Y(T8706_Y),     .A(T12608_Y), .B1(T205_Y));
KC_AOI31_X2 T8705 ( .B2(T743_Y), .B0(T212_Q), .Y(T8705_Y), .A(T7681_Y),     .B1(T15765_Y));
KC_AOI31_X2 T8778 ( .B2(T8108_Y), .B0(T8777_Y), .Y(T8778_Y),     .A(T11227_Y), .B1(T9381_Y));
KC_AOI31_X2 T8910 ( .B2(T9018_Y), .B0(T8865_Y), .Y(T8910_Y),     .A(T11271_Y), .B1(T8950_Y));
KC_AOI31_X2 T9114 ( .B2(T2392_Y), .B0(T15091_Y), .Y(T9114_Y),     .A(T4820_Y), .B1(T9117_Y));
KC_AOI31_X2 T8751 ( .B2(T550_Q), .B0(T541_Q), .Y(T8751_Y), .A(T8894_Y),     .B1(T544_Q));
KC_AOI31_X2 T1256 ( .B2(T7901_Y), .B0(T8900_Y), .Y(T1256_Y),     .A(T12720_Y), .B1(T8042_Y));
KC_AOI31_X2 T8941 ( .B2(T1328_Y), .B0(T566_Q), .Y(T8941_Y),     .A(T8071_Y), .B1(T8118_Y));
KC_AOI31_X2 T8906 ( .B2(T8908_Y), .B0(T16385_Y), .Y(T8906_Y),     .A(T12720_Y), .B1(T16408_Y));
KC_AOI31_X2 T8897 ( .B2(T8046_Y), .B0(T16408_Y), .Y(T8897_Y),     .A(T12720_Y), .B1(T8035_Y));
KC_AOI31_X2 T8896 ( .B2(T8035_Y), .B0(T8940_Y), .Y(T8896_Y),     .A(T12720_Y), .B1(T8900_Y));
KC_AOI31_X2 T8736 ( .B2(T12438_Y), .B0(T12611_Y), .Y(T8736_Y),     .A(T16387_Y), .B1(T7244_Y));
KC_AOI31_X2 T8940 ( .B2(T12456_Y), .B0(T9096_Y), .Y(T8940_Y),     .A(T12721_Y), .B1(T1198_Y));
KC_AOI31_X2 T8655 ( .B2(T1039_Y), .B0(T498_Y), .Y(T8655_Y),     .A(T8728_Y), .B1(T712_Q));
KC_AOI31_X2 T8724 ( .B2(T5360_Q), .B0(T638_Y), .Y(T8724_Y), .A(T719_Y),     .B1(T7558_Y));
KC_AOI31_X2 T945 ( .B2(T7840_Y), .B0(T8890_Y), .Y(T945_Y),     .A(T12884_Y), .B1(T7846_Y));
KC_AOI31_X2 T8844 ( .B2(T8849_Y), .B0(T8890_Y), .Y(T8844_Y),     .A(T12884_Y), .B1(T5347_Y));
KC_AOI31_X2 T8973 ( .B2(T1342_Y), .B0(T1197_Y), .Y(T8973_Y),     .A(T1341_Y), .B1(T15487_Y));
KC_AOI31_X2 T8789 ( .B2(T16117_Y), .B0(T8850_Y), .Y(T8789_Y),     .A(T15841_Y), .B1(T15455_Y));
KC_AOI31_X2 T8933 ( .B2(T1342_Y), .B0(T8974_Y), .Y(T8933_Y),     .A(T1341_Y), .B1(T1197_Y));
KC_AOI31_X2 T8932 ( .B2(T15486_Y), .B0(T1197_Y), .Y(T8932_Y),     .A(T1341_Y), .B1(T1458_Y));
KC_AOI31_X2 T10152 ( .B2(T86_Y), .B0(T15529_Y), .Y(T10152_Y),     .A(T16005_Y), .B1(T1362_Y));
KC_AOI31_X2 T10520 ( .B2(T1142_Y), .B0(T2023_Q), .Y(T10520_Y),     .A(T5363_Q), .B1(T9969_Y));
KC_AOI31_X2 T10099 ( .B2(T1548_Y), .B0(T10079_Y), .Y(T10099_Y),     .A(T12065_Y), .B1(T15814_Y));
KC_AOI31_X2 T8219 ( .B2(T11450_Y), .B0(T2162_Q), .Y(T8219_Y),     .A(T4010_Y), .B1(T2160_Q));
KC_AOI31_X2 T8242 ( .B2(T2172_Y), .B0(T2184_Y), .Y(T8242_Y),     .A(T2183_Y), .B1(T15959_Y));
KC_AOI31_X2 T8485 ( .B2(T2781_Y), .B0(T6280_Y), .Y(T8485_Y),     .A(T2854_Y), .B1(T12230_Y));
KC_AOI31_X2 T8298 ( .B2(T2194_Y), .B0(T6302_Y), .Y(T8298_Y),     .A(T2854_Y), .B1(T2174_Y));
KC_AOI31_X2 T8287 ( .B2(T2774_Y), .B0(T15983_Y), .Y(T8287_Y),     .A(T2854_Y), .B1(T12234_Y));
KC_AOI31_X2 T8283 ( .B2(T2772_Y), .B0(T6273_Y), .Y(T8283_Y),     .A(T2854_Y), .B1(T12218_Y));
KC_AOI31_X2 T9778 ( .B2(T634_Y), .B0(T15419_Y), .Y(T9778_Y),     .A(T6849_Y), .B1(T9744_Y));
KC_AOI31_X2 T9873 ( .B2(T15447_Y), .B0(T15447_Y), .Y(T9873_Y),     .A(T12085_Y), .B1(T15447_Y));
KC_AOI31_X2 T10056 ( .B2(T12091_Y), .B0(T10060_Y), .Y(T10056_Y),     .A(T15502_Y), .B1(T1509_Y));
KC_AOI31_X2 T10248 ( .B2(T5750_Y), .B0(T6729_Y), .Y(T10248_Y),     .A(T11355_Y), .B1(T10250_Y));
KC_AOI31_X2 T8228 ( .B2(T8496_Y), .B0(T12189_Y), .Y(T8228_Y),     .A(T3408_Y), .B1(T2727_Y));
KC_AOI31_X2 T8261 ( .B2(T5925_Y), .B0(T5465_Q), .Y(T8261_Y),     .A(T6011_Y), .B1(T5461_Q));
KC_AOI31_X2 T8250 ( .B2(T11597_Y), .B0(T11464_Y), .Y(T8250_Y),     .A(T5465_Q), .B1(T11449_Y));
KC_AOI31_X2 T8241 ( .B2(T15606_Y), .B0(T16156_Y), .Y(T8241_Y),     .A(T12203_Y), .B1(T2879_Y));
KC_AOI31_X2 T16025 ( .B2(T8261_Y), .B0(T15600_Y), .Y(T16025_Y),     .A(T6055_Y), .B1(T11996_Y));
KC_AOI31_X2 T8316 ( .B2(T3411_Y), .B0(T11603_Y), .Y(T8316_Y),     .A(T15942_Y), .B1(T6082_Y));
KC_AOI31_X2 T8306 ( .B2(T16038_Y), .B0(T15600_Y), .Y(T8306_Y),     .A(T6026_Y), .B1(T8261_Y));
KC_AOI31_X2 T8362 ( .B2(T3379_Y), .B0(T5539_Y), .Y(T8362_Y),     .A(T6066_Y), .B1(T11029_Y));
KC_AOI31_X2 T8346 ( .B2(T12005_Y), .B0(T15802_Q), .Y(T8346_Y),     .A(T2832_Q), .B1(T3396_Y));
KC_AOI31_X2 T6577 ( .B2(T2908_Y), .B0(T12311_Y), .Y(T6577_Y),     .A(T6578_Y), .B1(T2901_Y));
KC_AOI31_X2 T8515 ( .B2(T10559_Y), .B0(T2886_Y), .Y(T8515_Y),     .A(T2882_Y), .B1(T10561_Y));
KC_AOI31_X2 T8417 ( .B2(T6222_Y), .B0(T6223_Y), .Y(T8417_Y),     .A(T11768_Y), .B1(T11810_Y));
KC_AOI31_X2 T8416 ( .B2(T2894_Y), .B0(T11808_Y), .Y(T8416_Y),     .A(T2911_Y), .B1(T2318_Y));
KC_AOI31_X2 T8409 ( .B2(T2898_Y), .B0(T12106_Y), .Y(T8409_Y),     .A(T6080_Y), .B1(T12103_Y));
KC_AOI31_X2 T9752 ( .B2(T3062_Y), .B0(T3061_Y), .Y(T9752_Y),     .A(T15420_Y), .B1(T2494_Y));
KC_AOI31_X2 T8187 ( .B2(T3207_Y), .B0(T12130_Y), .Y(T8187_Y),     .A(T5774_Y), .B1(T3815_Y));
KC_AOI31_X2 T8257 ( .B2(T3300_Y), .B0(T5922_Y), .Y(T8257_Y),     .A(T12206_Y), .B1(T3300_Y));
KC_AOI31_X2 T8239 ( .B2(T5065_Y), .B0(T3307_Y), .Y(T8239_Y),     .A(T3299_Y), .B1(T5065_Y));
KC_AOI31_X2 T8324 ( .B2(T16015_Y), .B0(T3360_Y), .Y(T8324_Y),     .A(T15607_Y), .B1(T7915_Y));
KC_AOI31_X2 T8307 ( .B2(T5996_Y), .B0(T16102_Y), .Y(T8307_Y),     .A(T13148_Y), .B1(T16037_Y));
KC_AOI31_X2 T8469 ( .B2(T5059_Y), .B0(T6069_Y), .Y(T8469_Y),     .A(T6006_Y), .B1(T6051_Y));
KC_AOI31_X2 T8345 ( .B2(T16044_Y), .B0(T3375_Y), .Y(T8345_Y),     .A(T3395_Y), .B1(T10966_Y));
KC_AOI31_X2 T8377 ( .B2(T16167_Y), .B0(T15616_Y), .Y(T8377_Y),     .A(T11816_Y), .B1(T15234_Y));
KC_AOI31_X2 T8415 ( .B2(T3474_Y), .B0(T3471_Y), .Y(T8415_Y),     .A(T2865_Y), .B1(T3479_Y));
KC_AOI31_X2 T8170 ( .B2(T11822_Y), .B0(T6049_Y), .Y(T8170_Y),     .A(T3512_Y), .B1(T11746_Y));
KC_AOI31_X2 T8167 ( .B2(T8170_Y), .B0(T3523_Q), .Y(T8167_Y),     .A(T12875_Y), .B1(T11042_Y));
KC_AOI31_X2 T9861 ( .B2(T3657_Y), .B0(T3707_Y), .Y(T9861_Y),     .A(T3681_Y), .B1(T857_Y));
KC_AOI31_X2 T5779 ( .B2(T14942_Q), .B0(T11353_Y), .Y(T5779_Y),     .A(T11315_Y), .B1(T5826_Y));
KC_AOI31_X2 T8452 ( .B2(T5789_Y), .B0(T11969_Y), .Y(T8452_Y),     .A(T6746_Y), .B1(T14942_Q));
KC_AOI31_X2 T8451 ( .B2(T11982_Y), .B0(T14942_Q), .Y(T8451_Y),     .A(T11372_Y), .B1(T11393_Y));
KC_AOI31_X2 T8186 ( .B2(T11985_Y), .B0(T5830_Y), .Y(T8186_Y),     .A(T12956_Y), .B1(T11365_Y));
KC_AOI31_X2 T8185 ( .B2(T5838_Y), .B0(T11365_Y), .Y(T8185_Y),     .A(T8176_Y), .B1(T11985_Y));
KC_AOI31_X2 T8176 ( .B2(T3816_Y), .B0(T5781_Y), .Y(T8176_Y),     .A(T5780_Y), .B1(T5756_Y));
KC_AOI31_X2 T8204 ( .B2(T12167_Y), .B0(T11379_Y), .Y(T8204_Y),     .A(T6116_Y), .B1(T11402_Y));
KC_AOI31_X2 T8201 ( .B2(T15888_Y), .B0(T11367_Y), .Y(T8201_Y),     .A(T11407_Y), .B1(T3854_Y));
KC_AOI31_X2 T8196 ( .B2(T5822_Y), .B0(T15877_Y), .Y(T8196_Y),     .A(T11388_Y), .B1(T11378_Y));
KC_AOI31_X2 T8193 ( .B2(T5802_Y), .B0(T145_Q), .Y(T8193_Y),     .A(T13306_Y), .B1(T11428_Y));
KC_AOI31_X2 T8192 ( .B2(T4460_Y), .B0(T3848_Y), .Y(T8192_Y),     .A(T5803_Y), .B1(T10915_Y));
KC_AOI31_X2 T8190 ( .B2(T5837_Y), .B0(T145_Q), .Y(T8190_Y),     .A(T15901_Y), .B1(T4487_Q));
KC_AOI31_X2 T15933 ( .B2(T15903_Y), .B0(T2073_Y), .Y(T15933_Y),     .A(T5454_Y), .B1(T5457_Y));
KC_AOI31_X2 T8445 ( .B2(T3856_Y), .B0(T11969_Y), .Y(T8445_Y),     .A(T11968_Y), .B1(T5788_Y));
KC_AOI31_X2 T8444 ( .B2(T5788_Y), .B0(T11969_Y), .Y(T8444_Y),     .A(T11968_Y), .B1(T11367_Y));
KC_AOI31_X2 T5936 ( .B2(T10940_Y), .B0(T8264_Y), .Y(T5936_Y),     .A(T10940_Y), .B1(T10940_Y));
KC_AOI31_X2 T8272 ( .B2(T11616_Y), .B0(T3974_Q), .Y(T8272_Y),     .A(T5958_Y), .B1(T5981_Y));
KC_AOI31_X2 T8271 ( .B2(T6251_Y), .B0(T5905_Y), .Y(T8271_Y),     .A(T3975_Y), .B1(T8290_Y));
KC_AOI31_X2 T8373 ( .B2(T6048_Y), .B0(T6526_Q), .Y(T8373_Y),     .A(T4022_Y), .B1(T6062_Y));
KC_AOI31_X2 T8381 ( .B2(T4078_Y), .B0(T6111_Y), .Y(T8381_Y),     .A(T4083_Y), .B1(T4073_Y));
KC_AOI31_X2 T8376 ( .B2(T4088_Y), .B0(T10582_Y), .Y(T8376_Y),     .A(T6119_Y), .B1(T10578_Y));
KC_AOI31_X2 T8203 ( .B2(T5440_Y), .B0(T6113_Y), .Y(T8203_Y),     .A(T11423_Y), .B1(T11366_Y));
KC_AOI31_X2 T8200 ( .B2(T4441_Y), .B0(T5824_Y), .Y(T8200_Y),     .A(T8201_Y), .B1(T4446_Y));
KC_AOI31_X2 T8195 ( .B2(T3839_Y), .B0(T5816_Y), .Y(T8195_Y),     .A(T15908_Y), .B1(T10910_Y));
KC_AOI31_X2 T8194 ( .B2(T13090_Y), .B0(T11393_Y), .Y(T8194_Y),     .A(T11389_Y), .B1(T145_Q));
KC_AOI31_X2 T15937 ( .B2(T15936_Y), .B0(T10632_Y), .Y(T15937_Y),     .A(T2757_Y), .B1(T6217_Y));
KC_AOI31_X2 T8220 ( .B2(T1276_Y), .B0(T12183_Y), .Y(T8220_Y),     .A(T2757_Y), .B1(T147_Y));
KC_AOI31_X2 T8263 ( .B2(T12816_Y), .B0(T12207_Y), .Y(T8263_Y),     .A(T2757_Y), .B1(T1276_Y));
KC_AOI31_X2 T8254 ( .B2(T4525_Y), .B0(T5140_Y), .Y(T8254_Y),     .A(T12208_Y), .B1(T5917_Y));
KC_AOI31_X2 T8243 ( .B2(T4508_Y), .B0(T146_Y), .Y(T8243_Y),     .A(T2757_Y), .B1(T10937_Y));
KC_AOI31_X2 T8235 ( .B2(T4521_Y), .B0(T4568_Q), .Y(T8235_Y),     .A(T11506_Y), .B1(T4474_Y));
KC_AOI31_X2 T8474 ( .B2(T6241_Y), .B0(T8272_Y), .Y(T8474_Y),     .A(T2757_Y), .B1(T4584_Y));
KC_AOI31_X2 T8291 ( .B2(T3960_Y), .B0(T11570_Y), .Y(T8291_Y),     .A(T2757_Y), .B1(T12223_Y));
KC_AOI31_X2 T8288 ( .B2(T4559_Y), .B0(T12221_Y), .Y(T8288_Y),     .A(T2757_Y), .B1(T149_Y));
KC_AOI31_X2 T8284 ( .B2(T15586_Y), .B0(T11554_Y), .Y(T8284_Y),     .A(T2757_Y), .B1(T4551_Y));
KC_AOI31_X2 T8312 ( .B2(T3973_Y), .B0(T3982_Y), .Y(T8312_Y),     .A(T6326_Y), .B1(T12237_Y));
KC_AOI31_X2 T9455 ( .B2(T9080_S), .B0(T9080_Co), .Y(T9455_Y),     .A(T9024_Y), .B1(T4808_Y));
KC_AOI31_X2 T9262 ( .B2(T9283_Y), .B0(T6245_Y), .Y(T9262_Y),     .A(T8640_Y), .B1(T9278_Y));
KC_AOI31_X2 T8448 ( .B2(T2133_Y), .B0(T5444_Y), .Y(T8448_Y),     .A(T13303_Y), .B1(T6737_Y));
KC_AOI31_X2 T8508 ( .B2(T3447_Y), .B0(T11818_Y), .Y(T8508_Y),     .A(T13164_Y), .B1(T8361_Y));
KC_AOI31_X2 T8487 ( .B2(T3297_Y), .B0(T8488_Y), .Y(T8487_Y),     .A(T8486_Y), .B1(T3297_Y));
KC_AOI31_X2 T8466 ( .B2(T11018_Y), .B0(T3356_Y), .Y(T8466_Y),     .A(T6176_Y), .B1(T16043_Y));
KC_AOI31_X2 T8478 ( .B2(T10937_Y), .B0(T11577_Y), .Y(T8478_Y),     .A(T3981_Y), .B1(T11616_Y));
KC_AOI31_X2 T8166 ( .B2(T4175_Y), .B0(T4180_Y), .Y(T8166_Y),     .A(T8163_Y), .B1(T4761_Y));
KC_AOI31_X2 T8494 ( .B2(T15577_Y), .B0(T4531_Y), .Y(T8494_Y),     .A(T6194_S), .B1(T4529_Y));
KC_AOI31_X2 T10471 ( .B2(T2496_Y), .B0(T1535_Y), .Y(T10471_Y),     .A(T5270_Y), .B1(T15681_Y));
KC_AOI31_X2 T8888 ( .B2(T15487_Y), .B0(T8891_Y), .Y(T8888_Y),     .A(T12884_Y), .B1(T1458_Y));
KC_AOI31_X2 T8887 ( .B2(T937_Y), .B0(T128_Y), .Y(T8887_Y),     .A(T12884_Y), .B1(T16421_Y));
KC_AOI31_X2 T9132 ( .B2(T16158_Y), .B0(T15093_Y), .Y(T9132_Y),     .A(T9099_Y), .B1(T15109_Y));
KC_AOI31_X2 T8468 ( .B2(T11019_Y), .B0(T3377_Y), .Y(T8468_Y),     .A(T11675_Y), .B1(T2805_Y));
KC_AOI31_X2 T8349 ( .B2(T16099_Y), .B0(T11675_Y), .Y(T8349_Y),     .A(T11769_Y), .B1(T6050_Y));
KC_AOI31_X2 T8172 ( .B2(T11834_Y), .B0(T12102_Y), .Y(T8172_Y),     .A(T12875_Y), .B1(T11747_Y));
KC_AOI31_X2 T8154 ( .B2(T6491_Y), .B0(T2947_Y), .Y(T8154_Y),     .A(T8160_Y), .B1(T11844_Y));
KC_AOI31_X2 T8493 ( .B2(T11025_Y), .B0(T6007_Y), .Y(T8493_Y),     .A(T3411_Y), .B1(T2848_Y));
KC_AO2222_X1 T8638 ( .Y(T8638_Y), .A0(T12412_Y), .A1(T293_Q),     .B0(T12413_Y), .B1(T5226_Q), .C0(T12411_Y), .C1(T5241_Q),     .D0(T12440_Y), .D1(T288_Q));
KC_AO2222_X1 T8625 ( .Y(T8625_Y), .A0(T12412_Y), .A1(T313_Q),     .B0(T12413_Y), .B1(T158_Q), .C0(T12411_Y), .C1(T306_Q),     .D0(T12440_Y), .D1(T4822_Q));
KC_AO2222_X1 T8646 ( .Y(T8646_Y), .A0(T12412_Y), .A1(T5263_Q),     .B0(T12413_Y), .B1(T174_Q), .C0(T12411_Y), .C1(T326_Q),     .D0(T12440_Y), .D1(T5255_Q));
KC_AO2222_X1 T8669 ( .Y(T8669_Y), .A0(T12412_Y), .A1(T335_Q),     .B0(T12413_Y), .B1(T182_Q), .C0(T12411_Y), .C1(T344_Q),     .D0(T12440_Y), .D1(T5275_Q));
KC_AO2222_X1 T8666 ( .Y(T8666_Y), .A0(T12412_Y), .A1(T9350_Q),     .B0(T5281_Q), .B1(T12413_Y), .C0(T524_Q), .C1(T12411_Y),     .D0(T12440_Y), .D1(T337_Q));
KC_AO2222_X1 T8665 ( .Y(T8665_Y), .A0(T12412_Y), .A1(T9349_Q),     .B0(T12413_Y), .B1(T9352_Q), .C0(T12411_Y), .C1(T362_Q),     .D0(T12440_Y), .D1(T5277_Q));
KC_AO2222_X1 T7950 ( .Y(T7950_Y), .A0(T11893_Y), .A1(T8697_Y),     .B0(T8704_Y), .B1(T8741_Y), .C0(T9143_Y), .C1(T8742_Y),     .D0(T8740_Y), .D1(T8720_Y));
KC_AO2222_X1 T8723 ( .Y(T8723_Y), .A0(T11188_Y), .A1(T8697_Y),     .B0(T11214_Y), .B1(T8741_Y), .C0(T8742_Y), .C1(T9149_Y),     .D0(T8607_Y), .D1(T8740_Y));
KC_AO2222_X1 T8837 ( .Y(T8837_Y), .A0(T15451_Y), .A1(T8868_Y),     .B0(T8917_Y), .B1(T8812_Y), .C0(T9148_Y), .C1(T8867_Y),     .D0(T8638_Y), .D1(T8811_Y));
KC_AO2222_X1 T8836 ( .Y(T8836_Y), .A0(T11266_Y), .A1(T8812_Y),     .B0(T8951_Y), .B1(T8868_Y), .C0(T9017_Y), .C1(T8867_Y),     .D0(T8811_Y), .D1(T8711_Y));
KC_AO2222_X1 T8814 ( .Y(T8814_Y), .A0(T11270_Y), .A1(T8812_Y),     .B0(T11246_Y), .B1(T8868_Y), .C0(T8648_Y), .C1(T8811_Y),     .D0(T9101_Y), .D1(T8867_Y));
KC_AO2222_X1 T8813 ( .Y(T8813_Y), .A0(T11247_Y), .A1(T8812_Y),     .B0(T11270_Y), .B1(T8868_Y), .C0(T8867_Y), .C1(T9066_Y),     .D0(T8605_Y), .D1(T8811_Y));
KC_AO2222_X1 T8637 ( .Y(T8637_Y), .A0(T12412_Y), .A1(T459_Q),     .B0(T12440_Y), .B1(T5221_Q), .C0(T12413_Y), .C1(T5193_Q),     .D0(T12411_Y), .D1(T296_Q));
KC_AO2222_X1 T9511 ( .Y(T9511_Y), .A0(T12412_Y), .A1(T5254_Q),     .B0(T12440_Y), .B1(T489_Q), .C0(T12413_Y), .C1(T5261_Q),     .D0(T12411_Y), .D1(T329_Q));
KC_AO2222_X1 T8654 ( .Y(T8654_Y), .A0(T12412_Y), .A1(T5265_Q),     .B0(T12440_Y), .B1(T460_Q), .C0(T12413_Y), .C1(T4835_Q),     .D0(T12411_Y), .D1(T275_Q));
KC_AO2222_X1 T8651 ( .Y(T8651_Y), .A0(T12412_Y), .A1(T5257_Q),     .B0(T12440_Y), .B1(T5260_Q), .C0(T12413_Y), .C1(T672_Q),     .D0(T12411_Y), .D1(T323_Q));
KC_AO2222_X1 T8679 ( .Y(T8679_Y), .A0(T12412_Y), .A1(T519_Q),     .B0(T12440_Y), .B1(T501_Q), .C0(T12413_Y), .C1(T5282_Q),     .D0(T12411_Y), .D1(T5304_Q));
KC_AO2222_X1 T8663 ( .Y(T8663_Y), .A0(T12412_Y), .A1(T525_Q),     .B0(T12440_Y), .B1(T500_Q), .C0(T12413_Y), .C1(T5279_Q),     .D0(T12411_Y), .D1(T343_Q));
KC_AO2222_X1 T8738 ( .Y(T8738_Y), .A0(T12412_Y), .A1(T543_Q),     .B0(T12413_Y), .B1(T517_Q), .C0(T5346_Q), .C1(T12440_Y),     .D0(T12411_Y), .D1(T4840_Q));
KC_AO2222_X1 T8695 ( .Y(T8695_Y), .A0(T12412_Y), .A1(T5356_Q),     .B0(T12413_Y), .B1(T4827_Q), .C0(T551_Q), .C1(T12440_Y),     .D0(T529_Q), .D1(T12411_Y));
KC_AO2222_X1 T8694 ( .Y(T8694_Y), .A0(T12412_Y), .A1(T544_Q),     .B0(T12413_Y), .B1(T528_Q), .C0(T541_Q), .C1(T12440_Y),     .D0(T550_Q), .D1(T12411_Y));
KC_AO2222_X1 T8692 ( .Y(T8692_Y), .A0(T12416_Y), .A1(T5357_Q),     .B0(T12417_Y), .B1(T512_Q), .C0(T12414_Y), .C1(T5350_Q),     .D0(T12415_Y), .D1(T530_Q));
KC_AO2222_X1 T8691 ( .Y(T8691_Y), .A0(T12416_Y), .A1(T722_Q),     .B0(T12417_Y), .B1(T714_Q), .C0(T12414_Y), .C1(T5342_Q),     .D0(T12415_Y), .D1(T741_Q));
KC_AO2222_X1 T8861 ( .Y(T8861_Y), .A0(T571_Y), .A1(T8868_Y),     .B0(T8631_Y), .B1(T8811_Y), .C0(T969_Y), .C1(T8812_Y),     .D0(T8867_Y), .D1(T9488_Y));
KC_AO2222_X1 T8807 ( .Y(T8807_Y), .A0(T571_Y), .A1(T8812_Y),     .B0(T8907_Y), .B1(T8868_Y), .C0(T240_Y), .C1(T8867_Y),     .D0(T9320_Y), .D1(T8811_Y));
KC_AO2222_X1 T8635 ( .Y(T8635_Y), .A0(T12416_Y), .A1(T449_Q),     .B0(T12417_Y), .B1(T436_Q), .C0(T12415_Y), .C1(T657_Q),     .D0(T12414_Y), .D1(T453_Q));
KC_AO2222_X1 T8632 ( .Y(T8632_Y), .A0(T12416_Y), .A1(T838_Q),     .B0(T12414_Y), .B1(T848_Q), .C0(T12417_Y), .C1(T826_Q),     .D0(T12415_Y), .D1(T820_Q));
KC_AO2222_X1 T8631 ( .Y(T8631_Y), .A0(T12416_Y), .A1(T817_Q),     .B0(T12417_Y), .B1(T5229_Q), .C0(T12415_Y), .C1(T843_Q),     .D0(T12414_Y), .D1(T812_Q));
KC_AO2222_X1 T8610 ( .Y(T8610_Y), .A0(T12416_Y), .A1(T823_Q),     .B0(T12417_Y), .B1(T815_Q), .C0(T12415_Y), .C1(T834_Q),     .D0(T12414_Y), .D1(T824_Q));
KC_AO2222_X1 T8607 ( .Y(T8607_Y), .A0(T12416_Y), .A1(T4845_Q),     .B0(T12414_Y), .B1(T445_Q), .C0(T12417_Y), .C1(T5194_Q),     .D0(T12415_Y), .D1(T5223_Q));
KC_AO2222_X1 T8606 ( .Y(T8606_Y), .A0(T12416_Y), .A1(T4846_Q),     .B0(T12414_Y), .B1(T452_Q), .C0(T12417_Y), .C1(T432_Q),     .D0(T12415_Y), .D1(T456_Q));
KC_AO2222_X1 T8649 ( .Y(T8649_Y), .A0(T12416_Y), .A1(T828_Q),     .B0(T12414_Y), .B1(T4854_Q), .C0(T12417_Y), .C1(T5238_Q),     .D0(T12415_Y), .D1(T5259_Q));
KC_AO2222_X1 T8648 ( .Y(T8648_Y), .A0(T12416_Y), .A1(T861_Q),     .B0(T12417_Y), .B1(T860_Q), .C0(T12415_Y), .C1(T5258_Q),     .D0(T12414_Y), .D1(T5565_Q));
KC_AO2222_X1 T9310 ( .Y(T9310_Y), .A0(T12416_Y), .A1(T696_Q),     .B0(T12417_Y), .B1(T6487_Q), .C0(T12414_Y), .C1(T6486_Q),     .D0(T12415_Y), .D1(T865_Q));
KC_AO2222_X1 T8720 ( .Y(T8720_Y), .A0(T12416_Y), .A1(T5308_Q),     .B0(T12414_Y), .B1(T1044_Q), .C0(T12417_Y), .C1(T1037_Q),     .D0(T12415_Y), .D1(T1066_Q));
KC_AO2222_X1 T8711 ( .Y(T8711_Y), .A0(T12416_Y), .A1(T5309_Q),     .B0(T12417_Y), .B1(T4858_Q), .C0(T12415_Y), .C1(T5301_Q),     .D0(T12414_Y), .D1(T1048_Q));
KC_AO2222_X1 T8710 ( .Y(T8710_Y), .A0(T12416_Y), .A1(T935_Q),     .B0(T12417_Y), .B1(T1041_Q), .C0(T12415_Y), .C1(T8714_Q),     .D0(T12414_Y), .D1(T1045_Q));
KC_AO2222_X1 T8690 ( .Y(T8690_Y), .A0(T12416_Y), .A1(T724_Q),     .B0(T12417_Y), .B1(T701_Q), .C0(T12414_Y), .C1(T729_Q),     .D0(T12415_Y), .D1(T717_Q));
KC_AO2222_X1 T10127 ( .Y(T10127_Y), .A0(T1363_Y), .A1(T1369_Y),     .B0(T15527_Y), .B1(T1370_Y), .C0(T10129_Y), .C1(T1360_Y),     .D0(T10123_Y), .D1(T10128_Y));
KC_AO2222_X1 T8181 ( .Y(T8181_Y), .A0(T11499_Y), .A1(T16484_Q),     .B0(T5909_Y), .B1(T5429_Q), .C0(T5848_Y), .C1(T15891_Q),     .D0(T12248_Y), .D1(T16486_Q));
KC_AO2222_X1 T8180 ( .Y(T8180_Y), .A0(T11499_Y), .A1(T16485_Q),     .B0(T5909_Y), .B1(T2692_Q), .C0(T5848_Y), .C1(T15880_Q),     .D0(T12248_Y), .D1(T16487_Q));
KC_AO2222_X1 T8270 ( .Y(T8270_Y), .A0(T13128_Q), .A1(T11480_Y),     .B0(T5909_Y), .B1(T4971_Q), .C0(T11499_Y), .C1(T16481_Q),     .D0(T5944_Y), .D1(T2381_Q));
KC_AO2222_X1 T8249 ( .Y(T8249_Y), .A0(T5465_Q), .A1(T11480_Y),     .B0(T5909_Y), .B1(T2115_Q), .C0(T11499_Y), .C1(T1984_Q),     .D0(T5944_Y), .D1(T2385_Q));
KC_AO2222_X1 T8350 ( .Y(T8350_Y), .A0(T2278_Q), .A1(T4965_Y),     .B0(T2843_Q), .B1(T2876_Y), .C0(T12270_Y), .C1(T15815_Q),     .D0(T1820_Q), .D1(T6164_Y));
KC_AO2222_X1 T8159 ( .Y(T8159_Y), .A0(T2369_Y), .A1(T15142_Y),     .B0(T2383_Y), .B1(T2368_Y), .C0(T8156_Y), .C1(T6501_Y),     .D0(T13197_Y), .D1(T8155_Y));
KC_AO2222_X1 T9965 ( .Y(T9965_Y), .A0(T2576_Y), .A1(T2585_Y),     .B0(T9947_Y), .B1(T2562_Y), .C0(T2013_Y), .C1(T2586_Y),     .D0(T16412_Y), .D1(T2587_Y));
KC_AO2222_X1 T8260 ( .Y(T8260_Y), .A0(T3331_Y), .A1(T5011_Y),     .B0(T15960_Y), .B1(T2766_Y), .C0(T15844_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T3921_Y));
KC_AO2222_X1 T8259 ( .Y(T8259_Y), .A0(T3331_Y), .A1(T2765_Y),     .B0(T15960_Y), .B1(T421_Y), .C0(T964_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T2164_Y));
KC_AO2222_X1 T8481 ( .Y(T8481_Y), .A0(T15797_Q), .A1(T11546_Y),     .B0(T3331_Y), .B1(T16452_Y), .C0(T15960_Y), .C1(T3963_Y),     .D0(T15597_Y), .D1(T3338_Y));
KC_AO2222_X1 T8295 ( .Y(T8295_Y), .A0(T3331_Y), .A1(T3330_Y),     .B0(T15960_Y), .B1(T16152_Y), .C0(T15809_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T16456_Y));
KC_AO2222_X1 T8294 ( .Y(T8294_Y), .A0(T3331_Y), .A1(T3876_Y),     .B0(T15960_Y), .B1(T2122_Y), .C0(T15807_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T13142_Y));
KC_AO2222_X1 T8279 ( .Y(T8279_Y), .A0(T3331_Y), .A1(T2787_Y),     .B0(T15960_Y), .B1(T13055_Y), .C0(T15808_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T5012_Y));
KC_AO2222_X1 T8278 ( .Y(T8278_Y), .A0(T3331_Y), .A1(T2808_Y),     .B0(T15960_Y), .B1(T12460_Y), .C0(T5380_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T3992_Y));
KC_AO2222_X1 T8276 ( .Y(T8276_Y), .A0(T3331_Y), .A1(T2767_Y),     .B0(T15960_Y), .B1(T2785_Y), .C0(T15796_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T13139_Y));
KC_AO2222_X1 T8162 ( .Y(T8162_Y), .A0(T2930_Y), .A1(T2947_Y),     .B0(T2376_Y), .B1(T2933_Y), .C0(T2930_Y), .C1(T8154_Y),     .D0(T2930_Y), .D1(T2376_Y));
KC_AO2222_X1 T8223 ( .Y(T8223_Y), .A0(T3269_Y), .A1(T3252_Y),     .B0(T3267_Y), .B1(T3315_Y), .C0(T11455_Y), .C1(T2778_Y),     .D0(T3254_Y), .D1(T10638_Y));
KC_AO2222_X1 T8273 ( .Y(T8273_Y), .A0(T12817_Y), .A1(T16001_Y),     .B0(T3363_Y), .B1(T15591_Y), .C0(T3341_Y), .C1(T3316_Y),     .D0(T3328_Y), .D1(T5965_Y));
KC_AO2222_X1 T8424 ( .Y(T8424_Y), .A0(T6079_Y), .A1(T4169_Q),     .B0(T4176_Q), .B1(T6524_Y), .C0(T4168_Q), .C1(T6043_Y),     .D0(T4179_Q), .D1(T6517_Y));
KC_AO2222_X1 T8262 ( .Y(T8262_Y), .A0(T5884_Y), .A1(T15947_Y),     .B0(T12197_Y), .B1(T10938_Y), .C0(T5934_Y), .C1(T15946_Y),     .D0(T4522_Y), .D1(T11518_Y));
KC_AO2222_X1 T8320 ( .Y(T8320_Y), .A0(T4613_Y), .A1(T4600_Y),     .B0(T4600_Y), .B1(T4611_Y), .C0(T4582_Y), .C1(T4585_Y),     .D0(T4585_Y), .D1(T6019_Y));
KC_AO2222_X1 T9325 ( .Y(T9325_Y), .A0(T12412_Y), .A1(T5559_Q),     .B0(T12413_Y), .B1(T5251_Q), .C0(T12411_Y), .C1(T319_Q),     .D0(T12440_Y), .D1(T167_Q));
KC_AO2222_X1 T9259 ( .Y(T9259_Y), .A0(T12412_Y), .A1(T5239_Q),     .B0(T12413_Y), .B1(T5564_Q), .C0(T12411_Y), .C1(T4823_Q),     .D0(T12440_Y), .D1(T5237_Q));
KC_AO2222_X1 T9344 ( .Y(T9344_Y), .A0(T5305_Q), .A1(T12412_Y),     .B0(T699_Q), .B1(T12440_Y), .C0(T12413_Y), .C1(T5283_Q),     .D0(T12411_Y), .D1(T521_Q));
KC_AO2222_X1 T9321 ( .Y(T9321_Y), .A0(T12412_Y), .A1(T681_Q),     .B0(T12440_Y), .B1(T5276_Q), .C0(T12413_Y), .C1(T5560_Q),     .D0(T12411_Y), .D1(T320_Q));
KC_AO2222_X1 T9320 ( .Y(T9320_Y), .A0(T12412_Y), .A1(T863_Q),     .B0(T12413_Y), .B1(T5264_Q), .C0(T12411_Y), .C1(T862_Q),     .D0(T12440_Y), .D1(T5262_Q));
KC_AO2222_X1 T8171 ( .Y(T8171_Y), .A0(T15645_Y), .A1(T15646_Y),     .B0(T2340_Y), .B1(T15646_Y), .C0(T2365_Y), .C1(T15943_Y),     .D0(T15645_Y), .D1(T2375_Y));
KC_AO2222_X1 T8490 ( .Y(T8490_Y), .A0(T3331_Y), .A1(T4174_Y),     .B0(T15960_Y), .B1(T2760_Y), .C0(T15804_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T2741_Y));
KC_AO2222_X1 T8491 ( .Y(T8491_Y), .A0(T3331_Y), .A1(T16202_Y),     .B0(T15960_Y), .B1(T5569_Y), .C0(T16299_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T12462_Y));
KC_AO2222_X1 T8605 ( .Y(T8605_Y), .A0(T12416_Y), .A1(T5227_Q),     .B0(T12417_Y), .B1(T446_Q), .C0(T12415_Y), .C1(T5240_Q),     .D0(T12414_Y), .D1(T450_Q));
KC_AO2222_X1 T8739 ( .Y(T8739_Y), .A0(T4824_Y), .A1(T8741_Y),     .B0(T1143_Y), .B1(T8740_Y), .C0(T738_Y), .C1(T8697_Y),     .D0(T8742_Y), .D1(T8086_Y));
KC_AO2222_X1 T8722 ( .Y(T8722_Y), .A0(T8703_Y), .A1(T8741_Y),     .B0(T7814_Y), .B1(T8697_Y), .C0(T8742_Y), .C1(T8087_Y),     .D0(T8606_Y), .D1(T8740_Y));
KC_AO2222_X1 T8696 ( .Y(T8696_Y), .A0(T4824_Y), .A1(T8697_Y),     .B0(T8754_Y), .B1(T8741_Y), .C0(T8098_Y), .C1(T8742_Y),     .D0(T9310_Y), .D1(T8740_Y));
KC_AO2222_X1 T8689 ( .Y(T8689_Y), .A0(T12416_Y), .A1(T725_Q),     .B0(T12417_Y), .B1(T713_Q), .C0(T5348_Q), .C1(T12414_Y),     .D0(T716_Q), .D1(T12415_Y));
KC_AO2222_X1 T8833 ( .Y(T8833_Y), .A0(T8917_Y), .A1(T8868_Y),     .B0(T7912_Y), .B1(T8812_Y), .C0(T8867_Y), .C1(T231_Y),     .D0(T8635_Y), .D1(T8811_Y));
KC_AO2222_X1 T8258 ( .Y(T8258_Y), .A0(T3331_Y), .A1(T4177_Y),     .B0(T15960_Y), .B1(T13302_Y), .C0(T15005_Y), .C1(T11546_Y),     .D0(T15597_Y), .D1(T5483_Y));
KC_AO2222_X1 T8480 ( .Y(T8480_Y), .A0(T3331_Y), .A1(T16503_Y),     .B0(T15960_Y), .B1(T5067_Y), .C0(T15805_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T3335_Y));
KC_AO2222_X1 T8293 ( .Y(T8293_Y), .A0(T3331_Y), .A1(T3951_Y),     .B0(T15960_Y), .B1(T12461_Y), .C0(T16088_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T3268_Y));
KC_AO2222_X1 T8285 ( .Y(T8285_Y), .A0(T3331_Y), .A1(T12463_Y),     .B0(T15960_Y), .B1(T3329_Y), .C0(T15803_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T16083_Y));
KC_AO2222_X1 T8277 ( .Y(T8277_Y), .A0(T3331_Y), .A1(T3334_Y),     .B0(T15960_Y), .B1(T3991_Y), .C0(T15798_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T3451_Y));
KC_AO2222_X1 T8161 ( .Y(T8161_Y), .A0(T2930_Y), .A1(T2931_Y),     .B0(T2933_Y), .B1(T5535_Y), .C0(T2376_Y), .C1(T5535_Y),     .D0(T11844_Y), .D1(T8154_Y));
KC_AO2222_X1 T9333 ( .Y(T9333_Y), .A0(T12416_Y), .A1(T709_Q),     .B0(T12417_Y), .B1(T1040_Q), .C0(T12414_Y), .C1(T1046_Q),     .D0(T12415_Y), .D1(T1068_Q));
KC_AO2222_X1 T8489 ( .Y(T8489_Y), .A0(T3331_Y), .A1(T2747_Y),     .B0(T15960_Y), .B1(T3305_Y), .C0(T16301_Q), .C1(T11546_Y),     .D0(T15597_Y), .D1(T3310_Y));
KC_AOI21_X1 T5613 ( .A0(T8546_Y), .Y(T5613_Y), .B(T8544_Y),     .A1(T6862_Y));
KC_AOI21_X1 T5597 ( .A0(T5599_Y), .Y(T5597_Y), .B(T12470_Y),     .A1(T8541_Y));
KC_AOI21_X1 T6967 ( .A0(T6970_Y), .Y(T6967_Y), .B(T12475_Y),     .A1(T6911_Y));
KC_AOI21_X1 T6910 ( .A0(T123_Y), .Y(T6910_Y), .B(T12475_Y),     .A1(T8590_Y));
KC_AOI21_X1 T6909 ( .A0(T8600_Y), .Y(T6909_Y), .B(T12475_Y),     .A1(T6911_Y));
KC_AOI21_X1 T1367 ( .A0(T15490_Y), .Y(T1367_Y), .B(T1378_Y),     .A1(T15091_Y));
KC_AOI21_X1 T8142 ( .A0(T1428_Y), .Y(T8142_Y), .B(T8990_Y),     .A1(T1339_Y));
KC_AOI21_X1 T6316 ( .A0(T12398_Y), .Y(T6316_Y), .B(T13248_Y),     .A1(T156_Y));
KC_AOI21_X1 T6314 ( .A0(T12398_Y), .Y(T6314_Y), .B(T735_Y),     .A1(T7606_Y));
KC_AOI21_X1 T268 ( .A0(T7108_Y), .Y(T268_Y), .B(T13248_Y),     .A1(T6805_Y));
KC_AOI21_X1 T266 ( .A0(T16162_Y), .Y(T266_Y), .B(T735_Y),     .A1(T12398_Y));
KC_AOI21_X1 T6966 ( .A0(T6804_Y), .Y(T6966_Y), .B(T735_Y),     .A1(T7606_Y));
KC_AOI21_X1 T6964 ( .A0(T16162_Y), .Y(T6964_Y), .B(T735_Y),     .A1(T12401_Y));
KC_AOI21_X1 T6943 ( .A0(T284_Q), .Y(T6943_Y), .B(T8575_Y),     .A1(T264_Y));
KC_AOI21_X1 T6941 ( .A0(T12401_Y), .Y(T6941_Y), .B(T735_Y),     .A1(T7606_Y));
KC_AOI21_X1 T6930 ( .A0(T16162_Y), .Y(T6930_Y), .B(T735_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7107 ( .A0(T156_Y), .Y(T7107_Y), .B(T13248_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7106 ( .A0(T12401_Y), .Y(T7106_Y), .B(T13248_Y),     .A1(T156_Y));
KC_AOI21_X1 T7103 ( .A0(T7606_Y), .Y(T7103_Y), .B(T735_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7083 ( .A0(T294_Q), .Y(T7083_Y), .B(T8613_Y),     .A1(T331_Y));
KC_AOI21_X1 T7072 ( .A0(T6804_Y), .Y(T7072_Y), .B(T13248_Y),     .A1(T156_Y));
KC_AOI21_X1 T7071 ( .A0(T5243_Q), .Y(T7071_Y), .B(T8609_Y),     .A1(T15373_Y));
KC_AOI21_X1 T7317 ( .A0(T12398_Y), .Y(T7317_Y), .B(T13249_Y),     .A1(T16376_Y));
KC_AOI21_X1 T7316 ( .A0(T6804_Y), .Y(T7316_Y), .B(T13249_Y),     .A1(T16376_Y));
KC_AOI21_X1 T7315 ( .A0(T16376_Y), .Y(T7315_Y), .B(T13249_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7314 ( .A0(T12401_Y), .Y(T7314_Y), .B(T13249_Y),     .A1(T16376_Y));
KC_AOI21_X1 T7311 ( .A0(T176_Y), .Y(T7311_Y), .B(T13247_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7310 ( .A0(T7812_Y), .Y(T7310_Y), .B(T13249_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7258 ( .A0(T6804_Y), .Y(T7258_Y), .B(T13247_Y),     .A1(T186_Y));
KC_AOI21_X1 T7257 ( .A0(T12401_Y), .Y(T7257_Y), .B(T13247_Y),     .A1(T186_Y));
KC_AOI21_X1 T7256 ( .A0(T12398_Y), .Y(T7256_Y), .B(T13247_Y),     .A1(T186_Y));
KC_AOI21_X1 T7253 ( .A0(T186_Y), .Y(T7253_Y), .B(T13247_Y),     .A1(T6805_Y));
KC_AOI21_X1 T15724 ( .A0(T7813_Y), .Y(T15724_Y), .B(T13242_Y),     .A1(T6805_Y));
KC_AOI21_X1 T15723 ( .A0(T8808_Y), .Y(T15723_Y), .B(T13242_Y),     .A1(T6805_Y));
KC_AOI21_X1 T6814 ( .A0(T6804_Y), .Y(T6814_Y), .B(T13245_Y),     .A1(T214_Y));
KC_AOI21_X1 T6811 ( .A0(T214_Y), .Y(T6811_Y), .B(T13245_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7458 ( .A0(T357_Y), .Y(T7458_Y), .B(T13244_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7457 ( .A0(T6804_Y), .Y(T7457_Y), .B(T13242_Y),     .A1(T8808_Y));
KC_AOI21_X1 T7428 ( .A0(T16429_Y), .Y(T7428_Y), .B(T13243_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7427 ( .A0(T6804_Y), .Y(T7427_Y), .B(T13243_Y),     .A1(T16429_Y));
KC_AOI21_X1 T7426 ( .A0(T10264_Y), .Y(T7426_Y), .B(T13243_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7404 ( .A0(T12398_Y), .Y(T7404_Y), .B(T13243_Y),     .A1(T16429_Y));
KC_AOI21_X1 T7403 ( .A0(T12401_Y), .Y(T7403_Y), .B(T13243_Y),     .A1(T16429_Y));
KC_AOI21_X1 T7389 ( .A0(T12401_Y), .Y(T7389_Y), .B(T13244_Y),     .A1(T15425_Y));
KC_AOI21_X1 T7388 ( .A0(T12398_Y), .Y(T7388_Y), .B(T13244_Y),     .A1(T15425_Y));
KC_AOI21_X1 T7384 ( .A0(T8808_Y), .Y(T7384_Y), .B(T13242_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7383 ( .A0(T15425_Y), .Y(T7383_Y), .B(T13244_Y),     .A1(T6805_Y));
KC_AOI21_X1 T7382 ( .A0(T6804_Y), .Y(T7382_Y), .B(T13244_Y),     .A1(T15425_Y));
KC_AOI21_X1 T7381 ( .A0(T12398_Y), .Y(T7381_Y), .B(T13242_Y),     .A1(T8808_Y));
KC_AOI21_X1 T7576 ( .A0(T382_Y), .Y(T7576_Y), .B(T16334_Y),     .A1(T8720_Y));
KC_AOI21_X1 T7574 ( .A0(T382_Y), .Y(T7574_Y), .B(T8698_Y),     .A1(T8637_Y));
KC_AOI21_X1 T16390 ( .A0(T371_Y), .Y(T16390_Y), .B(T9424_Y),     .A1(T8638_Y));
KC_AOI21_X1 T16330 ( .A0(T382_Y), .Y(T16330_Y), .B(T16329_Y),     .A1(T612_Y));
KC_AOI21_X1 T16326 ( .A0(T7827_Y), .Y(T16326_Y), .B(T7570_Y),     .A1(T9388_Y));
KC_AOI21_X1 T7909 ( .A0(T371_Y), .Y(T7909_Y), .B(T970_Y),     .A1(T8711_Y));
KC_AOI21_X1 T7908 ( .A0(T371_Y), .Y(T7908_Y), .B(T8866_Y),     .A1(T9259_Y));
KC_AOI21_X1 T8097 ( .A0(T8078_Y), .Y(T8097_Y), .B(T7857_Y),     .A1(T7917_Y));
KC_AOI21_X1 T8076 ( .A0(T371_Y), .Y(T8076_Y), .B(T1272_Y),     .A1(T613_Y));
KC_AOI21_X1 T6861 ( .A0(T272_Q), .Y(T6861_Y), .B(T9295_Y),     .A1(T217_Y));
KC_AOI21_X1 T6305 ( .A0(T273_Q), .Y(T6305_Y), .B(T9265_Y),     .A1(T285_Y));
KC_AOI21_X1 T6965 ( .A0(T283_Q), .Y(T6965_Y), .B(T8587_Y),     .A1(T15357_Y));
KC_AOI21_X1 T6960 ( .A0(T7318_Y), .Y(T6960_Y), .B(T721_Y),     .A1(T9313_Y));
KC_AOI21_X1 T6959 ( .A0(T6809_Y), .Y(T6959_Y), .B(T733_Y),     .A1(T9313_Y));
KC_AOI21_X1 T6958 ( .A0(T9312_Y), .Y(T6958_Y), .B(T733_Y),     .A1(T7810_Y));
KC_AOI21_X1 T6957 ( .A0(T9312_Y), .Y(T6957_Y), .B(T721_Y),     .A1(T472_Y));
KC_AOI21_X1 T6942 ( .A0(T278_Q), .Y(T6942_Y), .B(T8586_Y),     .A1(T251_Y));
KC_AOI21_X1 T6927 ( .A0(T12398_Y), .Y(T6927_Y), .B(T733_Y),     .A1(T7810_Y));
KC_AOI21_X1 T6926 ( .A0(T12398_Y), .Y(T6926_Y), .B(T721_Y),     .A1(T472_Y));
KC_AOI21_X1 T6908 ( .A0(T6809_Y), .Y(T6908_Y), .B(T733_Y),     .A1(T692_Y));
KC_AOI21_X1 T6907 ( .A0(T692_Y), .Y(T6907_Y), .B(T733_Y),     .A1(T7810_Y));
KC_AOI21_X1 T6906 ( .A0(T692_Y), .Y(T6906_Y), .B(T721_Y), .A1(T472_Y));
KC_AOI21_X1 T6905 ( .A0(T7318_Y), .Y(T6905_Y), .B(T721_Y),     .A1(T692_Y));
KC_AOI21_X1 T6345 ( .A0(T7108_Y), .Y(T6345_Y), .B(T13248_Y),     .A1(T12401_Y));
KC_AOI21_X1 T6343 ( .A0(T6804_Y), .Y(T6343_Y), .B(T733_Y),     .A1(T6809_Y));
KC_AOI21_X1 T7096 ( .A0(T274_Q), .Y(T7096_Y), .B(T9257_Y),     .A1(T342_Y));
KC_AOI21_X1 T7095 ( .A0(T472_Y), .Y(T7095_Y), .B(T721_Y),     .A1(T6805_Y));
KC_AOI21_X1 T6732 ( .A0(T6804_Y), .Y(T6732_Y), .B(T13249_Y),     .A1(T7812_Y));
KC_AOI21_X1 T6731 ( .A0(T15028_Y), .Y(T6731_Y), .B(T13245_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7305 ( .A0(T176_Y), .Y(T7305_Y), .B(T13247_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7287 ( .A0(T6804_Y), .Y(T7287_Y), .B(T13247_Y),     .A1(T176_Y));
KC_AOI21_X1 T7286 ( .A0(T7812_Y), .Y(T7286_Y), .B(T13249_Y),     .A1(T12398_Y));
KC_AOI21_X1 T7282 ( .A0(T176_Y), .Y(T7282_Y), .B(T13247_Y),     .A1(T12398_Y));
KC_AOI21_X1 T7267 ( .A0(T7812_Y), .Y(T7267_Y), .B(T13249_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7248 ( .A0(T6804_Y), .Y(T7248_Y), .B(T13248_Y),     .A1(T7108_Y));
KC_AOI21_X1 T7450 ( .A0(T357_Y), .Y(T7450_Y), .B(T13244_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7449 ( .A0(T357_Y), .Y(T7449_Y), .B(T13244_Y),     .A1(T12398_Y));
KC_AOI21_X1 T7375 ( .A0(T10264_Y), .Y(T7375_Y), .B(T13243_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7374 ( .A0(T10264_Y), .Y(T7374_Y), .B(T13243_Y),     .A1(T12398_Y));
KC_AOI21_X1 T7688 ( .A0(T382_Y), .Y(T7688_Y), .B(T8752_Y),     .A1(T9310_Y));
KC_AOI21_X1 T7575 ( .A0(T382_Y), .Y(T7575_Y), .B(T8753_Y),     .A1(T8651_Y));
KC_AOI21_X1 T16391 ( .A0(T371_Y), .Y(T16391_Y), .B(T9421_Y),     .A1(T9320_Y));
KC_AOI21_X1 T16385 ( .A0(T16310_Y), .Y(T16385_Y), .B(T8943_Y),     .A1(T8041_Y));
KC_AOI21_X1 T1417 ( .A0(T13259_Y), .Y(T1417_Y), .B(T12888_Y),     .A1(T1426_Y));
KC_AOI21_X1 T8069 ( .A0(T8940_Y), .Y(T8069_Y), .B(T12720_Y),     .A1(T7901_Y));
KC_AOI21_X1 T8044 ( .A0(T16385_Y), .Y(T8044_Y), .B(T12720_Y),     .A1(T8909_Y));
KC_AOI21_X1 T1839 ( .A0(T8123_Y), .Y(T1839_Y), .B(T1594_Y),     .A1(T9112_Y));
KC_AOI21_X1 T5335 ( .A0(T4842_Y), .Y(T5335_Y), .B(T9166_Y),     .A1(T9193_Y));
KC_AOI21_X1 T5307 ( .A0(T567_Q), .Y(T5307_Y), .B(T13265_Y),     .A1(T9476_Y));
KC_AOI21_X1 T216 ( .A0(T1279_Y), .Y(T216_Y), .B(T9166_Y),     .A1(T15538_Y));
KC_AOI21_X1 T6951 ( .A0(T6350_Y), .Y(T6951_Y), .B(T16427_Y),     .A1(T9313_Y));
KC_AOI21_X1 T6900 ( .A0(T6350_Y), .Y(T6900_Y), .B(T16427_Y),     .A1(T692_Y));
KC_AOI21_X1 T15730 ( .A0(T7813_Y), .Y(T15730_Y), .B(T13242_Y),     .A1(T9334_Y));
KC_AOI21_X1 T7451 ( .A0(T6804_Y), .Y(T7451_Y), .B(T13242_Y),     .A1(T7813_Y));
KC_AOI21_X1 T7444 ( .A0(T7813_Y), .Y(T7444_Y), .B(T13242_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7392 ( .A0(T6804_Y), .Y(T7392_Y), .B(T13245_Y),     .A1(T15028_Y));
KC_AOI21_X1 T7652 ( .A0(T16352_Y), .Y(T7652_Y), .B(T931_Y),     .A1(T7803_Y));
KC_AOI21_X1 T7651 ( .A0(T16353_Y), .Y(T7651_Y), .B(T931_Y),     .A1(T16351_Y));
KC_AOI21_X1 T7650 ( .A0(T16347_Y), .Y(T7650_Y), .B(T931_Y),     .A1(T16349_Y));
KC_AOI21_X1 T7642 ( .A0(T703_Y), .Y(T7642_Y), .B(T16425_Y),     .A1(T690_Q));
KC_AOI21_X1 T7640 ( .A0(T16348_Y), .Y(T7640_Y), .B(T931_Y),     .A1(T16350_Y));
KC_AOI21_X1 T16386 ( .A0(T9416_Y), .Y(T16386_Y), .B(T8903_Y),     .A1(T1255_Y));
KC_AOI21_X1 T8036 ( .A0(T8905_Y), .Y(T8036_Y), .B(T9096_Y),     .A1(T16387_Y));
KC_AOI21_X1 T8035 ( .A0(T8072_Y), .Y(T8035_Y), .B(T5608_Y),     .A1(T8117_Y));
KC_AOI21_X1 T6274 ( .A0(T9334_Y), .Y(T6274_Y), .B(T732_Y),     .A1(T7607_Y));
KC_AOI21_X1 T6269 ( .A0(T15731_Y), .Y(T6269_Y), .B(T732_Y),     .A1(T9334_Y));
KC_AOI21_X1 T6952 ( .A0(T692_Y), .Y(T6952_Y), .B(T16427_Y),     .A1(T7603_Y));
KC_AOI21_X1 T6950 ( .A0(T15731_Y), .Y(T6950_Y), .B(T732_Y),     .A1(T692_Y));
KC_AOI21_X1 T6949 ( .A0(T9312_Y), .Y(T6949_Y), .B(T16427_Y),     .A1(T7603_Y));
KC_AOI21_X1 T6937 ( .A0(T692_Y), .Y(T6937_Y), .B(T732_Y),     .A1(T7607_Y));
KC_AOI21_X1 T6936 ( .A0(T15731_Y), .Y(T6936_Y), .B(T732_Y),     .A1(T9313_Y));
KC_AOI21_X1 T6918 ( .A0(T9312_Y), .Y(T6918_Y), .B(T732_Y),     .A1(T7607_Y));
KC_AOI21_X1 T7111 ( .A0(T7607_Y), .Y(T7111_Y), .B(T732_Y),     .A1(T9313_Y));
KC_AOI21_X1 T7092 ( .A0(T9312_Y), .Y(T7092_Y), .B(T732_Y),     .A1(T15731_Y));
KC_AOI21_X1 T7091 ( .A0(T7603_Y), .Y(T7091_Y), .B(T16427_Y),     .A1(T9313_Y));
KC_AOI21_X1 T7049 ( .A0(T6350_Y), .Y(T7049_Y), .B(T16427_Y),     .A1(T9334_Y));
KC_AOI21_X1 T7281 ( .A0(T16382_Y), .Y(T7281_Y), .B(T16426_Y),     .A1(T9313_Y));
KC_AOI21_X1 T7279 ( .A0(T736_Y), .Y(T7279_Y), .B(T16426_Y),     .A1(T12401_Y));
KC_AOI21_X1 T7278 ( .A0(T9312_Y), .Y(T7278_Y), .B(T16426_Y),     .A1(T16382_Y));
KC_AOI21_X1 T7262 ( .A0(T736_Y), .Y(T7262_Y), .B(T16426_Y),     .A1(T9334_Y));
KC_AOI21_X1 T7260 ( .A0(T736_Y), .Y(T7260_Y), .B(T16426_Y),     .A1(T9313_Y));
KC_AOI21_X1 T7259 ( .A0(T12401_Y), .Y(T7259_Y), .B(T16426_Y),     .A1(T16382_Y));
KC_AOI21_X1 T15745 ( .A0(T7637_Y), .Y(T15745_Y), .B(T6691_Y),     .A1(T919_Y));
KC_AOI21_X1 T7442 ( .A0(T552_Y), .Y(T7442_Y), .B(T16425_Y),     .A1(T697_Q));
KC_AOI21_X1 T7437 ( .A0(T497_Y), .Y(T7437_Y), .B(T929_Y), .A1(T909_Y));
KC_AOI21_X1 T7436 ( .A0(T548_Y), .Y(T7436_Y), .B(T16425_Y),     .A1(T7367_Q));
KC_AOI21_X1 T7435 ( .A0(T7637_Y), .Y(T7435_Y), .B(T497_Y),     .A1(T919_Y));
KC_AOI21_X1 T7415 ( .A0(T909_Y), .Y(T7415_Y), .B(T15770_Y),     .A1(T549_Y));
KC_AOI21_X1 T7363 ( .A0(T909_Y), .Y(T7363_Y), .B(T15770_Y),     .A1(T6691_Y));
KC_AOI21_X1 T7358 ( .A0(T545_Y), .Y(T7358_Y), .B(T16425_Y),     .A1(T5280_Q));
KC_AOI21_X1 T7357 ( .A0(T9370_Y), .Y(T7357_Y), .B(T929_Y),     .A1(T909_Y));
KC_AOI21_X1 T7356 ( .A0(T7637_Y), .Y(T7356_Y), .B(T549_Y),     .A1(T919_Y));
KC_AOI21_X1 T7683 ( .A0(T11181_Y), .Y(T7683_Y), .B(T15763_Y),     .A1(T9374_Y));
KC_AOI21_X1 T7641 ( .A0(T16163_Y), .Y(T7641_Y), .B(T16425_Y),     .A1(T698_Q));
KC_AOI21_X1 T7632 ( .A0(T7637_Y), .Y(T7632_Y), .B(T9374_Y),     .A1(T919_Y));
KC_AOI21_X1 T7631 ( .A0(T7637_Y), .Y(T7631_Y), .B(T727_Y),     .A1(T919_Y));
KC_AOI21_X1 T7630 ( .A0(T15223_Y), .Y(T7630_Y), .B(T7614_Y),     .A1(T15454_Y));
KC_AOI21_X1 T7596 ( .A0(T660_Y), .Y(T7596_Y), .B(T16425_Y),     .A1(T683_Q));
KC_AOI21_X1 T7587 ( .A0(T7637_Y), .Y(T7587_Y), .B(T9373_Y),     .A1(T919_Y));
KC_AOI21_X1 T7561 ( .A0(T11181_Y), .Y(T7561_Y), .B(T15763_Y),     .A1(T727_Y));
KC_AOI21_X1 T7560 ( .A0(T11181_Y), .Y(T7560_Y), .B(T15767_Y),     .A1(T9373_Y));
KC_AOI21_X1 T7554 ( .A0(T910_Q), .Y(T7554_Y), .B(T5309_Q),     .A1(T7558_Y));
KC_AOI21_X1 T7553 ( .A0(T11181_Y), .Y(T7553_Y), .B(T15767_Y),     .A1(T637_Y));
KC_AOI21_X1 T7875 ( .A0(T7846_Y), .Y(T7875_Y), .B(T12884_Y),     .A1(T9404_Y));
KC_AOI21_X1 T7800 ( .A0(T8792_Y), .Y(T7800_Y), .B(T8759_Y),     .A1(T15654_Y));
KC_AOI21_X1 T7549 ( .A0(T5359_Q), .Y(T7549_Y), .B(T1048_Q),     .A1(T7741_Y));
KC_AOI21_X1 T7634 ( .A0(T9507_Y), .Y(T7634_Y), .B(T11880_Y),     .A1(T15433_Y));
KC_AOI21_X1 T7633 ( .A0(T9503_Y), .Y(T7633_Y), .B(T11918_Y),     .A1(T718_Y));
KC_AOI21_X1 T7612 ( .A0(T5343_Q), .Y(T7612_Y), .B(T5301_Q),     .A1(T7638_Y));
KC_AOI21_X1 T7588 ( .A0(T9506_Y), .Y(T7588_Y), .B(T11193_Y),     .A1(T16381_Y));
KC_AOI21_X1 T7949 ( .A0(T8032_Y), .Y(T7949_Y), .B(T9891_Y),     .A1(T980_Q));
KC_AOI21_X1 T10737 ( .A0(T10315_Y), .Y(T10737_Y), .B(T10021_Y),     .A1(T7951_Y));
KC_AOI21_X1 T10652 ( .A0(T1586_Y), .Y(T10652_Y), .B(T16437_Y),     .A1(T7942_Y));
KC_AOI21_X1 T8017 ( .A0(T1586_Y), .Y(T8017_Y), .B(T16437_Y),     .A1(T7975_Y));
KC_AOI21_X1 T10725 ( .A0(T1738_Y), .Y(T10725_Y), .B(T1357_Y),     .A1(T4819_Y));
KC_AOI21_X1 T7217 ( .A0(T10263_Y), .Y(T7217_Y), .B(T6771_Y),     .A1(T7036_Y));
KC_AOI21_X1 T7194 ( .A0(T10263_Y), .Y(T7194_Y), .B(T6771_Y),     .A1(T7235_Y));
KC_AOI21_X1 T7193 ( .A0(T10263_Y), .Y(T7193_Y), .B(T6771_Y),     .A1(T7160_Y));
KC_AOI21_X1 T7191 ( .A0(T10263_Y), .Y(T7191_Y), .B(T6771_Y),     .A1(T6997_Y));
KC_AOI21_X1 T7181 ( .A0(T10263_Y), .Y(T7181_Y), .B(T6771_Y),     .A1(T7151_Y));
KC_AOI21_X1 T7180 ( .A0(T10263_Y), .Y(T7180_Y), .B(T6771_Y),     .A1(T7227_Y));
KC_AOI21_X1 T7143 ( .A0(T10263_Y), .Y(T7143_Y), .B(T6771_Y),     .A1(T7233_Y));
KC_AOI21_X1 T7142 ( .A0(T10263_Y), .Y(T7142_Y), .B(T6771_Y),     .A1(T7236_Y));
KC_AOI21_X1 T7138 ( .A0(T10263_Y), .Y(T7138_Y), .B(T6771_Y),     .A1(T10391_Y));
KC_AOI21_X1 T7137 ( .A0(T10263_Y), .Y(T7137_Y), .B(T6771_Y),     .A1(T7159_Y));
KC_AOI21_X1 T7136 ( .A0(T10263_Y), .Y(T7136_Y), .B(T6771_Y),     .A1(T6984_Y));
KC_AOI21_X1 T7135 ( .A0(T10263_Y), .Y(T7135_Y), .B(T6771_Y),     .A1(T7017_Y));
KC_AOI21_X1 T7134 ( .A0(T10263_Y), .Y(T7134_Y), .B(T6771_Y),     .A1(T7026_Y));
KC_AOI21_X1 T7133 ( .A0(T10263_Y), .Y(T7133_Y), .B(T6771_Y),     .A1(T7232_Y));
KC_AOI21_X1 T7349 ( .A0(T10263_Y), .Y(T7349_Y), .B(T15462_Y),     .A1(T5662_Y));
KC_AOI21_X1 T5672 ( .A0(T2564_Y), .Y(T5672_Y), .B(T6771_Y),     .A1(T5701_Y));
KC_AOI21_X1 T5671 ( .A0(T16164_Y), .Y(T5671_Y), .B(T6771_Y),     .A1(T5681_Y));
KC_AOI21_X1 T5670 ( .A0(T2564_Y), .Y(T5670_Y), .B(T6771_Y),     .A1(T7496_Y));
KC_AOI21_X1 T5669 ( .A0(T2564_Y), .Y(T5669_Y), .B(T15462_Y),     .A1(T10373_Y));
KC_AOI21_X1 T7540 ( .A0(T2564_Y), .Y(T7540_Y), .B(T15462_Y),     .A1(T7548_Y));
KC_AOI21_X1 T7509 ( .A0(T16164_Y), .Y(T7509_Y), .B(T15462_Y),     .A1(T5695_Y));
KC_AOI21_X1 T7793 ( .A0(T1586_Y), .Y(T7793_Y), .B(T16437_Y),     .A1(T7776_Y));
KC_AOI21_X1 T7789 ( .A0(T2564_Y), .Y(T7789_Y), .B(T15462_Y),     .A1(T7738_Y));
KC_AOI21_X1 T7788 ( .A0(T1586_Y), .Y(T7788_Y), .B(T16437_Y),     .A1(T9790_Y));
KC_AOI21_X1 T7787 ( .A0(T1586_Y), .Y(T7787_Y), .B(T16437_Y),     .A1(T7739_Y));
KC_AOI21_X1 T7786 ( .A0(T16164_Y), .Y(T7786_Y), .B(T15462_Y),     .A1(T10338_Y));
KC_AOI21_X1 T7701 ( .A0(T1586_Y), .Y(T7701_Y), .B(T16437_Y),     .A1(T7717_Y));
KC_AOI21_X1 T7700 ( .A0(T1586_Y), .Y(T7700_Y), .B(T16437_Y),     .A1(T7711_Y));
KC_AOI21_X1 T10760 ( .A0(T1586_Y), .Y(T10760_Y), .B(T16437_Y),     .A1(T7991_Y));
KC_AOI21_X1 T8013 ( .A0(T1586_Y), .Y(T8013_Y), .B(T16437_Y),     .A1(T7935_Y));
KC_AOI21_X1 T7971 ( .A0(T1586_Y), .Y(T7971_Y), .B(T16437_Y),     .A1(T7945_Y));
KC_AOI21_X1 T7963 ( .A0(T1586_Y), .Y(T7963_Y), .B(T16437_Y),     .A1(T10012_Y));
KC_AOI21_X1 T7962 ( .A0(T1586_Y), .Y(T7962_Y), .B(T16437_Y),     .A1(T7934_Y));
KC_AOI21_X1 T7961 ( .A0(T1586_Y), .Y(T7961_Y), .B(T16437_Y),     .A1(T9999_Y));
KC_AOI21_X1 T7960 ( .A0(T1586_Y), .Y(T7960_Y), .B(T16437_Y),     .A1(T9997_Y));
KC_AOI21_X1 T7953 ( .A0(T1586_Y), .Y(T7953_Y), .B(T16437_Y),     .A1(T7928_Y));
KC_AOI21_X1 T7177 ( .A0(T10263_Y), .Y(T7177_Y), .B(T6771_Y),     .A1(T7219_Y));
KC_AOI21_X1 T7176 ( .A0(T10263_Y), .Y(T7176_Y), .B(T6771_Y),     .A1(T7010_Y));
KC_AOI21_X1 T7778 ( .A0(T4919_Y), .Y(T7778_Y), .B(T835_Y),     .A1(T10757_Y));
KC_AOI21_X1 T8010 ( .A0(T16164_Y), .Y(T8010_Y), .B(T15462_Y),     .A1(T9994_Y));
KC_AOI21_X1 T7956 ( .A0(T1586_Y), .Y(T7956_Y), .B(T16437_Y),     .A1(T9992_Y));
KC_AOI21_X1 T7955 ( .A0(T1586_Y), .Y(T7955_Y), .B(T16437_Y),     .A1(T10010_Y));
KC_AOI21_X1 T7954 ( .A0(T1586_Y), .Y(T7954_Y), .B(T16437_Y),     .A1(T10310_Y));
KC_AOI21_X1 T6191 ( .A0(T5899_Y), .Y(T6191_Y), .B(T11494_Y),     .A1(T5911_Y));
KC_AOI21_X1 T6303 ( .A0(T10225_Y), .Y(T6303_Y), .B(T6006_Y),     .A1(T15973_Y));
KC_AOI21_X1 T6522 ( .A0(T2958_Y), .Y(T6522_Y), .B(T11766_Y),     .A1(T6199_Y));
KC_AOI21_X1 T6519 ( .A0(T2399_Y), .Y(T6519_Y), .B(T11766_Y),     .A1(T6201_Y));
KC_AOI21_X1 T6518 ( .A0(T6201_Y), .Y(T6518_Y), .B(T11766_Y),     .A1(T6199_Y));
KC_AOI21_X1 T5891 ( .A0(T868_Y), .Y(T5891_Y), .B(T11260_Y),     .A1(T2161_Q));
KC_AOI21_X1 T5881 ( .A0(T11949_Y), .Y(T5881_Y), .B(T10524_Y),     .A1(T1124_Y));
KC_AOI21_X1 T6280 ( .A0(T11586_Y), .Y(T6280_Y), .B(T12818_Y),     .A1(T15952_Y));
KC_AOI21_X1 T6273 ( .A0(T11586_Y), .Y(T6273_Y), .B(T12822_Y),     .A1(T2129_Q));
KC_AOI21_X1 T6817 ( .A0(T2315_Q), .Y(T6817_Y), .B(T13267_Y),     .A1(T6464_Y));
KC_AOI21_X1 T6404 ( .A0(T6419_Q), .Y(T6404_Y), .B(T13310_Y),     .A1(T12269_Y));
KC_AOI21_X1 T6388 ( .A0(T5494_Q), .Y(T6388_Y), .B(T13159_Y),     .A1(T12269_Y));
KC_AOI21_X1 T6387 ( .A0(T12270_Y), .Y(T6387_Y), .B(T13158_Y),     .A1(T1785_Q));
KC_AOI21_X1 T6370 ( .A0(T5571_Q), .Y(T6370_Y), .B(T13157_Y),     .A1(T12269_Y));
KC_AOI21_X1 T6464 ( .A0(T3482_Y), .Y(T6464_Y), .B(T2854_Y),     .A1(T2862_Y));
KC_AOI21_X1 T6588 ( .A0(T2349_Y), .Y(T6588_Y), .B(T2321_Y),     .A1(T2343_Y));
KC_AOI21_X1 T6523 ( .A0(T11772_Y), .Y(T6523_Y), .B(T1832_Q),     .A1(T6200_Y));
KC_AOI21_X1 T6521 ( .A0(T2364_Q), .Y(T6521_Y), .B(T2337_Y),     .A1(T11749_Y));
KC_AOI21_X1 T6632 ( .A0(T14984_Y), .Y(T6632_Y), .B(T6760_Y),     .A1(T3579_Y));
KC_AOI21_X1 T5805 ( .A0(T14995_Y), .Y(T5805_Y), .B(T6760_Y),     .A1(T10369_Y));
KC_AOI21_X1 T5792 ( .A0(T14995_Y), .Y(T5792_Y), .B(T6760_Y),     .A1(T4252_Y));
KC_AOI21_X1 T5847 ( .A0(T14995_Y), .Y(T5847_Y), .B(T875_Y),     .A1(T5083_Y));
KC_AOI21_X1 T5841 ( .A0(T14995_Y), .Y(T5841_Y), .B(T875_Y),     .A1(T4231_Y));
KC_AOI21_X1 T5839 ( .A0(T14995_Y), .Y(T5839_Y), .B(T875_Y),     .A1(T3627_Y));
KC_AOI21_X1 T5887 ( .A0(T14995_Y), .Y(T5887_Y), .B(T875_Y),     .A1(T5322_Y));
KC_AOI21_X1 T5886 ( .A0(T2564_Y), .Y(T5886_Y), .B(T875_Y),     .A1(T12089_Y));
KC_AOI21_X1 T5883 ( .A0(T2564_Y), .Y(T5883_Y), .B(T875_Y),     .A1(T4291_Y));
KC_AOI21_X1 T5866 ( .A0(T2564_Y), .Y(T5866_Y), .B(T875_Y),     .A1(T3137_Y));
KC_AOI21_X1 T5864 ( .A0(T14995_Y), .Y(T5864_Y), .B(T875_Y),     .A1(T3685_Y));
KC_AOI21_X1 T5856 ( .A0(T14995_Y), .Y(T5856_Y), .B(T875_Y),     .A1(T3713_Y));
KC_AOI21_X1 T5935 ( .A0(T2564_Y), .Y(T5935_Y), .B(T875_Y),     .A1(T3129_Y));
KC_AOI21_X1 T5920 ( .A0(T2598_Y), .Y(T5920_Y), .B(T1509_Y),     .A1(T2608_Y));
KC_AOI21_X1 T5979 ( .A0(T2640_Q), .Y(T5979_Y), .B(T4898_Y),     .A1(T2672_Y));
KC_AOI21_X1 T5962 ( .A0(T2564_Y), .Y(T5962_Y), .B(T15532_Y),     .A1(T3761_Y));
KC_AOI21_X1 T5961 ( .A0(T2564_Y), .Y(T5961_Y), .B(T15532_Y),     .A1(T3166_Y));
KC_AOI21_X1 T5960 ( .A0(T2564_Y), .Y(T5960_Y), .B(T15532_Y),     .A1(T3763_Y));
KC_AOI21_X1 T5959 ( .A0(T2564_Y), .Y(T5959_Y), .B(T15532_Y),     .A1(T3742_Y));
KC_AOI21_X1 T5951 ( .A0(T2564_Y), .Y(T5951_Y), .B(T15532_Y),     .A1(T3739_Y));
KC_AOI21_X1 T5950 ( .A0(T2564_Y), .Y(T5950_Y), .B(T15532_Y),     .A1(T3161_Y));
KC_AOI21_X1 T6017 ( .A0(T14954_Q), .Y(T6017_Y), .B(T10243_Y),     .A1(T10242_Y));
KC_AOI21_X1 T6063 ( .A0(T14525_Q), .Y(T6063_Y), .B(T15849_Y),     .A1(T2681_Y));
KC_AOI21_X1 T6061 ( .A0(T14526_Q), .Y(T6061_Y), .B(T11357_Y),     .A1(T5784_Y));
KC_AOI21_X1 T6037 ( .A0(T15696_Y), .Y(T6037_Y), .B(T15753_Y),     .A1(T5425_Q));
KC_AOI21_X1 T6186 ( .A0(T11490_Y), .Y(T6186_Y), .B(T3311_Y),     .A1(T11489_Y));
KC_AOI21_X1 T6295 ( .A0(T3335_Y), .Y(T6295_Y), .B(T2770_Y),     .A1(T5877_Y));
KC_AOI21_X1 T6399 ( .A0(T2630_Y), .Y(T6399_Y), .B(T6431_Q),     .A1(T6088_Y));
KC_AOI21_X1 T6383 ( .A0(T6119_Y), .Y(T6383_Y), .B(T2841_Q),     .A1(T6039_Y));
KC_AOI21_X1 T6493 ( .A0(T2906_Y), .Y(T6493_Y), .B(T3418_Y),     .A1(T16101_Y));
KC_AOI21_X1 T6478 ( .A0(T12285_Y), .Y(T6478_Y), .B(T2870_Y),     .A1(T2871_Y));
KC_AOI21_X1 T6513 ( .A0(T2325_Y), .Y(T6513_Y), .B(T5517_Y),     .A1(T10980_Y));
KC_AOI21_X1 T2931 ( .A0(T6491_Y), .Y(T2931_Y), .B(T6516_Y),     .A1(T2933_Y));
KC_AOI21_X1 T6637 ( .A0(T14984_Y), .Y(T6637_Y), .B(T6760_Y),     .A1(T5033_Y));
KC_AOI21_X1 T6636 ( .A0(T14984_Y), .Y(T6636_Y), .B(T6760_Y),     .A1(T3536_Y));
KC_AOI21_X1 T6635 ( .A0(T14984_Y), .Y(T6635_Y), .B(T6760_Y),     .A1(T3001_Y));
KC_AOI21_X1 T6634 ( .A0(T14984_Y), .Y(T6634_Y), .B(T6760_Y),     .A1(T2981_Y));
KC_AOI21_X1 T6633 ( .A0(T14984_Y), .Y(T6633_Y), .B(T6760_Y),     .A1(T2973_Y));
KC_AOI21_X1 T6631 ( .A0(T14984_Y), .Y(T6631_Y), .B(T6760_Y),     .A1(T3565_Y));
KC_AOI21_X1 T5752 ( .A0(T14984_Y), .Y(T5752_Y), .B(T6760_Y),     .A1(T3587_Y));
KC_AOI21_X1 T5811 ( .A0(T14995_Y), .Y(T5811_Y), .B(T15532_Y),     .A1(T5268_Y));
KC_AOI21_X1 T5865 ( .A0(T2564_Y), .Y(T5865_Y), .B(T875_Y),     .A1(T3082_Y));
KC_AOI21_X1 T6014 ( .A0(T14516_Q), .Y(T6014_Y), .B(T10266_Y),     .A1(T14515_Q));
KC_AOI21_X1 T6726 ( .A0(T12951_Y), .Y(T6726_Y), .B(T12776_Y),     .A1(T15819_Y));
KC_AOI21_X1 T6059 ( .A0(T11394_Y), .Y(T6059_Y), .B(T11335_Y),     .A1(T5431_Y));
KC_AOI21_X1 T6058 ( .A0(T11379_Y), .Y(T6058_Y), .B(T3202_Y),     .A1(T11370_Y));
KC_AOI21_X1 T6109 ( .A0(T15010_Y), .Y(T6109_Y), .B(T11412_Y),     .A1(T14544_Q));
KC_AOI21_X1 T6163 ( .A0(T5871_Y), .Y(T6163_Y), .B(T3252_Y),     .A1(T3267_Y));
KC_AOI21_X1 T6206 ( .A0(T3286_Y), .Y(T6206_Y), .B(T3287_Y),     .A1(T8257_Y));
KC_AOI21_X1 T6256 ( .A0(T16001_Y), .Y(T6256_Y), .B(T5964_Y),     .A1(T5964_Y));
KC_AOI21_X1 T6335 ( .A0(T3361_Y), .Y(T6335_Y), .B(T16015_Y),     .A1(T15607_Y));
KC_AOI21_X1 T6806 ( .A0(T15233_Y), .Y(T6806_Y), .B(T11663_Y),     .A1(T6083_Y));
KC_AOI21_X1 T6393 ( .A0(T10590_Y), .Y(T6393_Y), .B(T5052_Y),     .A1(T11997_Y));
KC_AOI21_X1 T6392 ( .A0(T15615_Y), .Y(T6392_Y), .B(T10962_Y),     .A1(T12253_Y));
KC_AOI21_X1 T6365 ( .A0(T6123_Y), .Y(T6365_Y), .B(T12002_Y),     .A1(T16139_Y));
KC_AOI21_X1 T6440 ( .A0(T15234_Y), .Y(T6440_Y), .B(T6124_Y),     .A1(T3443_Y));
KC_AOI21_X1 T6436 ( .A0(T10583_Y), .Y(T6436_Y), .B(T12845_Y),     .A1(T10587_Y));
KC_AOI21_X1 T6575 ( .A0(T6585_Y), .Y(T6575_Y), .B(T10568_Y),     .A1(T10996_Y));
KC_AOI21_X1 T6558 ( .A0(T11818_Y), .Y(T6558_Y), .B(T10990_Y),     .A1(T3495_Y));
KC_AOI21_X1 T6720 ( .A0(T3790_Y), .Y(T6720_Y), .B(T3202_Y),     .A1(T15835_Y));
KC_AOI21_X1 T6053 ( .A0(T4391_Y), .Y(T6053_Y), .B(T15867_Y),     .A1(T5772_Y));
KC_AOI21_X1 T6041 ( .A0(T3802_Y), .Y(T6041_Y), .B(T5780_Y),     .A1(T3803_Y));
KC_AOI21_X1 T6032 ( .A0(T3790_Y), .Y(T6032_Y), .B(T3202_Y),     .A1(T15825_Y));
KC_AOI21_X1 T6117 ( .A0(T15908_Y), .Y(T6117_Y), .B(T11423_Y),     .A1(T11426_Y));
KC_AOI21_X1 T6116 ( .A0(T10921_Y), .Y(T6116_Y), .B(T16154_Y),     .A1(T10920_Y));
KC_AOI21_X1 T6108 ( .A0(T15865_Y), .Y(T6108_Y), .B(T13092_Y),     .A1(T13093_Y));
KC_AOI21_X1 T6228 ( .A0(T5981_Y), .Y(T6228_Y), .B(T11587_Y),     .A1(T3913_Y));
KC_AOI21_X1 T6204 ( .A0(T11476_Y), .Y(T6204_Y), .B(T5459_Y),     .A1(T5989_Y));
KC_AOI21_X1 T6277 ( .A0(T5963_Y), .Y(T6277_Y), .B(T3950_Y),     .A1(T3883_Q));
KC_AOI21_X1 T6265 ( .A0(T4474_Y), .Y(T6265_Y), .B(T5457_Y),     .A1(T11533_Y));
KC_AOI21_X1 T6251 ( .A0(T4577_Y), .Y(T6251_Y), .B(T5981_Y),     .A1(T4517_Y));
KC_AOI21_X1 T6437 ( .A0(T16143_Y), .Y(T6437_Y), .B(T6080_Y),     .A1(T4027_Y));
KC_AOI21_X1 T6557 ( .A0(T8503_Y), .Y(T6557_Y), .B(T4150_Y),     .A1(T4098_Y));
KC_AOI21_X1 T6536 ( .A0(T4178_Q), .Y(T6536_Y), .B(T13187_Y),     .A1(T13325_Y));
KC_AOI21_X1 T5713 ( .A0(T9564_Y), .Y(T5713_Y), .B(T12473_Y),     .A1(T15365_Y));
KC_AOI21_X1 T6742 ( .A0(T15907_Y), .Y(T6742_Y), .B(T5778_Y),     .A1(T5760_Y));
KC_AOI21_X1 T6027 ( .A0(T3790_Y), .Y(T6027_Y), .B(T5762_Y),     .A1(T4392_Y));
KC_AOI21_X1 T6114 ( .A0(T5830_Y), .Y(T6114_Y), .B(T11401_Y),     .A1(T4464_Y));
KC_AOI21_X1 T6099 ( .A0(T4435_Y), .Y(T6099_Y), .B(T11423_Y),     .A1(T3836_Y));
KC_AOI21_X1 T6089 ( .A0(T15908_Y), .Y(T6089_Y), .B(T4446_Y),     .A1(T145_Q));
KC_AOI21_X1 T6074 ( .A0(T4447_Y), .Y(T6074_Y), .B(T5799_Y),     .A1(T4447_Y));
KC_AOI21_X1 T6165 ( .A0(T4469_Y), .Y(T6165_Y), .B(T5142_Y),     .A1(T15572_Y));
KC_AOI21_X1 T6128 ( .A0(T14547_Q), .Y(T6128_Y), .B(T11433_Y),     .A1(T10922_Y));
KC_AOI21_X1 T6218 ( .A0(T89_Y), .Y(T6218_Y), .B(T2757_Y),     .A1(T4515_Y));
KC_AOI21_X1 T6217 ( .A0(T4534_Y), .Y(T6217_Y), .B(T4509_Y),     .A1(T5930_Y));
KC_AOI21_X1 T6173 ( .A0(T4542_Y), .Y(T6173_Y), .B(T8236_Y),     .A1(T3939_Y));
KC_AOI21_X1 T6284 ( .A0(T11587_Y), .Y(T6284_Y), .B(T11588_Y),     .A1(T16013_Y));
KC_AOI21_X1 T6261 ( .A0(T12221_Y), .Y(T6261_Y), .B(T2757_Y),     .A1(T12224_Y));
KC_AOI21_X1 T6242 ( .A0(T8272_Y), .Y(T6242_Y), .B(T2757_Y),     .A1(T12213_Y));
KC_AOI21_X1 T6327 ( .A0(T16020_Y), .Y(T6327_Y), .B(T6008_Y),     .A1(T3986_Y));
KC_AOI21_X1 T6326 ( .A0(T3973_Y), .Y(T6326_Y), .B(T12237_Y),     .A1(T3982_Y));
KC_AOI21_X1 T6467 ( .A0(T10614_Y), .Y(T6467_Y), .B(T11779_Y),     .A1(T8498_Y));
KC_AOI21_X1 T6448 ( .A0(T10598_Y), .Y(T6448_Y), .B(T11778_Y),     .A1(T8498_Y));
KC_AOI21_X1 T16315 ( .A0(T230_Y), .Y(T16315_Y), .B(T12608_Y),     .A1(T7697_Y));
KC_AOI21_X1 T6813 ( .A0(T12401_Y), .Y(T6813_Y), .B(T13245_Y),     .A1(T214_Y));
KC_AOI21_X1 T6812 ( .A0(T12398_Y), .Y(T6812_Y), .B(T13245_Y),     .A1(T214_Y));
KC_AOI21_X1 T6810 ( .A0(T15028_Y), .Y(T6810_Y), .B(T13245_Y),     .A1(T6805_Y));
KC_AOI21_X1 T269 ( .A0(T7108_Y), .Y(T269_Y), .B(T13248_Y),     .A1(T12398_Y));
KC_AOI21_X1 T16185 ( .A0(T1599_Y), .Y(T16185_Y), .B(T9476_Y),     .A1(T9243_Y));
KC_AOI21_X1 T15729 ( .A0(T6804_Y), .Y(T15729_Y), .B(T13244_Y),     .A1(T357_Y));
KC_AOI21_X1 T15728 ( .A0(T6804_Y), .Y(T15728_Y), .B(T13243_Y),     .A1(T10264_Y));
KC_AOI21_X1 T6807 ( .A0(T15028_Y), .Y(T6807_Y), .B(T13245_Y),     .A1(T12398_Y));
KC_AOI21_X1 T6341 ( .A0(T6804_Y), .Y(T6341_Y), .B(T721_Y),     .A1(T7318_Y));
KC_AOI21_X1 T6339 ( .A0(T7810_Y), .Y(T6339_Y), .B(T733_Y),     .A1(T6805_Y));
KC_AOI21_X1 T520 ( .A0(T7318_Y), .Y(T520_Y), .B(T721_Y),     .A1(T12398_Y));
KC_AOI21_X1 T6260 ( .A0(T6809_Y), .Y(T6260_Y), .B(T733_Y),     .A1(T12398_Y));
KC_AOI21_X1 T16380 ( .A0(T8792_Y), .Y(T16380_Y), .B(T8759_Y),     .A1(T7868_Y));
KC_AOI21_X1 T16379 ( .A0(T8792_Y), .Y(T16379_Y), .B(T8759_Y),     .A1(T763_Y));
KC_AOI21_X1 T15746 ( .A0(T7637_Y), .Y(T15746_Y), .B(T637_Y),     .A1(T919_Y));
KC_AOI21_X1 T15736 ( .A0(T6659_Y), .Y(T15736_Y), .B(T16425_Y),     .A1(T688_Q));
KC_AOI21_X1 T6253 ( .A0(T9334_Y), .Y(T6253_Y), .B(T16427_Y),     .A1(T7603_Y));
KC_AOI21_X1 T10808 ( .A0(T2564_Y), .Y(T10808_Y), .B(T6771_Y),     .A1(T5680_Y));
KC_AOI21_X1 T10807 ( .A0(T2564_Y), .Y(T10807_Y), .B(T15462_Y),     .A1(T5696_Y));
KC_AOI21_X1 T10758 ( .A0(T16164_Y), .Y(T10758_Y), .B(T15462_Y),     .A1(T3656_Y));
KC_AOI21_X1 T6816 ( .A0(T2311_Q), .Y(T6816_Y), .B(T13163_Y),     .A1(T6464_Y));
KC_AOI21_X1 T6766 ( .A0(T5486_Q), .Y(T6766_Y), .B(T13311_Y),     .A1(T12269_Y));
KC_AOI21_X1 T6845 ( .A0(T1_Y), .Y(T6845_Y), .B(T6844_Y),     .A1(T11038_Y));
KC_AOI21_X1 T6831 ( .A0(T6100_Y), .Y(T6831_Y), .B(T2860_Y),     .A1(T10554_Y));
KC_AOI21_X1 T6790 ( .A0(T2879_Y), .Y(T6790_Y), .B(T15974_Y),     .A1(T15606_Y));
KC_AOI21_X1 T6729 ( .A0(T15752_Y), .Y(T6729_Y), .B(T4994_Y),     .A1(T10280_Y));
KC_AOI21_X1 T6692 ( .A0(T10060_Y), .Y(T6692_Y), .B(T15502_Y),     .A1(T2037_Y));
KC_AOI21_X1 T6676 ( .A0(T9778_Y), .Y(T6676_Y), .B(T15442_Y),     .A1(T11947_Y));
KC_AOI21_X1 T6673 ( .A0(T14995_Y), .Y(T6673_Y), .B(T15532_Y),     .A1(T4250_Y));
KC_AOI21_X1 T6820 ( .A0(T4132_Y), .Y(T6820_Y), .B(T6119_Y),     .A1(T4091_Y));
KC_AOI21_X1 T6769 ( .A0(T10958_Y), .Y(T6769_Y), .B(T10937_Y),     .A1(T4595_Y));
KC_AOI21_X1 T6746 ( .A0(T11349_Y), .Y(T6746_Y), .B(T5842_Y),     .A1(T5838_Y));
KC_AOI21_X1 T6780 ( .A0(T2073_Y), .Y(T6780_Y), .B(T11588_Y),     .A1(T15969_Y));
KC_AOI21_X1 T6741 ( .A0(T5821_Y), .Y(T6741_Y), .B(T11972_Y),     .A1(T11347_Y));
KC_AOI21_X1 T6740 ( .A0(T145_Q), .Y(T6740_Y), .B(T5798_Y),     .A1(T3856_Y));
KC_AOI21_X1 T6226 ( .A0(T6804_Y), .Y(T6226_Y), .B(T16427_Y),     .A1(T6350_Y));
KC_AOI21_X1 T7102 ( .A0(T6804_Y), .Y(T7102_Y), .B(T735_Y),     .A1(T16162_Y));
KC_AOI21_X1 T7280 ( .A0(T6804_Y), .Y(T7280_Y), .B(T16426_Y),     .A1(T736_Y));
KC_AOI21_X1 T7261 ( .A0(T12398_Y), .Y(T7261_Y), .B(T16426_Y),     .A1(T16382_Y));
KC_AOI21_X1 T5810 ( .A0(T14995_Y), .Y(T5810_Y), .B(T15532_Y),     .A1(T3614_Y));
KC_AOI21_X1 T7970 ( .A0(T1586_Y), .Y(T7970_Y), .B(T16437_Y),     .A1(T10037_Y));
KC_AOI21_X1 T6340 ( .A0(T5122_Y), .Y(T6340_Y), .B(T3978_Y),     .A1(T6025_Y));
KC_AOI21_X1 T6520 ( .A0(T2958_Y), .Y(T6520_Y), .B(T11766_Y),     .A1(T2399_Y));
KC_AOI21_X1 T6824 ( .A0(T6585_Y), .Y(T6824_Y), .B(T12041_Y),     .A1(T3473_Y));
KC_AOI21_X1 T6682 ( .A0(T14995_Y), .Y(T6682_Y), .B(T875_Y),     .A1(T3669_Y));
KC_NAND4_X1 T5630 ( .D(T5627_Y), .C(T80_Y), .B(T5190_Q), .A(T5589_Q),     .Y(T5630_Y));
KC_NAND4_X1 T5636 ( .D(T9255_Y), .C(T5611_Y), .B(T55_Y), .A(T12457_Y),     .Y(T5636_Y));
KC_NAND4_X1 T5631 ( .D(T13294_Y), .C(T5628_Y), .B(T5184_Q),     .A(T5611_Y), .Y(T5631_Y));
KC_NAND4_X1 T5633 ( .D(T98_Q), .C(T101_Q), .B(T83_Q), .A(T5185_Q),     .Y(T5633_Y));
KC_NAND4_X1 T5623 ( .D(T101_Q), .C(T81_Q), .B(T8548_Y), .A(T15213_Y),     .Y(T5623_Y));
KC_NAND4_X1 T5606 ( .D(T15320_Y), .C(T5615_Y), .B(T105_Q), .A(T40_Y),     .Y(T5606_Y));
KC_NAND4_X1 T5616 ( .D(T8542_Y), .C(T14971_Y), .B(T69_Y), .A(T112_Y),     .Y(T5616_Y));
KC_NAND4_X1 T5615 ( .D(T14971_Y), .C(T16478_Y), .B(T7901_Y),     .A(T112_Y), .Y(T5615_Y));
KC_NAND4_X1 T5614 ( .D(T16479_Y), .C(T9270_Y), .B(T8545_Y),     .A(T8543_Y), .Y(T5614_Y));
KC_NAND4_X1 T5603 ( .D(T16479_Y), .C(T15316_Y), .B(T8545_Y),     .A(T5202_Q), .Y(T5603_Y));
KC_NAND4_X1 T5602 ( .D(T8558_Y), .C(T8559_Y), .B(T106_Q), .A(T5202_Q),     .Y(T5602_Y));
KC_NAND4_X1 T5601 ( .D(T12379_Y), .C(T8541_Y), .B(T5602_Y),     .A(T8561_Y), .Y(T5601_Y));
KC_NAND4_X1 T6321 ( .D(T6317_Y), .C(T6319_Y), .B(T6318_Y), .A(T5192_Q),     .Y(T6321_Y));
KC_NAND4_X1 T9291 ( .D(T6319_Y), .C(T6318_Y), .B(T5192_Q), .A(T131_Q),     .Y(T9291_Y));
KC_NAND4_X1 T9289 ( .D(T6319_Y), .C(T6317_Y), .B(T5192_Q), .A(T5225_Q),     .Y(T9289_Y));
KC_NAND4_X1 T9288 ( .D(T6319_Y), .C(T6318_Y), .B(T131_Q), .A(T8579_Y),     .Y(T9288_Y));
KC_NAND4_X1 T6971 ( .D(T8603_Y), .C(T15356_Y), .B(T137_Y), .A(T8600_Y),     .Y(T6971_Y));
KC_NAND4_X1 T6945 ( .D(T9286_Y), .C(T15356_Y), .B(T9269_Y),     .A(T8596_Y), .Y(T6945_Y));
KC_NAND4_X1 T6935 ( .D(T8582_Y), .C(T137_Y), .B(T9290_Y), .A(T12383_Y),     .Y(T6935_Y));
KC_NAND4_X1 T6932 ( .D(T257_Y), .C(T6318_Y), .B(T8580_Y), .A(T150_Q),     .Y(T6932_Y));
KC_NAND4_X1 T6913 ( .D(T6914_Y), .C(T9269_Y), .B(T8600_Y), .A(T8597_Y),     .Y(T6913_Y));
KC_NAND4_X1 T6912 ( .D(T8603_Y), .C(T9286_Y), .B(T6970_Y), .A(T8596_Y),     .Y(T6912_Y));
KC_NAND4_X1 T7697 ( .D(T647_Y), .C(T7580_Y), .B(T208_Q), .A(T4803_Q),     .Y(T7697_Y));
KC_NAND4_X1 T7583 ( .D(T802_Y), .C(T7580_Y), .B(T208_Q), .A(T207_Q),     .Y(T7583_Y));
KC_NAND4_X1 T9395 ( .D(T12383_Y), .C(T15656_Y), .B(T941_Y), .A(T878_Y),     .Y(T9395_Y));
KC_NAND4_X1 T9138 ( .D(T9133_Y), .C(T15100_Y), .B(T15150_Y),     .A(T4818_Y), .Y(T9138_Y));
KC_NAND4_X1 T9090 ( .D(T4800_Y), .C(T16286_Y), .B(T4817_Y),     .A(T9087_Y), .Y(T9090_Y));
KC_NAND4_X1 T9089 ( .D(T9071_Y), .C(T15100_Y), .B(T4818_Y),     .A(T15150_Y), .Y(T9089_Y));
KC_NAND4_X1 T9088 ( .D(T9117_Y), .C(T15100_Y), .B(T4818_Y),     .A(T15150_Y), .Y(T9088_Y));
KC_NAND4_X1 T9285 ( .D(T270_Y), .C(T6923_Y), .B(T6267_Y), .A(T6929_Y),     .Y(T9285_Y));
KC_NAND4_X1 T7069 ( .D(T5242_Q), .C(T289_Q), .B(T282_Q), .A(T281_Q),     .Y(T7069_Y));
KC_NAND4_X1 T7067 ( .D(T7062_Y), .C(T7061_Y), .B(T7066_Y), .A(T7064_Y),     .Y(T7067_Y));
KC_NAND4_X1 T9515 ( .D(T171_Q), .C(T316_Q), .B(T177_Q), .A(T330_Q),     .Y(T9515_Y));
KC_NAND4_X1 T7275 ( .D(T8627_Y), .C(T8574_Y), .B(T8647_Y), .A(T9516_Y),     .Y(T7275_Y));
KC_NAND4_X1 T7254 ( .D(T157_Q), .C(T180_Q), .B(T154_Q), .A(T179_Q),     .Y(T7254_Y));
KC_NAND4_X1 T9326 ( .D(T6715_Y), .C(T6721_Y), .B(T6717_Y), .A(T6615_Y),     .Y(T9326_Y));
KC_NAND4_X1 T9124 ( .D(T9129_Y), .C(T9077_Y), .B(T9128_Y), .A(T9127_Y),     .Y(T9124_Y));
KC_NAND4_X1 T9073 ( .D(T388_Y), .C(T11294_Y), .B(T16288_Y),     .A(T11295_Y), .Y(T9073_Y));
KC_NAND4_X1 T9281 ( .D(T442_Q), .C(T5200_Q), .B(T434_Q), .A(T438_Q),     .Y(T9281_Y));
KC_NAND4_X1 T9280 ( .D(T6921_Y), .C(T6309_Y), .B(T6312_Y), .A(T6925_Y),     .Y(T9280_Y));
KC_NAND4_X1 T7068 ( .D(T7057_Y), .C(T7063_Y), .B(T7065_Y), .A(T7118_Y),     .Y(T7068_Y));
KC_NAND4_X1 T7060 ( .D(T7058_Y), .C(T6263_Y), .B(T7054_Y), .A(T7081_Y),     .Y(T7060_Y));
KC_NAND4_X1 T9513 ( .D(T6617_Y), .C(T7304_Y), .B(T6642_Y), .A(T7659_Y),     .Y(T9513_Y));
KC_NAND4_X1 T9512 ( .D(T6644_Y), .C(T6616_Y), .B(T6640_Y), .A(T7657_Y),     .Y(T9512_Y));
KC_NAND4_X1 T7289 ( .D(T7273_Y), .C(T7271_Y), .B(T7269_Y), .A(T7285_Y),     .Y(T7289_Y));
KC_NAND4_X1 T7268 ( .D(T6643_Y), .C(T7283_Y), .B(T6639_Y), .A(T7655_Y),     .Y(T7268_Y));
KC_NAND4_X1 T9346 ( .D(T9354_Q), .C(T359_Q), .B(T9355_Q), .A(T9338_Q),     .Y(T9346_Y));
KC_NAND4_X1 T7452 ( .D(T7425_Y), .C(T6660_Y), .B(T7378_Y), .A(T7455_Y),     .Y(T7452_Y));
KC_NAND4_X1 T7429 ( .D(T7398_Y), .C(T7400_Y), .B(T7422_Y), .A(T7419_Y),     .Y(T7429_Y));
KC_NAND4_X1 T7421 ( .D(T8673_Y), .C(T189_Q), .B(T181_Q), .A(T341_Q),     .Y(T7421_Y));
KC_NAND4_X1 T7397 ( .D(T12882_Y), .C(T12574_Y), .B(T12496_Y),     .A(T12890_Y), .Y(T7397_Y));
KC_NAND4_X1 T7396 ( .D(T6711_Y), .C(T7394_Y), .B(T7395_Y), .A(T7648_Y),     .Y(T7396_Y));
KC_NAND4_X1 T7386 ( .D(T7379_Y), .C(T7380_Y), .B(T7376_Y), .A(T7373_Y),     .Y(T7386_Y));
KC_NAND4_X1 T7625 ( .D(T7620_Y), .C(T6666_Y), .B(T7602_Y), .A(T7656_Y),     .Y(T7625_Y));
KC_NAND4_X1 T7624 ( .D(T7622_Y), .C(T6665_Y), .B(T7619_Y), .A(T7654_Y),     .Y(T7624_Y));
KC_NAND4_X1 T7605 ( .D(T5303_Q), .C(T522_Q), .B(T363_Q), .A(T9339_Q),     .Y(T7605_Y));
KC_NAND4_X1 T7604 ( .D(T7621_Y), .C(T6667_Y), .B(T7600_Y), .A(T7649_Y),     .Y(T7604_Y));
KC_NAND4_X1 T7566 ( .D(T6414_Y), .C(T8749_Y), .B(T15768_Y),     .A(T8737_Y), .Y(T7566_Y));
KC_NAND4_X1 T7565 ( .D(T12605_Y), .C(T516_Y), .B(T7660_Y),     .A(T12441_Y), .Y(T7565_Y));
KC_NAND4_X1 T9418 ( .D(T11272_Y), .C(T8036_Y), .B(T7845_Y), .A(T960_Y),     .Y(T9418_Y));
KC_NAND4_X1 T8124 ( .D(T558_Y), .C(T8984_Y), .B(T9015_Y), .A(T11276_Y),     .Y(T8124_Y));
KC_NAND4_X1 T8061 ( .D(T1200_Y), .C(T8945_Y), .B(T8045_Y), .A(T8940_Y),     .Y(T8061_Y));
KC_NAND4_X1 T9097 ( .D(T9102_Y), .C(T9469_Q), .B(T604_Q), .A(T5587_Y),     .Y(T9097_Y));
KC_NAND4_X1 T9277 ( .D(T814_Q), .C(T624_Q), .B(T831_Q), .A(T627_Q),     .Y(T9277_Y));
KC_NAND4_X1 T9276 ( .D(T8583_Y), .C(T9279_Y), .B(T9273_Y), .A(T9256_Y),     .Y(T9276_Y));
KC_NAND4_X1 T9275 ( .D(T6281_Y), .C(T6276_Y), .B(T6285_Y), .A(T6275_Y),     .Y(T9275_Y));
KC_NAND4_X1 T6922 ( .D(T626_Q), .C(T443_Q), .B(T5198_Q), .A(T5196_Q),     .Y(T6922_Y));
KC_NAND4_X1 T7115 ( .D(T6259_Y), .C(T704_Y), .B(T7077_Y), .A(T1442_Y),     .Y(T7115_Y));
KC_NAND4_X1 T7112 ( .D(T7109_Y), .C(T6255_Y), .B(T7048_Y), .A(T7089_Y),     .Y(T7112_Y));
KC_NAND4_X1 T7093 ( .D(T12491_Y), .C(T12525_Y), .B(T12492_Y),     .A(T12493_Y), .Y(T7093_Y));
KC_NAND4_X1 T7056 ( .D(T7055_Y), .C(T6298_Y), .B(T7053_Y), .A(T7114_Y),     .Y(T7056_Y));
KC_NAND4_X1 T7051 ( .D(T12389_Y), .C(T6254_Y), .B(T7047_Y),     .A(T7076_Y), .Y(T7051_Y));
KC_NAND4_X1 T7050 ( .D(T7046_Y), .C(T7110_Y), .B(T7044_Y), .A(T6282_Y),     .Y(T7050_Y));
KC_NAND4_X1 T9509 ( .D(T6623_Y), .C(T6697_Y), .B(T6624_Y), .A(T6696_Y),     .Y(T9509_Y));
KC_NAND4_X1 T7299 ( .D(T7294_Y), .C(T6323_Y), .B(T7277_Y), .A(T7296_Y),     .Y(T7299_Y));
KC_NAND4_X1 T7241 ( .D(T7240_Y), .C(T6322_Y), .B(T7293_Y),     .A(T16512_Y), .Y(T7241_Y));
KC_NAND4_X1 T9337 ( .D(T6653_Y), .C(T6655_Y), .B(T6657_Y), .A(T7440_Y),     .Y(T9337_Y));
KC_NAND4_X1 T7443 ( .D(T7441_Y), .C(T7438_Y), .B(T7361_Y), .A(T7439_Y),     .Y(T7443_Y));
KC_NAND4_X1 T7417 ( .D(T9311_Y), .C(T8661_Y), .B(T3277_Y), .A(T6834_Y),     .Y(T7417_Y));
KC_NAND4_X1 T7416 ( .D(T12575_Y), .C(T6830_Y), .B(T7263_Y),     .A(T12494_Y), .Y(T7416_Y));
KC_NAND4_X1 T7393 ( .D(T6403_Y), .C(T6394_Y), .B(T6815_Y), .A(T6395_Y),     .Y(T7393_Y));
KC_NAND4_X1 T7366 ( .D(T691_Y), .C(T15047_Y), .B(T12402_Y),     .A(T12609_Y), .Y(T7366_Y));
KC_NAND4_X1 T7365 ( .D(T698_Q), .C(T688_Q), .B(T683_Q), .A(T7367_Q),     .Y(T7365_Y));
KC_NAND4_X1 T7643 ( .D(T11200_Y), .C(T11202_Y), .B(T6402_Y),     .A(T7642_Y), .Y(T7643_Y));
KC_NAND4_X1 T7598 ( .D(T5300_Q), .C(T705_Q), .B(T710_Q), .A(T687_Q),     .Y(T7598_Y));
KC_NAND4_X1 T9004 ( .D(T746_Y), .C(T9009_Y), .B(T1399_Y), .A(T8133_Y),     .Y(T9004_Y));
KC_NAND4_X1 T9003 ( .D(T8126_Y), .C(T1402_Y), .B(T8135_Y),     .A(T16280_Y), .Y(T9003_Y));
KC_NAND4_X1 T8115 ( .D(T8121_Y), .C(T1400_Y), .B(T8132_Y), .A(T753_Y),     .Y(T8115_Y));
KC_NAND4_X1 T8095 ( .D(T8129_Y), .C(T8114_Y), .B(T8096_Y), .A(T8113_Y),     .Y(T8095_Y));
KC_NAND4_X1 T8060 ( .D(T1349_Y), .C(T977_Q), .B(T8978_Y), .A(T5378_Q),     .Y(T8060_Y));
KC_NAND4_X1 T9098 ( .D(T9444_Y), .C(T16359_Y), .B(T1838_Y),     .A(T1676_Y), .Y(T9098_Y));
KC_NAND4_X1 T9095 ( .D(T9045_Y), .C(T12454_Y), .B(T1574_Y),     .A(T1653_Y), .Y(T9095_Y));
KC_NAND4_X1 T9049 ( .D(T9042_Y), .C(T7895_Y), .B(T1568_Y), .A(T1635_Y),     .Y(T9049_Y));
KC_NAND4_X1 T9040 ( .D(T9043_Y), .C(T16355_Y), .B(T1576_Y),     .A(T1566_Y), .Y(T9040_Y));
KC_NAND4_X1 T9038 ( .D(T9051_Y), .C(T1631_Y), .B(T7894_Y), .A(T1558_Y),     .Y(T9038_Y));
KC_NAND4_X1 T9037 ( .D(T9052_Y), .C(T1561_Y), .B(T8134_Y), .A(T1562_Y),     .Y(T9037_Y));
KC_NAND4_X1 T9036 ( .D(T9044_Y), .C(T8033_Y), .B(T1575_Y), .A(T1666_Y),     .Y(T9036_Y));
KC_NAND4_X1 T9035 ( .D(T9041_Y), .C(T16357_Y), .B(T1741_Y),     .A(T1636_Y), .Y(T9035_Y));
KC_NAND4_X1 T9226 ( .D(T9462_Y), .C(T777_Y), .B(T778_Y), .A(T9240_Y),     .Y(T9226_Y));
KC_NAND4_X1 T7052 ( .D(T816_Q), .C(T793_Q), .B(T813_Q), .A(T5199_Q),     .Y(T7052_Y));
KC_NAND4_X1 T7300 ( .D(T4855_Q), .C(T670_Q), .B(T676_Q), .A(T679_Q),     .Y(T7300_Y));
KC_NAND4_X1 T7597 ( .D(T8396_Y), .C(T11194_Y), .B(T6382_Y),     .A(T7596_Y), .Y(T7597_Y));
KC_NAND4_X1 T7589 ( .D(T11189_Y), .C(T11878_Y), .B(T15738_Y),     .A(T15736_Y), .Y(T7589_Y));
KC_NAND4_X1 T7562 ( .D(T16115_Y), .C(T11178_Y), .B(T6381_Y),     .A(T7641_Y), .Y(T7562_Y));
KC_NAND4_X1 T9403 ( .D(T937_Y), .C(T9404_Y), .B(T7840_Y), .A(T9400_Y),     .Y(T9403_Y));
KC_NAND4_X1 T9402 ( .D(T15457_Y), .C(T992_Q), .B(T925_Y), .A(T938_Q),     .Y(T9402_Y));
KC_NAND4_X1 T9401 ( .D(T979_Y), .C(T7876_Y), .B(T9400_Y), .A(T8847_Y),     .Y(T9401_Y));
KC_NAND4_X1 T9400 ( .D(T948_Y), .C(T981_Q), .B(T992_Q), .A(T925_Y),     .Y(T9400_Y));
KC_NAND4_X1 T7880 ( .D(T8800_Y), .C(T7877_Y), .B(T7878_Y), .A(T7839_Y),     .Y(T7880_Y));
KC_NAND4_X1 T7879 ( .D(T9405_Y), .C(T979_Y), .B(T7877_Y), .A(T16383_Y),     .Y(T7879_Y));
KC_NAND4_X1 T7878 ( .D(T8846_Y), .C(T938_Q), .B(T8795_Y), .A(T940_Q),     .Y(T7878_Y));
KC_NAND4_X1 T7877 ( .D(T947_Y), .C(T8848_Y), .B(T8846_Y), .A(T938_Q),     .Y(T7877_Y));
KC_NAND4_X1 T7876 ( .D(T948_Y), .C(T947_Y), .B(T8845_Y), .A(T8796_Y),     .Y(T7876_Y));
KC_NAND4_X1 T7839 ( .D(T947_Y), .C(T8796_Y), .B(T8846_Y), .A(T938_Q),     .Y(T7839_Y));
KC_NAND4_X1 T9005 ( .D(T8131_Y), .C(T1405_Y), .B(T8122_Y), .A(T1415_Y),     .Y(T9005_Y));
KC_NAND4_X1 T8998 ( .D(T8999_Y), .C(T9006_Y), .B(T1391_Y), .A(T8982_Y),     .Y(T8998_Y));
KC_NAND4_X1 T9039 ( .D(T9050_Y), .C(T1565_Y), .B(T1425_Y), .A(T1550_Y),     .Y(T9039_Y));
KC_NAND4_X1 T9223 ( .D(T9219_Y), .C(T9221_Y), .B(T9220_Y),     .A(T10220_Y), .Y(T9223_Y));
KC_NAND4_X1 T10391 ( .D(T9562_Y), .C(T7029_Y), .B(T7032_Y),     .A(T10863_Y), .Y(T10391_Y));
KC_NAND4_X1 T7036 ( .D(T9555_Y), .C(T7003_Y), .B(T7033_Y),     .A(T10861_Y), .Y(T7036_Y));
KC_NAND4_X1 T7035 ( .D(T10645_Y), .C(T7031_Y), .B(T7030_Y),     .A(T10862_Y), .Y(T7035_Y));
KC_NAND4_X1 T7034 ( .D(T9558_Y), .C(T7028_Y), .B(T7021_Y),     .A(T10860_Y), .Y(T7034_Y));
KC_NAND4_X1 T7236 ( .D(T10646_Y), .C(T7237_Y), .B(T7161_Y),     .A(T10864_Y), .Y(T7236_Y));
KC_NAND4_X1 T7235 ( .D(T9560_Y), .C(T7164_Y), .B(T7229_Y),     .A(T10865_Y), .Y(T7235_Y));
KC_NAND4_X1 T7234 ( .D(T9538_Y), .C(T7163_Y), .B(T7230_Y),     .A(T10859_Y), .Y(T7234_Y));
KC_NAND4_X1 T7233 ( .D(T9559_Y), .C(T7203_Y), .B(T7162_Y),     .A(T10648_Y), .Y(T7233_Y));
KC_NAND4_X1 T7232 ( .D(T9554_Y), .C(T7204_Y), .B(T7166_Y),     .A(T10869_Y), .Y(T7232_Y));
KC_NAND4_X1 T7231 ( .D(T10644_Y), .C(T7168_Y), .B(T7167_Y),     .A(T10858_Y), .Y(T7231_Y));
KC_NAND4_X1 T7207 ( .D(T9561_Y), .C(T7205_Y), .B(T7165_Y), .A(T7228_Y),     .Y(T7207_Y));
KC_NAND4_X1 T7206 ( .D(T9553_Y), .C(T10879_Y), .B(T7202_Y),     .A(T10868_Y), .Y(T7206_Y));
KC_NAND4_X1 T10343 ( .D(T11917_Y), .C(T11165_Y), .B(T15741_Y),     .A(T7436_Y), .Y(T10343_Y));
KC_NAND4_X1 T7550 ( .D(T11170_Y), .C(T12079_Y), .B(T6646_Y),     .A(T899_Y), .Y(T7550_Y));
KC_NAND4_X1 T7499 ( .D(T515_Y), .C(T11880_Y), .B(T11918_Y),     .A(T8724_Y), .Y(T7499_Y));
KC_NAND4_X1 T7359 ( .D(T11138_Y), .C(T11142_Y), .B(T6380_Y),     .A(T7358_Y), .Y(T7359_Y));
KC_NAND4_X1 T7613 ( .D(T1052_Y), .C(T12432_Y), .B(T12430_Y),     .A(T12419_Y), .Y(T7613_Y));
KC_NAND4_X1 T7556 ( .D(T636_Y), .C(T15433_Y), .B(T8684_Y), .A(T8726_Y),     .Y(T7556_Y));
KC_NAND4_X1 T7951 ( .D(T1008_Y), .C(T16394_Y), .B(T1009_Y), .A(T987_Y),     .Y(T7951_Y));
KC_NAND4_X1 T10028 ( .D(T927_Y), .C(T980_Q), .B(T1469_Y), .A(T10049_Y),     .Y(T10028_Y));
KC_NAND4_X1 T10170 ( .D(T16414_Y), .C(T1457_Y), .B(T15497_Y),     .A(T16308_Y), .Y(T10170_Y));
KC_NAND4_X1 T1164 ( .D(T10235_Y), .C(T10222_Y), .B(T9185_Y),     .A(T10221_Y), .Y(T1164_Y));
KC_NAND4_X1 T1165 ( .D(T10236_Y), .C(T10237_Y), .B(T10234_Y),     .A(T13060_Y), .Y(T1165_Y));
KC_NAND4_X1 T1166 ( .D(T10215_Y), .C(T10212_Y), .B(T10230_Y),     .A(T10219_Y), .Y(T1166_Y));
KC_NAND4_X1 T7027 ( .D(T9535_Y), .C(T7023_Y), .B(T7002_Y),     .A(T10856_Y), .Y(T7027_Y));
KC_NAND4_X1 T7026 ( .D(T10382_Y), .C(T7018_Y), .B(T7022_Y),     .A(T10854_Y), .Y(T7026_Y));
KC_NAND4_X1 T7025 ( .D(T9556_Y), .C(T7024_Y), .B(T7019_Y),     .A(T10855_Y), .Y(T7025_Y));
KC_NAND4_X1 T6984 ( .D(T9549_Y), .C(T7020_Y), .B(T7001_Y),     .A(T10857_Y), .Y(T6984_Y));
KC_NAND4_X1 T7227 ( .D(T9552_Y), .C(T7223_Y), .B(T7152_Y), .A(T7146_Y),     .Y(T7227_Y));
KC_NAND4_X1 T7201 ( .D(T9557_Y), .C(T7156_Y), .B(T7198_Y), .A(T7196_Y),     .Y(T7201_Y));
KC_NAND4_X1 T7200 ( .D(T9534_Y), .C(T7224_Y), .B(T7199_Y), .A(T7197_Y),     .Y(T7200_Y));
KC_NAND4_X1 T7160 ( .D(T9547_Y), .C(T7225_Y), .B(T7153_Y), .A(T7147_Y),     .Y(T7160_Y));
KC_NAND4_X1 T7159 ( .D(T10383_Y), .C(T7154_Y), .B(T7155_Y),     .A(T7149_Y), .Y(T7159_Y));
KC_NAND4_X1 T7158 ( .D(T9537_Y), .C(T7226_Y), .B(T7157_Y), .A(T7195_Y),     .Y(T7158_Y));
KC_NAND4_X1 T7150 ( .D(T9548_Y), .C(T7222_Y), .B(T7145_Y), .A(T7148_Y),     .Y(T7150_Y));
KC_NAND4_X1 T5701 ( .D(T9628_Y), .C(T10832_Y), .B(T5689_Y),     .A(T10827_Y), .Y(T5701_Y));
KC_NAND4_X1 T5696 ( .D(T9627_Y), .C(T10830_Y), .B(T5687_Y),     .A(T5685_Y), .Y(T5696_Y));
KC_NAND4_X1 T5695 ( .D(T9616_Y), .C(T5700_Y), .B(T5683_Y), .A(T5692_Y),     .Y(T5695_Y));
KC_NAND4_X1 T5694 ( .D(T10429_Y), .C(T10831_Y), .B(T7342_Y),     .A(T5684_Y), .Y(T5694_Y));
KC_NAND4_X1 T5693 ( .D(T9626_Y), .C(T5699_Y), .B(T5686_Y), .A(T5690_Y),     .Y(T5693_Y));
KC_NAND4_X1 T5681 ( .D(T9615_Y), .C(T10814_Y), .B(T5688_Y),     .A(T7512_Y), .Y(T5681_Y));
KC_NAND4_X1 T5678 ( .D(T9625_Y), .C(T5691_Y), .B(T7341_Y), .A(T7513_Y),     .Y(T5678_Y));
KC_NAND4_X1 T7548 ( .D(T9703_Y), .C(T7470_Y), .B(T7494_Y), .A(T7543_Y),     .Y(T7548_Y));
KC_NAND4_X1 T7547 ( .D(T9722_Y), .C(T7471_Y), .B(T7495_Y), .A(T7546_Y),     .Y(T7547_Y));
KC_NAND4_X1 T7518 ( .D(T9701_Y), .C(T7520_Y), .B(T10824_Y),     .A(T7517_Y), .Y(T7518_Y));
KC_NAND4_X1 T7496 ( .D(T9702_Y), .C(T7519_Y), .B(T10825_Y),     .A(T7493_Y), .Y(T7496_Y));
KC_NAND4_X1 T7472 ( .D(T10341_Y), .C(T7469_Y), .B(T10791_Y),     .A(T7773_Y), .Y(T7472_Y));
KC_NAND4_X1 T7777 ( .D(T10342_Y), .C(T7734_Y), .B(T7770_Y),     .A(T7766_Y), .Y(T7777_Y));
KC_NAND4_X1 T7776 ( .D(T10340_Y), .C(T7468_Y), .B(T7771_Y),     .A(T7765_Y), .Y(T7776_Y));
KC_NAND4_X1 T7775 ( .D(T9807_Y), .C(T7769_Y), .B(T7772_Y), .A(T7774_Y),     .Y(T7775_Y));
KC_NAND4_X1 T7739 ( .D(T9805_Y), .C(T7736_Y), .B(T10790_Y),     .A(T7737_Y), .Y(T7739_Y));
KC_NAND4_X1 T7738 ( .D(T9806_Y), .C(T7718_Y), .B(T7735_Y), .A(T7728_Y),     .Y(T7738_Y));
KC_NAND4_X1 T10314 ( .D(T1224_Q), .C(T1195_Q), .B(T1221_Q),     .A(T1231_Q), .Y(T10314_Y));
KC_NAND4_X1 T8024 ( .D(T1202_Q), .C(T4869_Q), .B(T1188_Q), .A(T1209_Q),     .Y(T8024_Y));
KC_NAND4_X1 T8023 ( .D(T1203_Q), .C(T1215_Q), .B(T1216_Q), .A(T1190_Q),     .Y(T8023_Y));
KC_NAND4_X1 T10041 ( .D(T1193_Y), .C(T5370_Y), .B(T1218_Y),     .A(T16126_Y), .Y(T10041_Y));
KC_NAND4_X1 T10025 ( .D(T1238_Y), .C(T5372_Y), .B(T1239_Y),     .A(T1237_Y), .Y(T10025_Y));
KC_NAND4_X1 T9986 ( .D(T16276_Y), .C(T10163_Y), .B(T1365_Y),     .A(T10293_Y), .Y(T9986_Y));
KC_NAND4_X1 T10171 ( .D(T10154_Y), .C(T10298_Y), .B(T4868_Y),     .A(T10157_Y), .Y(T10171_Y));
KC_NAND4_X1 T10169 ( .D(T2103_Y), .C(T9984_Y), .B(T10141_Y),     .A(T15817_Y), .Y(T10169_Y));
KC_NAND4_X1 T10158 ( .D(T4902_Y), .C(T1365_Y), .B(T10139_Y),     .A(T15529_Y), .Y(T10158_Y));
KC_NAND4_X1 T1277 ( .D(T10209_Y), .C(T10287_Y), .B(T10213_Y),     .A(T10124_Y), .Y(T1277_Y));
KC_NAND4_X1 T10390 ( .D(T9536_Y), .C(T10851_Y), .B(T7000_Y),     .A(T10853_Y), .Y(T10390_Y));
KC_NAND4_X1 T7017 ( .D(T9551_Y), .C(T7013_Y), .B(T6998_Y),     .A(T10852_Y), .Y(T7017_Y));
KC_NAND4_X1 T7016 ( .D(T9544_Y), .C(T7014_Y), .B(T6999_Y), .A(T7008_Y),     .Y(T7016_Y));
KC_NAND4_X1 T7011 ( .D(T9533_Y), .C(T7015_Y), .B(T6996_Y),     .A(T10850_Y), .Y(T7011_Y));
KC_NAND4_X1 T7010 ( .D(T9545_Y), .C(T7012_Y), .B(T6994_Y), .A(T7009_Y),     .Y(T7010_Y));
KC_NAND4_X1 T6997 ( .D(T10381_Y), .C(T7007_Y), .B(T6995_Y),     .A(T10849_Y), .Y(T6997_Y));
KC_NAND4_X1 T7219 ( .D(T9546_Y), .C(T7213_Y), .B(T7211_Y), .A(T7214_Y),     .Y(T7219_Y));
KC_NAND4_X1 T7218 ( .D(T9532_Y), .C(T7221_Y), .B(T7216_Y), .A(T7212_Y),     .Y(T7218_Y));
KC_NAND4_X1 T7151 ( .D(T9550_Y), .C(T7220_Y), .B(T7144_Y),     .A(T10647_Y), .Y(T7151_Y));
KC_NAND4_X1 T5680 ( .D(T9621_Y), .C(T10820_Y), .B(T10811_Y),     .A(T7511_Y), .Y(T5680_Y));
KC_NAND4_X1 T10370 ( .D(T9619_Y), .C(T10823_Y), .B(T6792_Y),     .A(T7515_Y), .Y(T10370_Y));
KC_NAND4_X1 T10369 ( .D(T9620_Y), .C(T10821_Y), .B(T10810_Y),     .A(T7510_Y), .Y(T10369_Y));
KC_NAND4_X1 T7467 ( .D(T10339_Y), .C(T7465_Y), .B(T7491_Y),     .A(T7544_Y), .Y(T7467_Y));
KC_NAND4_X1 T9790 ( .D(T9804_Y), .C(T7712_Y), .B(T7715_Y), .A(T7795_Y),     .Y(T9790_Y));
KC_NAND4_X1 T7757 ( .D(T9800_Y), .C(T7722_Y), .B(T7723_Y), .A(T7710_Y),     .Y(T7757_Y));
KC_NAND4_X1 T7733 ( .D(T9799_Y), .C(T7730_Y), .B(T7729_Y), .A(T7794_Y),     .Y(T7733_Y));
KC_NAND4_X1 T7732 ( .D(T9802_Y), .C(T7731_Y), .B(T7727_Y), .A(T7716_Y),     .Y(T7732_Y));
KC_NAND4_X1 T7717 ( .D(T9798_Y), .C(T7714_Y), .B(T7713_Y), .A(T7796_Y),     .Y(T7717_Y));
KC_NAND4_X1 T7711 ( .D(T9801_Y), .C(T7709_Y), .B(T7724_Y), .A(T7791_Y),     .Y(T7711_Y));
KC_NAND4_X1 T8022 ( .D(T9908_Y), .C(T8018_Y), .B(T8020_Y), .A(T8016_Y),     .Y(T8022_Y));
KC_NAND4_X1 T7996 ( .D(T9887_Y), .C(T7988_Y), .B(T7995_Y), .A(T7969_Y),     .Y(T7996_Y));
KC_NAND4_X1 T7991 ( .D(T10292_Y), .C(T8021_Y), .B(T7994_Y),     .A(T7965_Y), .Y(T7991_Y));
KC_NAND4_X1 T7990 ( .D(T9885_Y), .C(T7973_Y), .B(T7993_Y), .A(T7966_Y),     .Y(T7990_Y));
KC_NAND4_X1 T7989 ( .D(T10290_Y), .C(T7974_Y), .B(T7992_Y),     .A(T7964_Y), .Y(T7989_Y));
KC_NAND4_X1 T7975 ( .D(T9909_Y), .C(T8019_Y), .B(T7972_Y), .A(T7968_Y),     .Y(T7975_Y));
KC_NAND4_X1 T7948 ( .D(T1212_Q), .C(T1211_Q), .B(T1207_Q), .A(T1208_Q),     .Y(T7948_Y));
KC_NAND4_X1 T7943 ( .D(T9886_Y), .C(T7937_Y), .B(T10754_Y),     .A(T7938_Y), .Y(T7943_Y));
KC_NAND4_X1 T7942 ( .D(T10312_Y), .C(T7936_Y), .B(T10721_Y),     .A(T7941_Y), .Y(T7942_Y));
KC_NAND4_X1 T10038 ( .D(T10036_Y), .C(T10720_Y), .B(T10691_Y),     .A(T10718_Y), .Y(T10038_Y));
KC_NAND4_X1 T10037 ( .D(T10019_Y), .C(T10719_Y), .B(T10696_Y),     .A(T10717_Y), .Y(T10037_Y));
KC_NAND4_X1 T9999 ( .D(T9979_Y), .C(T10671_Y), .B(T10682_Y),     .A(T10694_Y), .Y(T9999_Y));
KC_NAND4_X1 T9997 ( .D(T9978_Y), .C(T10672_Y), .B(T10675_Y),     .A(T10681_Y), .Y(T9997_Y));
KC_NAND4_X1 T9996 ( .D(T10291_Y), .C(T10673_Y), .B(T10674_Y),     .A(T10690_Y), .Y(T9996_Y));
KC_NAND4_X1 T9980 ( .D(T10151_Y), .C(T10656_Y), .B(T10658_Y),     .A(T10693_Y), .Y(T9980_Y));
KC_NAND4_X1 T1358 ( .D(T10725_Y), .C(T1368_Y), .B(T1372_Y),     .A(T4819_Y), .Y(T1358_Y));
KC_NAND4_X1 T5662 ( .D(T10357_Y), .C(T5656_Y), .B(T5665_Y),     .A(T5653_Y), .Y(T5662_Y));
KC_NAND4_X1 T10363 ( .D(T9708_Y), .C(T10804_Y), .B(T5655_Y),     .A(T5658_Y), .Y(T10363_Y));
KC_NAND4_X1 T7945 ( .D(T10311_Y), .C(T7987_Y), .B(T1480_Y),     .A(T7939_Y), .Y(T7945_Y));
KC_NAND4_X1 T7944 ( .D(T9884_Y), .C(T7929_Y), .B(T10752_Y),     .A(T7940_Y), .Y(T7944_Y));
KC_NAND4_X1 T7935 ( .D(T10148_Y), .C(T7930_Y), .B(T10705_Y),     .A(T10749_Y), .Y(T7935_Y));
KC_NAND4_X1 T7934 ( .D(T10150_Y), .C(T7931_Y), .B(T10714_Y),     .A(T10750_Y), .Y(T7934_Y));
KC_NAND4_X1 T10035 ( .D(T10149_Y), .C(T7933_Y), .B(T10715_Y),     .A(T10713_Y), .Y(T10035_Y));
KC_NAND4_X1 T10034 ( .D(T10134_Y), .C(T7932_Y), .B(T10706_Y),     .A(T10748_Y), .Y(T10034_Y));
KC_NAND4_X1 T7039 ( .D(T10375_Y), .C(T6988_Y), .B(T10836_Y),     .A(T6977_Y), .Y(T7039_Y));
KC_NAND4_X1 T5661 ( .D(T9710_Y), .C(T10803_Y), .B(T5652_Y),     .A(T5654_Y), .Y(T5661_Y));
KC_NAND4_X1 T10364 ( .D(T9711_Y), .C(T7506_Y), .B(T10806_Y),     .A(T5660_Y), .Y(T10364_Y));
KC_NAND4_X1 T10353 ( .D(T9715_Y), .C(T7500_Y), .B(T10800_Y),     .A(T10796_Y), .Y(T10353_Y));
KC_NAND4_X1 T10335 ( .D(T10332_Y), .C(T10775_Y), .B(T10773_Y),     .A(T10774_Y), .Y(T10335_Y));
KC_NAND4_X1 T10334 ( .D(T9796_Y), .C(T10772_Y), .B(T10778_Y),     .A(T10780_Y), .Y(T10334_Y));
KC_NAND4_X1 T7533 ( .D(T9717_Y), .C(T7485_Y), .B(T7484_Y), .A(T7527_Y),     .Y(T7533_Y));
KC_NAND4_X1 T7507 ( .D(T9697_Y), .C(T7505_Y), .B(T10805_Y),     .A(T5659_Y), .Y(T7507_Y));
KC_NAND4_X1 T7504 ( .D(T9716_Y), .C(T7501_Y), .B(T10798_Y),     .A(T10797_Y), .Y(T7504_Y));
KC_NAND4_X1 T7463 ( .D(T9718_Y), .C(T7483_Y), .B(T7486_Y), .A(T7530_Y),     .Y(T7463_Y));
KC_NAND4_X1 T7754 ( .D(T9794_Y), .C(T10776_Y), .B(T7744_Y),     .A(T7742_Y), .Y(T7754_Y));
KC_NAND4_X1 T7753 ( .D(T9797_Y), .C(T7749_Y), .B(T7746_Y), .A(T7752_Y),     .Y(T7753_Y));
KC_NAND4_X1 T7721 ( .D(T9791_Y), .C(T10782_Y), .B(T7745_Y),     .A(T7747_Y), .Y(T7721_Y));
KC_NAND4_X1 T10310 ( .D(T10133_Y), .C(T7926_Y), .B(T10704_Y),     .A(T10744_Y), .Y(T10310_Y));
KC_NAND4_X1 T10307 ( .D(T10145_Y), .C(T10710_Y), .B(T10703_Y),     .A(T10699_Y), .Y(T10307_Y));
KC_NAND4_X1 T7928 ( .D(T10146_Y), .C(T7927_Y), .B(T10707_Y),     .A(T10746_Y), .Y(T7928_Y));
KC_NAND4_X1 T10012 ( .D(T10126_Y), .C(T10667_Y), .B(T10685_Y),     .A(T10679_Y), .Y(T10012_Y));
KC_NAND4_X1 T10011 ( .D(T10147_Y), .C(T10745_Y), .B(T10708_Y),     .A(T10709_Y), .Y(T10011_Y));
KC_NAND4_X1 T10010 ( .D(T10121_Y), .C(T10686_Y), .B(T10684_Y),     .A(T10687_Y), .Y(T10010_Y));
KC_NAND4_X1 T9994 ( .D(T10125_Y), .C(T10670_Y), .B(T10653_Y),     .A(T10680_Y), .Y(T9994_Y));
KC_NAND4_X1 T9993 ( .D(T10135_Y), .C(T10666_Y), .B(T10688_Y),     .A(T10665_Y), .Y(T9993_Y));
KC_NAND4_X1 T9992 ( .D(T10289_Y), .C(T10654_Y), .B(T10662_Y),     .A(T10678_Y), .Y(T9992_Y));
KC_NAND4_X1 T9991 ( .D(T10728_Y), .C(T10711_Y), .B(T10677_Y),     .A(T10683_Y), .Y(T9991_Y));
KC_NAND4_X1 T9989 ( .D(T10288_Y), .C(T10655_Y), .B(T10663_Y),     .A(T10676_Y), .Y(T9989_Y));
KC_NAND4_X1 T10387 ( .D(T10384_Y), .C(T7004_Y), .B(T10847_Y),     .A(T1619_Y), .Y(T10387_Y));
KC_NAND4_X1 T10386 ( .D(T10385_Y), .C(T7005_Y), .B(T7006_Y),     .A(T4910_Y), .Y(T10386_Y));
KC_NAND4_X1 T7038 ( .D(T9521_Y), .C(T6978_Y), .B(T1623_Y), .A(T1624_Y),     .Y(T7038_Y));
KC_NAND4_X1 T6989 ( .D(T10376_Y), .C(T6985_Y), .B(T7037_Y),     .A(T6986_Y), .Y(T6989_Y));
KC_NAND4_X1 T6981 ( .D(T10377_Y), .C(T6974_Y), .B(T6976_Y),     .A(T6973_Y), .Y(T6981_Y));
KC_NAND4_X1 T6980 ( .D(T10378_Y), .C(T6975_Y), .B(T6972_Y),     .A(T6979_Y), .Y(T6980_Y));
KC_NAND4_X1 T1620 ( .D(T9519_Y), .C(T6987_Y), .B(T5718_Y), .A(T5720_Y),     .Y(T1620_Y));
KC_NAND4_X1 T1621 ( .D(T9517_Y), .C(T5211_Y), .B(T5207_Y), .A(T1884_Y),     .Y(T1621_Y));
KC_NAND4_X1 T1622 ( .D(T9518_Y), .C(T5726_Y), .B(T1872_Y), .A(T5719_Y),     .Y(T1622_Y));
KC_NAND4_X1 T7185 ( .D(T9583_Y), .C(T7209_Y), .B(T7124_Y), .A(T7125_Y),     .Y(T7185_Y));
KC_NAND4_X1 T7126 ( .D(T9584_Y), .C(T7210_Y), .B(T7123_Y), .A(T1625_Y),     .Y(T7126_Y));
KC_NAND4_X1 T1627 ( .D(T10392_Y), .C(T5233_Y), .B(T1626_Y),     .A(T1630_Y), .Y(T1627_Y));
KC_NAND4_X1 T1628 ( .D(T10393_Y), .C(T1928_Y), .B(T5232_Y),     .A(T1629_Y), .Y(T1628_Y));
KC_NAND4_X1 T7347 ( .D(T9629_Y), .C(T7174_Y), .B(T7344_Y), .A(T7319_Y),     .Y(T7347_Y));
KC_NAND4_X1 T7346 ( .D(T9630_Y), .C(T7171_Y), .B(T7345_Y),     .A(T10876_Y), .Y(T7346_Y));
KC_NAND4_X1 T10352 ( .D(T9689_Y), .C(T7476_Y), .B(T10799_Y),     .A(T4909_Y), .Y(T10352_Y));
KC_NAND4_X1 T7528 ( .D(T9691_Y), .C(T7522_Y), .B(T7475_Y), .A(T1642_Y),     .Y(T7528_Y));
KC_NAND4_X1 T7482 ( .D(T9695_Y), .C(T7480_Y), .B(T10650_Y),     .A(T7474_Y), .Y(T7482_Y));
KC_NAND4_X1 T7481 ( .D(T9690_Y), .C(T7525_Y), .B(T7479_Y), .A(T1643_Y),     .Y(T7481_Y));
KC_NAND4_X1 T1640 ( .D(T9694_Y), .C(T7478_Y), .B(T7502_Y), .A(T1644_Y),     .Y(T1640_Y));
KC_NAND4_X1 T1645 ( .D(T9750_Y), .C(T7477_Y), .B(T7503_Y), .A(T1646_Y),     .Y(T1645_Y));
KC_NAND4_X1 T1647 ( .D(T9693_Y), .C(T7526_Y), .B(T7523_Y), .A(T5808_Y),     .Y(T1647_Y));
KC_NAND4_X1 T1648 ( .D(T9692_Y), .C(T7461_Y), .B(T1641_Y), .A(T1649_Y),     .Y(T1648_Y));
KC_NAND4_X1 T9990 ( .D(T10132_Y), .C(T10668_Y), .B(T10664_Y),     .A(T10669_Y), .Y(T9990_Y));
KC_NAND4_X1 T1720 ( .D(T3786_Y), .C(T3898_Y), .B(T10063_Y),     .A(T10066_Y), .Y(T1720_Y));
KC_NAND4_X1 T1721 ( .D(T10067_Y), .C(T10532_Y), .B(T9976_Y),     .A(T10068_Y), .Y(T1721_Y));
KC_NAND4_X1 T1744 ( .D(T1748_Y), .C(T15856_Y), .B(T15854_Y),     .A(T15853_Y), .Y(T1744_Y));
KC_NAND4_X1 T1771 ( .D(T2240_Y), .C(T5927_Y), .B(T16041_Y),     .A(T15611_Y), .Y(T1771_Y));
KC_NAND4_X1 T1780 ( .D(T2247_Y), .C(T1786_Y), .B(T1788_Y), .A(T6028_Y),     .Y(T1780_Y));
KC_NAND4_X1 T1781 ( .D(T2245_Y), .C(T16042_Y), .B(T2280_Y),     .A(T16017_Y), .Y(T1781_Y));
KC_NAND4_X1 T1783 ( .D(T1793_Y), .C(T1782_Y), .B(T2271_Y), .A(T4914_Y),     .Y(T1783_Y));
KC_NAND4_X1 T1792 ( .D(T1791_Y), .C(T1797_Y), .B(T2284_Y), .A(T1795_Y),     .Y(T1792_Y));
KC_NAND4_X1 T1815 ( .D(T1814_Y), .C(T1810_Y), .B(T2299_Y), .A(T4913_Y),     .Y(T1815_Y));
KC_NAND4_X1 T1816 ( .D(T1813_Y), .C(T1818_Y), .B(T2300_Y), .A(T1809_Y),     .Y(T1816_Y));
KC_NAND4_X1 T1873 ( .D(T9531_Y), .C(T1882_Y), .B(T1898_Y), .A(T1894_Y),     .Y(T1873_Y));
KC_NAND4_X1 T1874 ( .D(T9530_Y), .C(T1880_Y), .B(T1895_Y), .A(T2424_Y),     .Y(T1874_Y));
KC_NAND4_X1 T1875 ( .D(T9520_Y), .C(T1876_Y), .B(T1883_Y), .A(T1893_Y),     .Y(T1875_Y));
KC_NAND4_X1 T1885 ( .D(T10463_Y), .C(T1877_Y), .B(T1896_Y),     .A(T1888_Y), .Y(T1885_Y));
KC_NAND4_X1 T1886 ( .D(T10464_Y), .C(T1890_Y), .B(T1897_Y),     .A(T1889_Y), .Y(T1886_Y));
KC_NAND4_X1 T1892 ( .D(T10379_Y), .C(T1891_Y), .B(T1878_Y),     .A(T1887_Y), .Y(T1892_Y));
KC_NAND4_X1 T1899 ( .D(T9595_Y), .C(T1926_Y), .B(T1905_Y), .A(T1907_Y),     .Y(T1899_Y));
KC_NAND4_X1 T1913 ( .D(T9597_Y), .C(T1923_Y), .B(T1915_Y), .A(T1902_Y),     .Y(T1913_Y));
KC_NAND4_X1 T1914 ( .D(T9596_Y), .C(T1925_Y), .B(T1901_Y), .A(T1900_Y),     .Y(T1914_Y));
KC_NAND4_X1 T1916 ( .D(T9594_Y), .C(T1927_Y), .B(T1906_Y), .A(T1919_Y),     .Y(T1916_Y));
KC_NAND4_X1 T1917 ( .D(T9598_Y), .C(T1922_Y), .B(T1903_Y), .A(T1920_Y),     .Y(T1917_Y));
KC_NAND4_X1 T1918 ( .D(T9603_Y), .C(T1924_Y), .B(T1904_Y), .A(T1921_Y),     .Y(T1918_Y));
KC_NAND4_X1 T1931 ( .D(T10494_Y), .C(T6679_Y), .B(T1945_Y),     .A(T1946_Y), .Y(T1931_Y));
KC_NAND4_X1 T1937 ( .D(T10498_Y), .C(T1934_Y), .B(T1944_Y),     .A(T1956_Y), .Y(T1937_Y));
KC_NAND4_X1 T1938 ( .D(T9850_Y), .C(T1936_Y), .B(T1943_Y), .A(T1951_Y),     .Y(T1938_Y));
KC_NAND4_X1 T1939 ( .D(T10495_Y), .C(T6678_Y), .B(T1953_Y),     .A(T1948_Y), .Y(T1939_Y));
KC_NAND4_X1 T1940 ( .D(T9751_Y), .C(T1932_Y), .B(T1942_Y), .A(T1957_Y),     .Y(T1940_Y));
KC_NAND4_X1 T1941 ( .D(T10497_Y), .C(T1935_Y), .B(T1952_Y),     .A(T1947_Y), .Y(T1941_Y));
KC_NAND4_X1 T1949 ( .D(T9851_Y), .C(T1969_Y), .B(T5797_Y), .A(T1955_Y),     .Y(T1949_Y));
KC_NAND4_X1 T1950 ( .D(T10496_Y), .C(T1933_Y), .B(T1954_Y),     .A(T1958_Y), .Y(T1950_Y));
KC_NAND4_X1 T1986 ( .D(T9950_Y), .C(T5367_Y), .B(T2015_Q), .A(T2028_Q),     .Y(T1986_Y));
KC_NAND4_X1 T1987 ( .D(T1116_Y), .C(T15478_Y), .B(T2008_Q),     .A(T1997_Y), .Y(T1987_Y));
KC_NAND4_X1 T1988 ( .D(T16364_Y), .C(T2008_Q), .B(T2016_Q),     .A(T1997_Y), .Y(T1988_Y));
KC_NAND4_X1 T1995 ( .D(T16370_Y), .C(T11915_Y), .B(T10527_Y),     .A(T9972_Y), .Y(T1995_Y));
KC_NAND4_X1 T1996 ( .D(T1990_Y), .C(T15478_Y), .B(T1116_Y), .A(T868_Y),     .Y(T1996_Y));
KC_NAND4_X1 T2029 ( .D(T10111_Y), .C(T10110_Y), .B(T16291_Y),     .A(T10120_Y), .Y(T2029_Y));
KC_NAND4_X1 T2032 ( .D(T10109_Y), .C(T10108_Y), .B(T10113_Y),     .A(T10112_Y), .Y(T2032_Y));
KC_NAND4_X1 T2036 ( .D(T1506_Y), .C(T1485_Y), .B(T15503_Y),     .A(T13048_Q), .Y(T2036_Y));
KC_NAND4_X1 T2064 ( .D(T12982_Y), .C(T10934_Y), .B(T10205_Y),     .A(T1365_Y), .Y(T2064_Y));
KC_NAND4_X1 T2065 ( .D(T12750_Y), .C(T12982_Y), .B(T15535_Y),     .A(T10205_Y), .Y(T2065_Y));
KC_NAND4_X1 T2066 ( .D(T10936_Y), .C(T10942_Y), .B(T13131_Y),     .A(T15529_Y), .Y(T2066_Y));
KC_NAND4_X1 T2067 ( .D(T13125_Y), .C(T5508_Y), .B(T10184_Y),     .A(T15529_Y), .Y(T2067_Y));
KC_NAND4_X1 T2069 ( .D(T16237_Y), .C(T6593_Y), .B(T6593_Y),     .A(T16234_Y), .Y(T2069_Y));
KC_NAND4_X1 T2074 ( .D(T8313_Y), .C(T13028_Q), .B(T13292_Q),     .A(T13070_Q), .Y(T2074_Y));
KC_NAND4_X1 T2106 ( .D(T5070_Y), .C(T11489_Y), .B(T2105_Y),     .A(T12794_Y), .Y(T2106_Y));
KC_NAND4_X1 T2134 ( .D(T2137_Y), .C(T2135_Y), .B(T2136_Y), .A(T4941_Y),     .Y(T2134_Y));
KC_NAND4_X1 T2141 ( .D(T2144_Y), .C(T2143_Y), .B(T2102_Y), .A(T4945_Y),     .Y(T2141_Y));
KC_NAND4_X1 T2146 ( .D(T2142_Y), .C(T2139_Y), .B(T2147_Y), .A(T2101_Y),     .Y(T2146_Y));
KC_NAND4_X1 T2167 ( .D(T5926_Y), .C(T5924_Y), .B(T2172_Y), .A(T2172_Y),     .Y(T2167_Y));
KC_NAND4_X1 T2191 ( .D(T11026_Y), .C(T2776_Y), .B(T8297_Y),     .A(T2193_Y), .Y(T2191_Y));
KC_NAND4_X1 T2199 ( .D(T11568_Y), .C(T2775_Y), .B(T2204_Y),     .A(T2224_Y), .Y(T2199_Y));
KC_NAND4_X1 T2205 ( .D(T2780_Y), .C(T2209_Y), .B(T2196_Y), .A(T2234_Y),     .Y(T2205_Y));
KC_NAND4_X1 T2206 ( .D(T2771_Y), .C(T12217_Y), .B(T8307_Y),     .A(T4938_Y), .Y(T2206_Y));
KC_NAND4_X1 T2218 ( .D(T2797_Y), .C(T2215_Y), .B(T4959_Y), .A(T2226_Y),     .Y(T2218_Y));
KC_NAND4_X1 T2227 ( .D(T8341_Y), .C(T8315_Y), .B(T8339_Y), .A(T8327_Y),     .Y(T2227_Y));
KC_NAND4_X1 T2228 ( .D(T8309_Y), .C(T8310_Y), .B(T8282_Y), .A(T8319_Y),     .Y(T2228_Y));
KC_NAND4_X1 T2229 ( .D(T8240_Y), .C(T8473_Y), .B(T8328_Y), .A(T8343_Y),     .Y(T2229_Y));
KC_NAND4_X1 T2256 ( .D(T2283_Y), .C(T2260_Y), .B(T2253_Y), .A(T2257_Y),     .Y(T2256_Y));
KC_NAND4_X1 T2262 ( .D(T2268_Y), .C(T2267_Y), .B(T2252_Y), .A(T2258_Y),     .Y(T2262_Y));
KC_NAND4_X1 T2294 ( .D(T2274_Y), .C(T2289_Y), .B(T2288_Y), .A(T2297_Y),     .Y(T2294_Y));
KC_NAND4_X1 T2301 ( .D(T2300_Y), .C(T2303_Y), .B(T2302_Y), .A(T2265_Y),     .Y(T2301_Y));
KC_NAND4_X1 T2304 ( .D(T2299_Y), .C(T2306_Y), .B(T2305_Y), .A(T2255_Y),     .Y(T2304_Y));
KC_NAND4_X1 T2318 ( .D(T16130_Y), .C(T6225_Y), .B(T16270_Y),     .A(T10558_Y), .Y(T2318_Y));
KC_NAND4_X1 T2323 ( .D(T6243_Y), .C(T2357_Y), .B(T8410_Y), .A(T2350_Y),     .Y(T2323_Y));
KC_NAND4_X1 T2324 ( .D(T11774_Y), .C(T6232_Y), .B(T16270_Y),     .A(T12101_Y), .Y(T2324_Y));
KC_NAND4_X1 T2336 ( .D(T1832_Q), .C(T1833_Q), .B(T5527_Q), .A(T2364_Q),     .Y(T2336_Y));
KC_NAND4_X1 T2366 ( .D(T8157_Y), .C(T8436_Y), .B(T2367_Y), .A(T8436_Y),     .Y(T2366_Y));
KC_NAND4_X1 T2370 ( .D(T6505_Y), .C(T2387_Y), .B(T12319_Y),     .A(T12320_Y), .Y(T2370_Y));
KC_NAND4_X1 T2373 ( .D(T5529_Q), .C(T1857_Q), .B(T1856_Q), .A(T2388_Q),     .Y(T2373_Y));
KC_NAND4_X1 T2412 ( .D(T10465_Y), .C(T1879_Y), .B(T2402_Y),     .A(T2422_Y), .Y(T2412_Y));
KC_NAND4_X1 T2425 ( .D(T10460_Y), .C(T2419_Y), .B(T2405_Y),     .A(T2964_Y), .Y(T2425_Y));
KC_NAND4_X1 T2426 ( .D(T9527_Y), .C(T2415_Y), .B(T2404_Y), .A(T2992_Y),     .Y(T2426_Y));
KC_NAND4_X1 T2455 ( .D(T2546_Y), .C(T10812_Y), .B(T2456_Y),     .A(T2431_Y), .Y(T2455_Y));
KC_NAND4_X1 T2461 ( .D(T2617_Y), .C(T6793_Y), .B(T2463_Y), .A(T2411_Y),     .Y(T2461_Y));
KC_NAND4_X1 T2468 ( .D(T2616_Y), .C(T10828_Y), .B(T2473_Y),     .A(T2418_Y), .Y(T2468_Y));
KC_NAND4_X1 T2469 ( .D(T2603_Y), .C(T10829_Y), .B(T2471_Y),     .A(T2423_Y), .Y(T2469_Y));
KC_NAND4_X1 T2470 ( .D(T2605_Y), .C(T10833_Y), .B(T2472_Y),     .A(T2430_Y), .Y(T2470_Y));
KC_NAND4_X1 T2483 ( .D(T2600_Y), .C(T7516_Y), .B(T2487_Y), .A(T2432_Y),     .Y(T2483_Y));
KC_NAND4_X1 T2484 ( .D(T2602_Y), .C(T10813_Y), .B(T2462_Y),     .A(T2410_Y), .Y(T2484_Y));
KC_NAND4_X1 T2485 ( .D(T2606_Y), .C(T10817_Y), .B(T2486_Y),     .A(T2433_Y), .Y(T2485_Y));
KC_NAND4_X1 T2509 ( .D(T9845_Y), .C(T7725_Y), .B(T7751_Y), .A(T3664_Y),     .Y(T2509_Y));
KC_NAND4_X1 T2511 ( .D(T2555_Y), .C(T7760_Y), .B(T2519_Y), .A(T4989_Y),     .Y(T2511_Y));
KC_NAND4_X1 T2512 ( .D(T9848_Y), .C(T7708_Y), .B(T7748_Y), .A(T5287_Y),     .Y(T2512_Y));
KC_NAND4_X1 T2513 ( .D(T9847_Y), .C(T7726_Y), .B(T10781_Y),     .A(T3663_Y), .Y(T2513_Y));
KC_NAND4_X1 T2514 ( .D(T2601_Y), .C(T7762_Y), .B(T2518_Y), .A(T2421_Y),     .Y(T2514_Y));
KC_NAND4_X1 T2515 ( .D(T2594_Y), .C(T7761_Y), .B(T2517_Y), .A(T2417_Y),     .Y(T2515_Y));
KC_NAND4_X1 T2516 ( .D(T9846_Y), .C(T7767_Y), .B(T7750_Y), .A(T3665_Y),     .Y(T2516_Y));
KC_NAND4_X1 T2561 ( .D(T2547_Y), .C(T5869_S), .B(T2547_Y), .A(T2573_Y),     .Y(T2561_Y));
KC_NAND4_X1 T2567 ( .D(T5025_Q), .C(T2572_Q), .B(T2592_Q), .A(T2591_Q),     .Y(T2567_Y));
KC_NAND4_X1 T2612 ( .D(T2598_Y), .C(T13032_Y), .B(T10526_Y),     .A(T2550_Y), .Y(T2612_Y));
KC_NAND4_X1 T2679 ( .D(T2675_Y), .C(T12141_Y), .B(T11962_Y),     .A(T5020_Y), .Y(T2679_Y));
KC_NAND4_X1 T2685 ( .D(T11339_Y), .C(T5776_Y), .B(T10272_Y),     .A(T2695_Y), .Y(T2685_Y));
KC_NAND4_X1 T2699 ( .D(T15851_Y), .C(T16088_Q), .B(T15796_Q),     .A(T15809_Q), .Y(T2699_Y));
KC_NAND4_X1 T2700 ( .D(T1743_Y), .C(T15807_Q), .B(T15804_Q),     .A(T15803_Q), .Y(T2700_Y));
KC_NAND4_X1 T2701 ( .D(T15005_Y), .C(T15797_Q), .B(T964_Q),     .A(T15798_Q), .Y(T2701_Y));
KC_NAND4_X1 T2704 ( .D(T15805_Q), .C(T15808_Q), .B(T16299_Q),     .A(T15844_Q), .Y(T2704_Y));
KC_NAND4_X1 T2721 ( .D(T2748_Q), .C(T2738_Q), .B(T2749_Q), .A(T2737_Q),     .Y(T2721_Y));
KC_NAND4_X1 T2725 ( .D(T8232_Y), .C(T8233_Y), .B(T8248_Y), .A(T8227_Y),     .Y(T2725_Y));
KC_NAND4_X1 T2726 ( .D(T8495_Y), .C(T13105_Y), .B(T8225_Y),     .A(T8226_Y), .Y(T2726_Y));
KC_NAND4_X1 T2728 ( .D(T8207_Y), .C(T8216_Y), .B(T8217_Y), .A(T8218_Y),     .Y(T2728_Y));
KC_NAND4_X1 T2729 ( .D(T15895_Y), .C(T10245_Y), .B(T16299_Q),     .A(T15809_Q), .Y(T2729_Y));
KC_NAND4_X1 T2732 ( .D(T15856_Y), .C(T15805_Q), .B(T15798_Q),     .A(T15807_Q), .Y(T2732_Y));
KC_NAND4_X1 T2755 ( .D(T11464_Y), .C(T11448_Y), .B(T964_Q),     .A(T11637_Y), .Y(T2755_Y));
KC_NAND4_X1 T2770 ( .D(T5877_Y), .C(T8492_Y), .B(T11491_Y),     .A(T2791_Y), .Y(T2770_Y));
KC_NAND4_X1 T2798 ( .D(T6776_Co), .C(T12961_Y), .B(T5068_Y),     .A(T3327_Y), .Y(T2798_Y));
KC_NAND4_X1 T2818 ( .D(T5002_Y), .C(T6119_Y), .B(T15622_Y),     .A(T2841_Q), .Y(T2818_Y));
KC_NAND4_X1 T2822 ( .D(T6511_Y), .C(T6039_Y), .B(T6087_Y),     .A(T11660_Y), .Y(T2822_Y));
KC_NAND4_X1 T2825 ( .D(T16056_Y), .C(T10596_Y), .B(T2735_Q),     .A(T2830_Y), .Y(T2825_Y));
KC_NAND4_X1 T2826 ( .D(T2817_Y), .C(T11629_Y), .B(T2282_Y),     .A(T2221_Y), .Y(T2826_Y));
KC_NAND4_X1 T2827 ( .D(T11628_Y), .C(T16156_Y), .B(T11818_Y),     .A(T15802_Q), .Y(T2827_Y));
KC_NAND4_X1 T2850 ( .D(T6515_Y), .C(T11731_Y), .B(T2856_Y),     .A(T11729_Y), .Y(T2850_Y));
KC_NAND4_X1 T2868 ( .D(T5539_Y), .C(T12064_Y), .B(T3514_Y),     .A(T16135_Y), .Y(T2868_Y));
KC_NAND4_X1 T2882 ( .D(T6240_Y), .C(T12106_Y), .B(T10557_Y),     .A(T12107_Y), .Y(T2882_Y));
KC_NAND4_X1 T2883 ( .D(T12062_Y), .C(T12310_Y), .B(T5001_Y),     .A(T12364_Y), .Y(T2883_Y));
KC_NAND4_X1 T2884 ( .D(T12974_Y), .C(T12259_Y), .B(T12266_Y),     .A(T2919_Y), .Y(T2884_Y));
KC_NAND4_X1 T2885 ( .D(T2893_Y), .C(T11808_Y), .B(T12106_Y),     .A(T12306_Y), .Y(T2885_Y));
KC_NAND4_X1 T2889 ( .D(T5518_Y), .C(T2890_Y), .B(T2887_Y),     .A(T12312_Y), .Y(T2889_Y));
KC_NAND4_X1 T2890 ( .D(T4999_Y), .C(T6572_Y), .B(T16131_Y),     .A(T2354_Y), .Y(T2890_Y));
KC_NAND4_X1 T2893 ( .D(T15633_Y), .C(T16131_Y), .B(T6232_Y),     .A(T12108_Y), .Y(T2893_Y));
KC_NAND4_X1 T2894 ( .D(T6225_Y), .C(T10573_Y), .B(T12108_Y),     .A(T12101_Y), .Y(T2894_Y));
KC_NAND4_X1 T2904 ( .D(T5518_Y), .C(T2893_Y), .B(T2903_Y), .A(T5520_Y),     .Y(T2904_Y));
KC_NAND4_X1 T2905 ( .D(T2901_Y), .C(T2887_Y), .B(T2907_Y), .A(T2356_Y),     .Y(T2905_Y));
KC_NAND4_X1 T2913 ( .D(T2320_Y), .C(T12106_Y), .B(T6221_Y),     .A(T6197_Y), .Y(T2913_Y));
KC_NAND4_X1 T2917 ( .D(T11822_Y), .C(T4096_Y), .B(T4055_Y),     .A(T2941_Y), .Y(T2917_Y));
KC_NAND4_X1 T2918 ( .D(T290_Y), .C(T6531_Y), .B(T2948_Y), .A(T4055_Y),     .Y(T2918_Y));
KC_NAND4_X1 T2940 ( .D(T2935_Y), .C(T12861_Y), .B(T2916_Y),     .A(T2939_Y), .Y(T2940_Y));
KC_NAND4_X1 T2962 ( .D(T10461_Y), .C(T2427_Y), .B(T2407_Y),     .A(T2972_Y), .Y(T2962_Y));
KC_NAND4_X1 T2966 ( .D(T9528_Y), .C(T2416_Y), .B(T2406_Y), .A(T2971_Y),     .Y(T2966_Y));
KC_NAND4_X1 T2973 ( .D(T9572_Y), .C(T2977_Y), .B(T2976_Y), .A(T2986_Y),     .Y(T2973_Y));
KC_NAND4_X1 T2980 ( .D(T9571_Y), .C(T2984_Y), .B(T2979_Y), .A(T2970_Y),     .Y(T2980_Y));
KC_NAND4_X1 T2981 ( .D(T9570_Y), .C(T2983_Y), .B(T2994_Y), .A(T2967_Y),     .Y(T2981_Y));
KC_NAND4_X1 T2985 ( .D(T9569_Y), .C(T2978_Y), .B(T2987_Y), .A(T2989_Y),     .Y(T2985_Y));
KC_NAND4_X1 T2990 ( .D(T9526_Y), .C(T2420_Y), .B(T2403_Y), .A(T2995_Y),     .Y(T2990_Y));
KC_NAND4_X1 T2991 ( .D(T9529_Y), .C(T5209_Y), .B(T2965_Y), .A(T2963_Y),     .Y(T2991_Y));
KC_NAND4_X1 T3000 ( .D(T10452_Y), .C(T3007_Y), .B(T3006_Y),     .A(T3002_Y), .Y(T3000_Y));
KC_NAND4_X1 T3001 ( .D(T10451_Y), .C(T3003_Y), .B(T5552_Y),     .A(T5234_Y), .Y(T3001_Y));
KC_NAND4_X1 T3011 ( .D(T473_Y), .C(T2998_Y), .B(T5249_Y), .A(T3596_Y),     .Y(T3011_Y));
KC_NAND4_X1 T3035 ( .D(T10489_Y), .C(T3055_Y), .B(T3033_Y),     .A(T3630_Y), .Y(T3035_Y));
KC_NAND4_X1 T3036 ( .D(T10487_Y), .C(T3058_Y), .B(T3044_Y),     .A(T3042_Y), .Y(T3036_Y));
KC_NAND4_X1 T3037 ( .D(T10486_Y), .C(T3040_Y), .B(T3049_Y),     .A(T3629_Y), .Y(T3037_Y));
KC_NAND4_X1 T3038 ( .D(T9776_Y), .C(T3041_Y), .B(T3048_Y), .A(T5271_Y),     .Y(T3038_Y));
KC_NAND4_X1 T3039 ( .D(T10488_Y), .C(T3059_Y), .B(T3043_Y),     .A(T5269_Y), .Y(T3039_Y));
KC_NAND4_X1 T3052 ( .D(T10490_Y), .C(T3057_Y), .B(T3050_Y),     .A(T3046_Y), .Y(T3052_Y));
KC_NAND4_X1 T3053 ( .D(T9777_Y), .C(T3060_Y), .B(T3034_Y), .A(T3047_Y),     .Y(T3053_Y));
KC_NAND4_X1 T3082 ( .D(T10513_Y), .C(T3085_Y), .B(T3086_Y),     .A(T3084_Y), .Y(T3082_Y));
KC_NAND4_X1 T3087 ( .D(T9934_Y), .C(T3114_Y), .B(T3091_Y), .A(T3090_Y),     .Y(T3087_Y));
KC_NAND4_X1 T3094 ( .D(T9963_Y), .C(T3083_Y), .B(T3096_Y), .A(T3097_Y),     .Y(T3094_Y));
KC_NAND4_X1 T3102 ( .D(T9945_Y), .C(T3107_Y), .B(T3095_Y), .A(T3105_Y),     .Y(T3102_Y));
KC_NAND4_X1 T3103 ( .D(T9944_Y), .C(T3106_Y), .B(T3098_Y), .A(T3104_Y),     .Y(T3103_Y));
KC_NAND4_X1 T3108 ( .D(T9935_Y), .C(T3111_Y), .B(T3092_Y), .A(T3113_Y),     .Y(T3108_Y));
KC_NAND4_X1 T3109 ( .D(T9956_Y), .C(T3100_Y), .B(T3088_Y), .A(T3089_Y),     .Y(T3109_Y));
KC_NAND4_X1 T3110 ( .D(T9955_Y), .C(T3101_Y), .B(T3115_Y), .A(T3112_Y),     .Y(T3110_Y));
KC_NAND4_X1 T3129 ( .D(T10098_Y), .C(T3125_Y), .B(T3124_Y),     .A(T3135_Y), .Y(T3129_Y));
KC_NAND4_X1 T3130 ( .D(T10097_Y), .C(T3128_Y), .B(T16259_Y),     .A(T3134_Y), .Y(T3130_Y));
KC_NAND4_X1 T3137 ( .D(T10074_Y), .C(T3132_Y), .B(T3136_Y),     .A(T3139_Y), .Y(T3137_Y));
KC_NAND4_X1 T3138 ( .D(T10075_Y), .C(T3131_Y), .B(T3133_Y),     .A(T3140_Y), .Y(T3138_Y));
KC_NAND4_X1 T3145 ( .D(T10076_Y), .C(T3143_Y), .B(T3141_Y),     .A(T3731_Y), .Y(T3145_Y));
KC_NAND4_X1 T3146 ( .D(T10053_Y), .C(T3144_Y), .B(T3142_Y),     .A(T5368_Y), .Y(T3146_Y));
KC_NAND4_X1 T3161 ( .D(T10200_Y), .C(T3170_Y), .B(T3164_Y),     .A(T3165_Y), .Y(T3161_Y));
KC_NAND4_X1 T3166 ( .D(T10190_Y), .C(T3175_Y), .B(T3168_Y),     .A(T3172_Y), .Y(T3166_Y));
KC_NAND4_X1 T3167 ( .D(T10189_Y), .C(T3169_Y), .B(T3162_Y),     .A(T5401_Y), .Y(T3167_Y));
KC_NAND4_X1 T3171 ( .D(T10192_Y), .C(T3174_Y), .B(T3173_Y),     .A(T5403_Y), .Y(T3171_Y));
KC_NAND4_X1 T3176 ( .D(T16249_Y), .C(T3182_Y), .B(T3181_Y),     .A(T3179_Y), .Y(T3176_Y));
KC_NAND4_X1 T3177 ( .D(T10114_Y), .C(T3178_Y), .B(T3183_Y),     .A(T3180_Y), .Y(T3177_Y));
KC_NAND4_X1 T3248 ( .D(T15911_Y), .C(T3282_Y), .B(T8206_Y),     .A(T4384_Y), .Y(T3248_Y));
KC_NAND4_X1 T3284 ( .D(T5940_Y), .C(T15928_Y), .B(T2734_Y),     .A(T2762_Y), .Y(T3284_Y));
KC_NAND4_X1 T3319 ( .D(T15978_Y), .C(T15976_Y), .B(T2719_Y),     .A(T15977_Y), .Y(T3319_Y));
KC_NAND4_X1 T3325 ( .D(T15980_Y), .C(T3326_Y), .B(T3451_Y),     .A(T3323_Y), .Y(T3325_Y));
KC_NAND4_X1 T3348 ( .D(T6776_Co), .C(T12961_Y), .B(T5068_Y),     .A(T6776_Co), .Y(T3348_Y));
KC_NAND4_X1 T3349 ( .D(T3347_Y), .C(T3350_Y), .B(T3340_Y), .A(T5478_Y),     .Y(T3349_Y));
KC_NAND4_X1 T3371 ( .D(T10965_Y), .C(T3405_Y), .B(T3368_Y),     .A(T12247_Y), .Y(T3371_Y));
KC_NAND4_X1 T3372 ( .D(T6084_Y), .C(T6065_Y), .B(T6158_Y),     .A(T11818_Y), .Y(T3372_Y));
KC_NAND4_X1 T3373 ( .D(T12858_Y), .C(T2850_Y), .B(T11998_Y),     .A(T15622_Y), .Y(T3373_Y));
KC_NAND4_X1 T3377 ( .D(T10979_Y), .C(T16302_Y), .B(T16034_Y),     .A(T11996_Y), .Y(T3377_Y));
KC_NAND4_X1 T3378 ( .D(T6044_Y), .C(T11604_Y), .B(T12004_Y),     .A(T5525_Q), .Y(T3378_Y));
KC_NAND4_X1 T3380 ( .D(T12039_Y), .C(T12003_Y), .B(T12248_Y),     .A(T6062_Y), .Y(T3380_Y));
KC_NAND4_X1 T3381 ( .D(T6069_Y), .C(T3516_Y), .B(T6393_Y), .A(T6086_Y),     .Y(T3381_Y));
KC_NAND4_X1 T3385 ( .D(T6043_Y), .C(T6044_Y), .B(T4147_Q), .A(T6526_Q),     .Y(T3385_Y));
KC_NAND4_X1 T3386 ( .D(T11659_Y), .C(T11661_Y), .B(T11630_Y),     .A(T10590_Y), .Y(T3386_Y));
KC_NAND4_X1 T3387 ( .D(T3413_Y), .C(T10590_Y), .B(T12000_Y),     .A(T3517_Y), .Y(T3387_Y));
KC_NAND4_X1 T3388 ( .D(T8353_Y), .C(T5532_Q), .B(T3528_Q), .A(T4178_Q),     .Y(T3388_Y));
KC_NAND4_X1 T3389 ( .D(T16035_Y), .C(T6048_Y), .B(T11626_Y),     .A(T6549_Q), .Y(T3389_Y));
KC_NAND4_X1 T3390 ( .D(T6064_Y), .C(T16035_Y), .B(T12003_Y),     .A(T16148_Y), .Y(T3390_Y));
KC_NAND4_X1 T3398 ( .D(T11631_Y), .C(T16167_Y), .B(T15616_Y),     .A(T11658_Y), .Y(T3398_Y));
KC_NAND4_X1 T3402 ( .D(T6175_Y), .C(T6034_Y), .B(T11996_Y),     .A(T15760_Q), .Y(T3402_Y));
KC_NAND4_X1 T3430 ( .D(T3460_Y), .C(T12852_Y), .B(T11695_Y),     .A(T2857_Y), .Y(T3430_Y));
KC_NAND4_X1 T3431 ( .D(T3457_Y), .C(T6532_Y), .B(T3482_Y),     .A(T15622_Y), .Y(T3431_Y));
KC_NAND4_X1 T3432 ( .D(T12273_Y), .C(T2864_Y), .B(T12274_Y),     .A(T3434_Y), .Y(T3432_Y));
KC_NAND4_X1 T3433 ( .D(T2850_Y), .C(T2911_Y), .B(T16138_Y),     .A(T6087_Y), .Y(T3433_Y));
KC_NAND4_X1 T3440 ( .D(T3452_Y), .C(T3423_Y), .B(T8377_Y),     .A(T12264_Y), .Y(T3440_Y));
KC_NAND4_X1 T3441 ( .D(T2850_Y), .C(T6582_Y), .B(T16137_Y),     .A(T12264_Y), .Y(T3441_Y));
KC_NAND4_X1 T3449 ( .D(T3448_Y), .C(T16135_Y), .B(T5506_Y),     .A(T6440_Y), .Y(T3449_Y));
KC_NAND4_X1 T3462 ( .D(T2888_Y), .C(T12258_Y), .B(T3463_Y),     .A(T12364_Y), .Y(T3462_Y));
KC_NAND4_X1 T3470 ( .D(T2922_Y), .C(T3494_Y), .B(T12272_Y),     .A(T6584_Y), .Y(T3470_Y));
KC_NAND4_X1 T3482 ( .D(T6550_Y), .C(T15255_Y), .B(T6214_Y),     .A(T4164_Q), .Y(T3482_Y));
KC_NAND4_X1 T3483 ( .D(T3424_Y), .C(T6214_Y), .B(T4178_Q), .A(T3528_Q),     .Y(T3483_Y));
KC_NAND4_X1 T3484 ( .D(T6582_Y), .C(T4142_Y), .B(T12293_Y),     .A(T6564_Y), .Y(T3484_Y));
KC_NAND4_X1 T3485 ( .D(T11761_Y), .C(T3526_Y), .B(T3479_Y),     .A(T3488_Y), .Y(T3485_Y));
KC_NAND4_X1 T3486 ( .D(T6559_Y), .C(T3424_Y), .B(T15640_Y),     .A(T6550_Y), .Y(T3486_Y));
KC_NAND4_X1 T3487 ( .D(T3387_Y), .C(T6213_Y), .B(T3476_Y), .A(T3492_Y),     .Y(T3487_Y));
KC_NAND4_X1 T3513 ( .D(T6512_Y), .C(T3523_Q), .B(T3519_Q), .A(T3525_Q),     .Y(T3513_Y));
KC_NAND4_X1 T3516 ( .D(T6529_Y), .C(T11041_Y), .B(T11823_Y),     .A(T11043_Y), .Y(T3516_Y));
KC_NAND4_X1 T3536 ( .D(T9522_Y), .C(T3550_Y), .B(T3572_Y), .A(T3540_Y),     .Y(T3536_Y));
KC_NAND4_X1 T3544 ( .D(T10450_Y), .C(T3546_Y), .B(T3563_Y),     .A(T5089_Y), .Y(T3544_Y));
KC_NAND4_X1 T3545 ( .D(T9566_Y), .C(T3547_Y), .B(T3556_Y), .A(T5090_Y),     .Y(T3545_Y));
KC_NAND4_X1 T3548 ( .D(T10458_Y), .C(T3561_Y), .B(T3552_Y),     .A(T3569_Y), .Y(T3548_Y));
KC_NAND4_X1 T3549 ( .D(T10459_Y), .C(T3558_Y), .B(T3551_Y),     .A(T3568_Y), .Y(T3549_Y));
KC_NAND4_X1 T3564 ( .D(T9523_Y), .C(T3553_Y), .B(T3570_Y), .A(T3541_Y),     .Y(T3564_Y));
KC_NAND4_X1 T3565 ( .D(T9524_Y), .C(T3554_Y), .B(T3571_Y), .A(T3537_Y),     .Y(T3565_Y));
KC_NAND4_X1 T3566 ( .D(T9525_Y), .C(T3555_Y), .B(T3567_Y), .A(T3538_Y),     .Y(T3566_Y));
KC_NAND4_X1 T3578 ( .D(T9565_Y), .C(T3583_Y), .B(T5091_Y), .A(T3581_Y),     .Y(T3578_Y));
KC_NAND4_X1 T3579 ( .D(T10449_Y), .C(T3580_Y), .B(T5092_Y),     .A(T3582_Y), .Y(T3579_Y));
KC_NAND4_X1 T3586 ( .D(T9662_Y), .C(T5733_Y), .B(T5098_Y), .A(T3597_Y),     .Y(T3586_Y));
KC_NAND4_X1 T3587 ( .D(T474_Y), .C(T3577_Y), .B(T5096_Y), .A(T3601_Y),     .Y(T3587_Y));
KC_NAND4_X1 T3588 ( .D(T9660_Y), .C(T3576_Y), .B(T5095_Y), .A(T3602_Y),     .Y(T3588_Y));
KC_NAND4_X1 T3589 ( .D(T9661_Y), .C(T5231_Y), .B(T3606_Y), .A(T3598_Y),     .Y(T3589_Y));
KC_NAND4_X1 T3603 ( .D(T9634_Y), .C(T3573_Y), .B(T5094_Y), .A(T3600_Y),     .Y(T3603_Y));
KC_NAND4_X1 T3604 ( .D(T10435_Y), .C(T3574_Y), .B(T5093_Y),     .A(T3590_Y), .Y(T3604_Y));
KC_NAND4_X1 T3605 ( .D(T10434_Y), .C(T3575_Y), .B(T5097_Y),     .A(T3595_Y), .Y(T3605_Y));
KC_NAND4_X1 T3614 ( .D(T10466_Y), .C(T6847_Y), .B(T4230_Y),     .A(T3616_Y), .Y(T3614_Y));
KC_NAND4_X1 T3617 ( .D(T9724_Y), .C(T3618_Y), .B(T4239_Y), .A(T3620_Y),     .Y(T3617_Y));
KC_NAND4_X1 T3622 ( .D(T8518_Y), .C(T3624_Y), .B(T3632_Y), .A(T3615_Y),     .Y(T3622_Y));
KC_NAND4_X1 T3627 ( .D(T10469_Y), .C(T3625_Y), .B(T4249_Y),     .A(T3633_Y), .Y(T3627_Y));
KC_NAND4_X1 T3628 ( .D(T8519_Y), .C(T3637_Y), .B(T5551_Y), .A(T5085_Y),     .Y(T3628_Y));
KC_NAND4_X1 T3655 ( .D(T9856_Y), .C(T3660_Y), .B(T3661_Y), .A(T3658_Y),     .Y(T3655_Y));
KC_NAND4_X1 T3656 ( .D(T9857_Y), .C(T3659_Y), .B(T4273_Y), .A(T3662_Y),     .Y(T3656_Y));
KC_NAND4_X1 T3669 ( .D(T9820_Y), .C(T3652_Y), .B(T3674_Y), .A(T3672_Y),     .Y(T3669_Y));
KC_NAND4_X1 T3670 ( .D(T9821_Y), .C(T3671_Y), .B(T3675_Y), .A(T3673_Y),     .Y(T3670_Y));
KC_NAND4_X1 T3685 ( .D(T10051_Y), .C(T6688_Y), .B(T3702_Y),     .A(T3686_Y), .Y(T3685_Y));
KC_NAND4_X1 T3688 ( .D(T10499_Y), .C(T3689_Y), .B(T3716_Y),     .A(T3691_Y), .Y(T3688_Y));
KC_NAND4_X1 T3692 ( .D(T10073_Y), .C(T3697_Y), .B(T3706_Y),     .A(T3693_Y), .Y(T3692_Y));
KC_NAND4_X1 T3708 ( .D(T10072_Y), .C(T3710_Y), .B(T3705_Y),     .A(T6689_Y), .Y(T3708_Y));
KC_NAND4_X1 T3709 ( .D(T10512_Y), .C(T3696_Y), .B(T3711_Y),     .A(T3700_Y), .Y(T3709_Y));
KC_NAND4_X1 T3713 ( .D(T9929_Y), .C(T3690_Y), .B(T3714_Y), .A(T3717_Y),     .Y(T3713_Y));
KC_NAND4_X1 T3720 ( .D(T10117_Y), .C(T3126_Y), .B(T3721_Y),     .A(T3725_Y), .Y(T3720_Y));
KC_NAND4_X1 T3738 ( .D(T10191_Y), .C(T3753_Y), .B(T3747_Y),     .A(T5402_Y), .Y(T3738_Y));
KC_NAND4_X1 T3739 ( .D(T10198_Y), .C(T3751_Y), .B(T3744_Y),     .A(T3163_Y), .Y(T3739_Y));
KC_NAND4_X1 T3740 ( .D(T10197_Y), .C(T5976_Y), .B(T3737_Y),     .A(T3755_Y), .Y(T3740_Y));
KC_NAND4_X1 T3741 ( .D(T10196_Y), .C(T3748_Y), .B(T3745_Y),     .A(T3752_Y), .Y(T3741_Y));
KC_NAND4_X1 T3742 ( .D(T10199_Y), .C(T3743_Y), .B(T3746_Y),     .A(T3749_Y), .Y(T3742_Y));
KC_NAND4_X1 T3750 ( .D(T10533_Y), .C(T5977_Y), .B(T3736_Y),     .A(T3754_Y), .Y(T3750_Y));
KC_NAND4_X1 T3760 ( .D(T10177_Y), .C(T3770_Y), .B(T3767_Y),     .A(T3758_Y), .Y(T3760_Y));
KC_NAND4_X1 T3761 ( .D(T10176_Y), .C(T3765_Y), .B(T3764_Y),     .A(T3757_Y), .Y(T3761_Y));
KC_NAND4_X1 T3762 ( .D(T10179_Y), .C(T3772_Y), .B(T3768_Y),     .A(T3756_Y), .Y(T3762_Y));
KC_NAND4_X1 T3763 ( .D(T10178_Y), .C(T3766_Y), .B(T3771_Y),     .A(T3759_Y), .Y(T3763_Y));
KC_NAND4_X1 T3798 ( .D(T10893_Y), .C(T3796_Y), .B(T5840_Y),     .A(T8186_Y), .Y(T3798_Y));
KC_NAND4_X1 T3799 ( .D(T15847_Y), .C(T15846_Y), .B(T12130_Y),     .A(T8186_Y), .Y(T3799_Y));
KC_NAND4_X1 T3807 ( .D(T3805_Y), .C(T3818_Y), .B(T5769_Y),     .A(T12139_Y), .Y(T3807_Y));
KC_NAND4_X1 T3808 ( .D(T3801_Y), .C(T5755_Y), .B(T3811_Y), .A(T3820_Y),     .Y(T3808_Y));
KC_NAND4_X1 T3809 ( .D(T11329_Y), .C(T10892_Y), .B(T4400_Y),     .A(T5104_Y), .Y(T3809_Y));
KC_NAND4_X1 T3810 ( .D(T3804_Y), .C(T15835_Y), .B(T12145_Y),     .A(T3823_Y), .Y(T3810_Y));
KC_NAND4_X1 T3812 ( .D(T3818_Y), .C(T15825_Y), .B(T15833_Y),     .A(T15836_Y), .Y(T3812_Y));
KC_NAND4_X1 T3837 ( .D(T10911_Y), .C(T3832_Y), .B(T3841_Y),     .A(T3836_Y), .Y(T3837_Y));
KC_NAND4_X1 T3844 ( .D(T11374_Y), .C(T10903_Y), .B(T12158_Y),     .A(T4390_Y), .Y(T3844_Y));
KC_NAND4_X1 T3845 ( .D(T4461_Y), .C(T3846_Y), .B(T6740_Y),     .A(T11427_Y), .Y(T3845_Y));
KC_NAND4_X1 T3861 ( .D(T3872_Y), .C(T3889_Q), .B(T3890_Q), .A(T3873_Q),     .Y(T3861_Y));
KC_NAND4_X1 T3870 ( .D(T3884_Q), .C(T3889_Q), .B(T3890_Q), .A(T3873_Q),     .Y(T3870_Y));
KC_NAND4_X1 T3903 ( .D(T11021_Y), .C(T5889_Y), .B(T3901_Y),     .A(T11524_Y), .Y(T3903_Y));
KC_NAND4_X1 T3907 ( .D(T5986_Y), .C(T12205_Y), .B(T11556_Y),     .A(T3965_Q), .Y(T3907_Y));
KC_NAND4_X1 T3908 ( .D(T12025_Y), .C(T15580_Y), .B(T12200_Y),     .A(T8254_Y), .Y(T3908_Y));
KC_NAND4_X1 T3909 ( .D(T11510_Y), .C(T15956_Y), .B(T11495_Y),     .A(T5905_Y), .Y(T3909_Y));
KC_NAND4_X1 T3910 ( .D(T3930_Y), .C(T11496_Y), .B(T11513_Y),     .A(T11523_Y), .Y(T3910_Y));
KC_NAND4_X1 T3979 ( .D(T6025_Y), .C(T15996_Y), .B(T5122_Y),     .A(T5022_Y), .Y(T3979_Y));
KC_NAND4_X1 T4018 ( .D(T11671_Y), .C(T12045_Y), .B(T5525_Q),     .A(T6555_Q), .Y(T4018_Y));
KC_NAND4_X1 T4019 ( .D(T8509_Y), .C(T8359_Y), .B(T6045_Y),     .A(T12043_Y), .Y(T4019_Y));
KC_NAND4_X1 T4020 ( .D(T8391_Y), .C(T8506_Y), .B(T8274_Y), .A(T8372_Y),     .Y(T4020_Y));
KC_NAND4_X1 T4021 ( .D(T6079_Y), .C(T6034_Y), .B(T6062_Y), .A(T5525_Q),     .Y(T4021_Y));
KC_NAND4_X1 T4026 ( .D(T8360_Y), .C(T8357_Y), .B(T8371_Y), .A(T8356_Y),     .Y(T4026_Y));
KC_NAND4_X1 T4027 ( .D(T6045_Y), .C(T6047_Y), .B(T4147_Q), .A(T5530_Q),     .Y(T4027_Y));
KC_NAND4_X1 T4063 ( .D(T4069_Y), .C(T6181_Y), .B(T6176_Y), .A(T6155_Y),     .Y(T4063_Y));
KC_NAND4_X1 T4064 ( .D(T4105_Y), .C(T15613_Y), .B(T3382_Y),     .A(T4112_Y), .Y(T4064_Y));
KC_NAND4_X1 T4070 ( .D(T6175_Y), .C(T6043_Y), .B(T15760_Q),     .A(T6526_Q), .Y(T4070_Y));
KC_NAND4_X1 T4072 ( .D(T6148_Y), .C(T4103_Y), .B(T4698_Y), .A(T4716_Y),     .Y(T4072_Y));
KC_NAND4_X1 T4080 ( .D(T6111_Y), .C(T6134_Y), .B(T6107_Y),     .A(T11710_Y), .Y(T4080_Y));
KC_NAND4_X1 T4086 ( .D(T4099_Y), .C(T10580_Y), .B(T10582_Y),     .A(T12262_Y), .Y(T4086_Y));
KC_NAND4_X1 T4094 ( .D(T4092_Y), .C(T16141_Y), .B(T12262_Y),     .A(T10579_Y), .Y(T4094_Y));
KC_NAND4_X1 T4107 ( .D(T4136_Y), .C(T10565_Y), .B(T16128_Y),     .A(T4090_Y), .Y(T4107_Y));
KC_NAND4_X1 T4108 ( .D(T4082_Y), .C(T12857_Y), .B(T12865_Y),     .A(T4118_Y), .Y(T4108_Y));
KC_NAND4_X1 T4109 ( .D(T8512_Y), .C(T8514_Y), .B(T6560_Y),     .A(T11814_Y), .Y(T4109_Y));
KC_NAND4_X1 T4145 ( .D(T4141_Y), .C(T3464_Y), .B(T4115_Y), .A(T6536_Y),     .Y(T4145_Y));
KC_NAND4_X1 T4161 ( .D(T4166_Y), .C(T4173_Y), .B(T4165_Y), .A(T4150_Y),     .Y(T4161_Y));
KC_NAND4_X1 T4231 ( .D(T9726_Y), .C(T4238_Y), .B(T4236_Y), .A(T4237_Y),     .Y(T4231_Y));
KC_NAND4_X1 T4232 ( .D(T9775_Y), .C(T4253_Y), .B(T4235_Y), .A(T5136_Y),     .Y(T4232_Y));
KC_NAND4_X1 T4240 ( .D(T9762_Y), .C(T4241_Y), .B(T4245_Y), .A(T4247_Y),     .Y(T4240_Y));
KC_NAND4_X1 T4250 ( .D(T9761_Y), .C(T4242_Y), .B(T4243_Y), .A(T4246_Y),     .Y(T4250_Y));
KC_NAND4_X1 T4251 ( .D(T10468_Y), .C(T4254_Y), .B(T4258_Y),     .A(T4259_Y), .Y(T4251_Y));
KC_NAND4_X1 T4252 ( .D(T10467_Y), .C(T4261_Y), .B(T4262_Y),     .A(T4255_Y), .Y(T4252_Y));
KC_NAND4_X1 T5882 ( .D(T9959_Y), .C(T4297_Y), .B(T4303_Y), .A(T4313_Y),     .Y(T5882_Y));
KC_NAND4_X1 T4290 ( .D(T9952_Y), .C(T4298_Y), .B(T4302_Y), .A(T4292_Y),     .Y(T4290_Y));
KC_NAND4_X1 T4291 ( .D(T9960_Y), .C(T4296_Y), .B(T4305_Y), .A(T4312_Y),     .Y(T4291_Y));
KC_NAND4_X1 T4306 ( .D(T9930_Y), .C(T5323_Y), .B(T5855_Y), .A(T4314_Y),     .Y(T4306_Y));
KC_NAND4_X1 T4307 ( .D(T9931_Y), .C(T5332_Y), .B(T4308_Y), .A(T4309_Y),     .Y(T4307_Y));
KC_NAND4_X1 T4395 ( .D(T420_Y), .C(T420_Y), .B(T420_Y), .A(T4397_Y),     .Y(T4395_Y));
KC_NAND4_X1 T4396 ( .D(T4387_Y), .C(T4393_Y), .B(T5781_Y), .A(T4398_Y),     .Y(T4396_Y));
KC_NAND4_X1 T4433 ( .D(T3831_Y), .C(T5840_Y), .B(T12172_Y),     .A(T8194_Y), .Y(T4433_Y));
KC_NAND4_X1 T4442 ( .D(T4458_Y), .C(T12156_Y), .B(T4443_Y),     .A(T6117_Y), .Y(T4442_Y));
KC_NAND4_X1 T4453 ( .D(T5821_Y), .C(T11428_Y), .B(T14550_Q),     .A(T4463_Y), .Y(T4453_Y));
KC_NAND4_X1 T4472 ( .D(T15570_Y), .C(T4483_Y), .B(T5932_Y),     .A(T4497_Y), .Y(T4472_Y));
KC_NAND4_X1 T4473 ( .D(T15570_Y), .C(T10629_Y), .B(T4497_Y),     .A(T4484_Q), .Y(T4473_Y));
KC_NAND4_X1 T4509 ( .D(T11021_Y), .C(T12816_Y), .B(T15968_Y),     .A(T4508_Y), .Y(T4509_Y));
KC_NAND4_X1 T4511 ( .D(T11504_Y), .C(T12355_Y), .B(T5946_Y),     .A(T4475_Y), .Y(T4511_Y));
KC_NAND4_X1 T4546 ( .D(T15703_Y), .C(T15584_Y), .B(T4573_Q),     .A(T4572_Q), .Y(T4546_Y));
KC_NAND4_X1 T4548 ( .D(T4549_Y), .C(T4551_Y), .B(T11570_Y),     .A(T11534_Y), .Y(T4548_Y));
KC_NAND4_X1 T4551 ( .D(T12016_Y), .C(T4575_Q), .B(T4572_Q),     .A(T11538_Y), .Y(T4551_Y));
KC_NAND4_X1 T4554 ( .D(T3860_Y), .C(T4559_Y), .B(T12212_Y),     .A(T12222_Y), .Y(T4554_Y));
KC_NAND4_X1 T4555 ( .D(T5149_Y), .C(T3960_Y), .B(T159_Y), .A(T11534_Y),     .Y(T4555_Y));
KC_NAND4_X1 T4559 ( .D(T5954_Y), .C(T11540_Y), .B(T12016_Y),     .A(T4578_Q), .Y(T4559_Y));
KC_NAND4_X1 T4560 ( .D(T11541_Y), .C(T4579_Q), .B(T4573_Q),     .A(T4578_Q), .Y(T4560_Y));
KC_NAND4_X1 T4583 ( .D(T4587_Y), .C(T4607_Q), .B(T5158_Q), .A(T4606_Q),     .Y(T4583_Y));
KC_NAND4_X1 T4584 ( .D(T6021_Y), .C(T4586_Y), .B(T4602_Q), .A(T4607_Q),     .Y(T4584_Y));
KC_NAND4_X1 T4593 ( .D(T4594_Y), .C(T8331_Y), .B(T6012_Y), .A(T3308_Y),     .Y(T4593_Y));
KC_NAND4_X1 T4641 ( .D(T4661_Y), .C(T8366_Y), .B(T4665_Y), .A(T4668_Y),     .Y(T4641_Y));
KC_NAND4_X1 T4649 ( .D(T4631_Y), .C(T6166_Y), .B(T8458_Y),     .A(T12031_Y), .Y(T4649_Y));
KC_NAND4_X1 T4650 ( .D(T4636_Y), .C(T6166_Y), .B(T8462_Y),     .A(T12031_Y), .Y(T4650_Y));
KC_NAND4_X1 T4651 ( .D(T4635_Y), .C(T6166_Y), .B(T8461_Y),     .A(T12031_Y), .Y(T4651_Y));
KC_NAND4_X1 T4695 ( .D(T8499_Y), .C(T392_Y), .B(T8501_Y), .A(T2642_Y),     .Y(T4695_Y));
KC_NAND4_X1 T4696 ( .D(T262_Y), .C(T394_Y), .B(T258_Y), .A(T408_Y),     .Y(T4696_Y));
KC_NAND4_X1 T4699 ( .D(T4648_Y), .C(T4710_Y), .B(T4724_Y),     .A(T16122_Y), .Y(T4699_Y));
KC_NAND4_X1 T4701 ( .D(T8500_Y), .C(T412_Y), .B(T263_Y), .A(T267_Y),     .Y(T4701_Y));
KC_NAND4_X1 T4704 ( .D(T11706_Y), .C(T4719_Q), .B(T4722_Q),     .A(T4720_Q), .Y(T4704_Y));
KC_NAND4_X1 T4707 ( .D(T15141_Y), .C(T6103_Y), .B(T12033_Y),     .A(T16145_Y), .Y(T4707_Y));
KC_NAND4_X1 T4730 ( .D(T15634_Y), .C(T6103_Y), .B(T10599_Y),     .A(T6244_Y), .Y(T4730_Y));
KC_NAND4_X1 T4734 ( .D(T15630_Y), .C(T15625_Y), .B(T4757_Q),     .A(T4758_Q), .Y(T4734_Y));
KC_NAND4_X1 T4735 ( .D(T6202_Y), .C(T4756_Q), .B(T4743_Y), .A(T4755_Q),     .Y(T4735_Y));
KC_NAND4_X1 T4736 ( .D(T15630_Y), .C(T4757_Q), .B(T4756_Q),     .A(T4743_Y), .Y(T4736_Y));
KC_NAND4_X1 T4739 ( .D(T15625_Y), .C(T4740_Y), .B(T4759_Q),     .A(T4758_Q), .Y(T4739_Y));
KC_NAND4_X1 T4742 ( .D(T286_Y), .C(T4740_Y), .B(T4759_Q), .A(T4760_Q),     .Y(T4742_Y));
KC_NAND4_X1 T9396 ( .D(T9399_Y), .C(T15656_Y), .B(T9392_Y),     .A(T9390_Y), .Y(T9396_Y));
KC_NAND4_X1 T9336 ( .D(T7360_Y), .C(T7368_Y), .B(T6658_Y), .A(T7595_Y),     .Y(T9336_Y));
KC_NAND4_X1 T9335 ( .D(T6654_Y), .C(T7362_Y), .B(T6656_Y), .A(T7594_Y),     .Y(T9335_Y));
KC_NAND4_X1 T9315 ( .D(T6702_Y), .C(T6622_Y), .B(T6698_Y), .A(T6695_Y),     .Y(T9315_Y));
KC_NAND4_X1 T9443 ( .D(T1416_Y), .C(T16279_Y), .B(T15799_Y),     .A(T1554_Y), .Y(T9443_Y));
KC_NAND4_X1 T9327 ( .D(T11873_Y), .C(T11874_Y), .B(T15742_Y),     .A(T7442_Y), .Y(T9327_Y));
KC_NAND4_X1 T9314 ( .D(T6638_Y), .C(T6629_Y), .B(T6625_Y),     .A(T15659_Y), .Y(T9314_Y));
KC_NAND4_X1 T10301 ( .D(T10880_Y), .C(T10942_Y), .B(T4872_Y),     .A(T10161_Y), .Y(T10301_Y));
KC_NAND4_X1 T10374 ( .D(T10430_Y), .C(T10834_Y), .B(T5682_Y),     .A(T10826_Y), .Y(T10374_Y));
KC_NAND4_X1 T10302 ( .D(T10934_Y), .C(T10163_Y), .B(T10155_Y),     .A(T1362_Y), .Y(T10302_Y));
KC_NAND4_X1 T10373 ( .D(T9623_Y), .C(T10815_Y), .B(T5675_Y),     .A(T10818_Y), .Y(T10373_Y));
KC_NAND4_X1 T10371 ( .D(T9624_Y), .C(T10819_Y), .B(T10816_Y),     .A(T7514_Y), .Y(T10371_Y));
KC_NAND4_X1 T10338 ( .D(T10337_Y), .C(T7464_Y), .B(T7492_Y),     .A(T7545_Y), .Y(T10338_Y));
KC_NAND4_X1 T10365 ( .D(T9709_Y), .C(T10801_Y), .B(T5657_Y),     .A(T10802_Y), .Y(T10365_Y));
KC_NAND4_X1 T10333 ( .D(T9795_Y), .C(T10777_Y), .B(T10779_Y),     .A(T10765_Y), .Y(T10333_Y));
KC_NAND4_X1 T10399 ( .D(T10395_Y), .C(T7173_Y), .B(T10874_Y),     .A(T10872_Y), .Y(T10399_Y));
KC_NAND4_X1 T10398 ( .D(T10396_Y), .C(T7172_Y), .B(T10875_Y),     .A(T10873_Y), .Y(T10398_Y));
KC_NAND4_X1 T4911 ( .D(T2279_Y), .C(T2250_Y), .B(T2246_Y), .A(T4968_Y),     .Y(T4911_Y));
KC_NAND4_X1 T4936 ( .D(T10521_Y), .C(T1142_Y), .B(T5891_Y),     .A(T16365_Y), .Y(T4936_Y));
KC_NAND4_X1 T4947 ( .D(T2816_Y), .C(T2282_Y), .B(T2254_Y), .A(T4953_Y),     .Y(T4947_Y));
KC_NAND4_X1 T4948 ( .D(T2284_Y), .C(T2292_Y), .B(T2291_Y), .A(T2270_Y),     .Y(T4948_Y));
KC_NAND4_X1 T4949 ( .D(T2266_Y), .C(T4946_Y), .B(T5489_Y), .A(T4952_Y),     .Y(T4949_Y));
KC_NAND4_X1 T4950 ( .D(T2271_Y), .C(T2290_Y), .B(T2286_Y), .A(T2269_Y),     .Y(T4950_Y));
KC_NAND4_X1 T4955 ( .D(T2769_Y), .C(T4958_Y), .B(T4940_Y), .A(T2233_Y),     .Y(T4955_Y));
KC_NAND4_X1 T4987 ( .D(T2553_Y), .C(T7466_Y), .B(T4988_Y), .A(T2414_Y),     .Y(T4987_Y));
KC_NAND4_X1 T4996 ( .D(T5019_Y), .C(T15755_Y), .B(T6017_Y),     .A(T5020_Y), .Y(T4996_Y));
KC_NAND4_X1 T5004 ( .D(T5003_Y), .C(T3415_Y), .B(T6077_Y),     .A(T12048_Y), .Y(T5004_Y));
KC_NAND4_X1 T5033 ( .D(T9567_Y), .C(T5035_Y), .B(T2975_Y), .A(T3005_Y),     .Y(T5033_Y));
KC_NAND4_X1 T5034 ( .D(T9568_Y), .C(T5036_Y), .B(T2974_Y), .A(T3004_Y),     .Y(T5034_Y));
KC_NAND4_X1 T5053 ( .D(T11703_Y), .C(T5004_Y), .B(T3376_Y),     .A(T3397_Y), .Y(T5053_Y));
KC_NAND4_X1 T5054 ( .D(T5522_Y), .C(T5523_Y), .B(T12046_Y),     .A(T11676_Y), .Y(T5054_Y));
KC_NAND4_X1 T5055 ( .D(T4104_Y), .C(T5004_Y), .B(T10610_Y),     .A(T16107_Y), .Y(T5055_Y));
KC_NAND4_X1 T16258 ( .D(T10116_Y), .C(T3127_Y), .B(T3769_Y),     .A(T3724_Y), .Y(T16258_Y));
KC_NAND4_X1 T5083 ( .D(T8517_Y), .C(T3634_Y), .B(T5267_Y), .A(T3609_Y),     .Y(T5083_Y));
KC_NAND4_X1 T5084 ( .D(T8516_Y), .C(T3631_Y), .B(T5086_Y), .A(T5087_Y),     .Y(T5084_Y));
KC_NAND4_X1 T5100 ( .D(T5986_Y), .C(T15587_Y), .B(T15961_Y),     .A(T3974_Q), .Y(T5100_Y));
KC_NAND4_X1 T5113 ( .D(T16027_Y), .C(T4009_Y), .B(T4030_Y),     .A(T12235_Y), .Y(T5113_Y));
KC_NAND4_X1 T5146 ( .D(T259_Y), .C(T261_Y), .B(T4157_Y), .A(T241_Y),     .Y(T5146_Y));
KC_NAND4_X1 T5149 ( .D(T15703_Y), .C(T5952_Y), .B(T11541_Y),     .A(T4573_Q), .Y(T5149_Y));
KC_NAND4_X1 T5150 ( .D(T4688_Y), .C(T4688_Y), .B(T12345_Y),     .A(T16045_Y), .Y(T5150_Y));
KC_NAND4_X1 T5629 ( .D(T54_Q), .C(T5220_Q), .B(T5611_Y), .A(T55_Y),     .Y(T5629_Y));
KC_NAND4_X1 T9290 ( .D(T6318_Y), .C(T9271_Y), .B(T150_Q), .A(T5222_Q),     .Y(T9290_Y));
KC_NAND4_X1 T9282 ( .D(T6292_Y), .C(T6291_Y), .B(T6296_Y), .A(T6294_Y),     .Y(T9282_Y));
KC_NAND4_X1 T6944 ( .D(T236_Y), .C(T9271_Y), .B(T5225_Q), .A(T5222_Q),     .Y(T6944_Y));
KC_NAND4_X1 T6933 ( .D(T236_Y), .C(T8577_Y), .B(T8580_Y), .A(T5225_Q),     .Y(T6933_Y));
KC_NAND4_X1 T6931 ( .D(T284_Q), .C(T278_Q), .B(T294_Q), .A(T272_Q),     .Y(T6931_Y));
KC_NAND4_X1 T5208 ( .D(T10462_Y), .C(T2413_Y), .B(T1881_Y),     .A(T5212_Y), .Y(T5208_Y));
KC_NAND4_X1 T7119 ( .D(T12403_Y), .C(T8626_Y), .B(T8572_Y),     .A(T12477_Y), .Y(T7119_Y));
KC_NAND4_X1 T9510 ( .D(T668_Q), .C(T665_Q), .B(T694_Q), .A(T663_Q),     .Y(T9510_Y));
KC_NAND4_X1 T7255 ( .D(T7308_Y), .C(T6472_Y), .B(T7251_Y), .A(T7247_Y),     .Y(T7255_Y));
KC_NAND4_X1 T5679 ( .D(T9622_Y), .C(T5677_Y), .B(T5676_Y),     .A(T10822_Y), .Y(T5679_Y));
KC_NAND4_X1 T5268 ( .D(T9725_Y), .C(T3619_Y), .B(T4260_Y), .A(T3613_Y),     .Y(T5268_Y));
KC_NAND4_X1 T5270 ( .D(T16201_Y), .C(T15681_Y), .B(T15681_Y),     .A(T15681_Y), .Y(T5270_Y));
KC_NAND4_X1 T7653 ( .D(T7647_Y), .C(T518_Y), .B(T12437_Y),     .A(T12615_Y), .Y(T7653_Y));
KC_NAND4_X1 T5321 ( .D(T10516_Y), .C(T2631_Q), .B(T10523_Y),     .A(T1997_Y), .Y(T5321_Y));
KC_NAND4_X1 T5322 ( .D(T10050_Y), .C(T3687_Y), .B(T3701_Y),     .A(T4289_Y), .Y(T5322_Y));
KC_NAND4_X1 T5325 ( .D(T1508_Y), .C(T5365_Q), .B(T9969_Y),     .A(T10523_Y), .Y(T5325_Y));
KC_NAND4_X1 T5327 ( .D(T10052_Y), .C(T3695_Y), .B(T5328_Y),     .A(T4299_Y), .Y(T5327_Y));
KC_NAND4_X1 T5411 ( .D(T10217_Y), .C(T10231_Y), .B(T10233_Y),     .A(T10232_Y), .Y(T5411_Y));
KC_NAND4_X1 T5412 ( .D(T10214_Y), .C(T10286_Y), .B(T10216_Y),     .A(T10208_Y), .Y(T5412_Y));
KC_NAND4_X1 T5426 ( .D(T10242_Y), .C(T3793_Y), .B(T6031_Co),     .A(T15554_Y), .Y(T5426_Y));
KC_NAND4_X1 T5446 ( .D(T5854_Y), .C(T5838_Y), .B(T11365_Y),     .A(T14548_Q), .Y(T5446_Y));
KC_NAND4_X1 T5477 ( .D(T10956_Y), .C(T6020_Y), .B(T4584_Y),     .A(T11617_Y), .Y(T5477_Y));
KC_NAND4_X1 T5492 ( .D(T2230_Y), .C(T11650_Y), .B(T8347_Y),     .A(T8470_Y), .Y(T5492_Y));
KC_NAND4_X1 T5503 ( .D(T6159_Y), .C(T3436_Y), .B(T6120_Y), .A(T5522_Y),     .Y(T5503_Y));
KC_NAND4_X1 T5518 ( .D(T16130_Y), .C(T6225_Y), .B(T6240_Y),     .A(T11774_Y), .Y(T5518_Y));
KC_NAND4_X1 T5523 ( .D(T6530_Y), .C(T11037_Y), .B(T11041_Y),     .A(T2941_Y), .Y(T5523_Y));
KC_NAND4_X1 T5549 ( .D(T10528_Y), .C(T4905_Y), .B(T1989_Y),     .A(T15811_Y), .Y(T5549_Y));
KC_AOI22_X1 T7671 ( .Y(T7671_Y), .B1(T743_Y), .B0(T212_Q),     .A1(T7833_Y), .A0(T7677_Y));
KC_AOI22_X1 T4804 ( .Y(T4804_Y), .B1(T9135_Y), .B0(T4818_Y),     .A1(T15100_Y), .A0(T15150_Y));
KC_AOI22_X1 T6315 ( .Y(T6315_Y), .B1(T7364_Y), .B0(T284_Q),     .A1(T8384_Y), .A0(T293_Q));
KC_AOI22_X1 T6963 ( .Y(T6963_Y), .B1(T15311_Y), .B0(T289_Q),     .A1(T15737_Y), .A0(T275_Q));
KC_AOI22_X1 T6962 ( .Y(T6962_Y), .B1(T15311_Y), .B0(T278_Q),     .A1(T15737_Y), .A0(T296_Q));
KC_AOI22_X1 T6928 ( .Y(T6928_Y), .B1(T6801_Y), .B0(T277_Q),     .A1(T6821_Y), .A0(T288_Q));
KC_AOI22_X1 T6475 ( .Y(T6475_Y), .B1(T6801_Y), .B0(T151_Q),     .A1(T6821_Y), .A0(T5237_Q));
KC_AOI22_X1 T6474 ( .Y(T6474_Y), .B1(T15739_Y), .B0(T154_Q),     .A1(T8389_Y), .A0(T4823_Q));
KC_AOI22_X1 T6473 ( .Y(T6473_Y), .B1(T15739_Y), .B0(T282_Q),     .A1(T8389_Y), .A0(T306_Q));
KC_AOI22_X1 T7100 ( .Y(T7100_Y), .B1(T12409_Y), .B0(T4822_Q),     .A1(T12408_Y), .A0(T158_Q));
KC_AOI22_X1 T7099 ( .Y(T7099_Y), .B1(T15739_Y), .B0(T294_Q),     .A1(T8389_Y), .A0(T5241_Q));
KC_AOI22_X1 T7098 ( .Y(T7098_Y), .B1(T7364_Y), .B0(T157_Q),     .A1(T8384_Y), .A0(T5239_Q));
KC_AOI22_X1 T7086 ( .Y(T7086_Y), .B1(T6818_Y), .B0(T5562_Q),     .A1(T6828_Y), .A0(T158_Q));
KC_AOI22_X1 T7070 ( .Y(T7070_Y), .B1(T7364_Y), .B0(T5242_Q),     .A1(T8384_Y), .A0(T313_Q));
KC_AOI22_X1 T7066 ( .Y(T7066_Y), .B1(T12426_Y), .B0(T313_Q),     .A1(T12424_Y), .A0(T275_Q));
KC_AOI22_X1 T7065 ( .Y(T7065_Y), .B1(T12426_Y), .B0(T293_Q),     .A1(T12424_Y), .A0(T296_Q));
KC_AOI22_X1 T7062 ( .Y(T7062_Y), .B1(T12399_Y), .B0(T5243_Q),     .A1(T12425_Y), .A0(T289_Q));
KC_AOI22_X1 T7061 ( .Y(T7061_Y), .B1(T12423_Y), .B0(T5242_Q),     .A1(T12407_Y), .A0(T5562_Q));
KC_AOI22_X1 T6606 ( .Y(T6606_Y), .B1(T12409_Y), .B0(T167_Q),     .A1(T12408_Y), .A0(T5251_Q));
KC_AOI22_X1 T6600 ( .Y(T6600_Y), .B1(T8384_Y), .B0(T5559_Q),     .A1(T7364_Y), .A0(T164_Q));
KC_AOI22_X1 T6599 ( .Y(T6599_Y), .B1(T6828_Y), .B0(T5251_Q),     .A1(T6818_Y), .A0(T173_Q));
KC_AOI22_X1 T7313 ( .Y(T7313_Y), .B1(T7364_Y), .B0(T171_Q),     .A1(T8384_Y), .A0(T5263_Q));
KC_AOI22_X1 T7312 ( .Y(T7312_Y), .B1(T6801_Y), .B0(T169_Q),     .A1(T11864_Y), .A0(T5255_Q));
KC_AOI22_X1 T7309 ( .Y(T7309_Y), .B1(T15311_Y), .B0(T180_Q),     .A1(T15737_Y), .A0(T323_Q));
KC_AOI22_X1 T7308 ( .Y(T7308_Y), .B1(T12399_Y), .B0(T151_Q),     .A1(T12425_Y), .A0(T180_Q));
KC_AOI22_X1 T7290 ( .Y(T7290_Y), .B1(T6818_Y), .B0(T172_Q),     .A1(T6828_Y), .A0(T174_Q));
KC_AOI22_X1 T7288 ( .Y(T7288_Y), .B1(T15311_Y), .B0(T316_Q),     .A1(T15737_Y), .A0(T329_Q));
KC_AOI22_X1 T7274 ( .Y(T7274_Y), .B1(T15739_Y), .B0(T177_Q),     .A1(T8389_Y), .A0(T326_Q));
KC_AOI22_X1 T7273 ( .Y(T7273_Y), .B1(T12399_Y), .B0(T169_Q),     .A1(T12425_Y), .A0(T316_Q));
KC_AOI22_X1 T7271 ( .Y(T7271_Y), .B1(T12423_Y), .B0(T171_Q),     .A1(T12407_Y), .A0(T172_Q));
KC_AOI22_X1 T7270 ( .Y(T7270_Y), .B1(T12409_Y), .B0(T5255_Q),     .A1(T12408_Y), .A0(T174_Q));
KC_AOI22_X1 T7269 ( .Y(T7269_Y), .B1(T12426_Y), .B0(T5263_Q),     .A1(T12424_Y), .A0(T329_Q));
KC_AOI22_X1 T7252 ( .Y(T7252_Y), .B1(T12409_Y), .B0(T5237_Q),     .A1(T12408_Y), .A0(T5564_Q));
KC_AOI22_X1 T7251 ( .Y(T7251_Y), .B1(T12426_Y), .B0(T5239_Q),     .A1(T12424_Y), .A0(T323_Q));
KC_AOI22_X1 T6721 ( .Y(T6721_Y), .B1(T12423_Y), .B0(T164_Q),     .A1(T12407_Y), .A0(T173_Q));
KC_AOI22_X1 T6719 ( .Y(T6719_Y), .B1(T6828_Y), .B0(T182_Q),     .A1(T6818_Y), .A0(T166_Q));
KC_AOI22_X1 T6674 ( .Y(T6674_Y), .B1(T15739_Y), .B0(T9355_Q),     .A1(T8389_Y), .A0(T362_Q));
KC_AOI22_X1 T7456 ( .Y(T7456_Y), .B1(T7364_Y), .B0(T5303_Q),     .A1(T8384_Y), .A0(T9350_Q));
KC_AOI22_X1 T7455 ( .Y(T7455_Y), .B1(T12423_Y), .B0(T5303_Q),     .A1(T12407_Y), .A0(T204_Q));
KC_AOI22_X1 T7454 ( .Y(T7454_Y), .B1(T7364_Y), .B0(T9354_Q),     .A1(T8384_Y), .A0(T9349_Q));
KC_AOI22_X1 T7432 ( .Y(T7432_Y), .B1(T6818_Y), .B0(T5278_Q),     .A1(T6828_Y), .A0(T9352_Q));
KC_AOI22_X1 T7431 ( .Y(T7431_Y), .B1(T6818_Y), .B0(T204_Q),     .A1(T6828_Y), .A0(T5281_Q));
KC_AOI22_X1 T7430 ( .Y(T7430_Y), .B1(T6801_Y), .B0(T9353_Q),     .A1(T6821_Y), .A0(T337_Q));
KC_AOI22_X1 T7425 ( .Y(T7425_Y), .B1(T12409_Y), .B0(T337_Q),     .A1(T12408_Y), .A0(T5281_Q));
KC_AOI22_X1 T7423 ( .Y(T7423_Y), .B1(T8389_Y), .B0(T344_Q),     .A1(T15739_Y), .A0(T189_Q));
KC_AOI22_X1 T7422 ( .Y(T7422_Y), .B1(T12426_Y), .B0(T335_Q),     .A1(T12424_Y), .A0(T343_Q));
KC_AOI22_X1 T7402 ( .Y(T7402_Y), .B1(T11864_Y), .B0(T5275_Q),     .A1(T6801_Y), .A0(T183_Q));
KC_AOI22_X1 T7401 ( .Y(T7401_Y), .B1(T12409_Y), .B0(T5275_Q),     .A1(T12408_Y), .A0(T182_Q));
KC_AOI22_X1 T7400 ( .Y(T7400_Y), .B1(T12423_Y), .B0(T191_Q),     .A1(T12407_Y), .A0(T166_Q));
KC_AOI22_X1 T7399 ( .Y(T7399_Y), .B1(T8384_Y), .B0(T335_Q),     .A1(T7364_Y), .A0(T191_Q));
KC_AOI22_X1 T7398 ( .Y(T7398_Y), .B1(T12399_Y), .B0(T183_Q),     .A1(T12425_Y), .A0(T190_Q));
KC_AOI22_X1 T7387 ( .Y(T7387_Y), .B1(T6801_Y), .B0(T184_Q),     .A1(T11864_Y), .A0(T5277_Q));
KC_AOI22_X1 T7380 ( .Y(T7380_Y), .B1(T12423_Y), .B0(T9354_Q),     .A1(T12407_Y), .A0(T5278_Q));
KC_AOI22_X1 T7379 ( .Y(T7379_Y), .B1(T12399_Y), .B0(T184_Q),     .A1(T12425_Y), .A0(T359_Q));
KC_AOI22_X1 T7377 ( .Y(T7377_Y), .B1(T12409_Y), .B0(T5277_Q),     .A1(T12408_Y), .A0(T9352_Q));
KC_AOI22_X1 T7376 ( .Y(T7376_Y), .B1(T12426_Y), .B0(T9349_Q),     .A1(T12424_Y), .A0(T5304_Q));
KC_AOI22_X1 T7694 ( .Y(T7694_Y), .B1(T7670_Y), .B0(T9375_Y),     .A1(T16319_Y), .A0(T16332_Y));
KC_AOI22_X1 T7693 ( .Y(T7693_Y), .B1(T7830_Y), .B0(T9384_Y),     .A1(T7672_Y), .A0(T918_Y));
KC_AOI22_X1 T7692 ( .Y(T7692_Y), .B1(T7576_Y), .B0(T918_Y),     .A1(T9384_Y), .A0(T8698_Y));
KC_AOI22_X1 T7691 ( .Y(T7691_Y), .B1(T797_Y), .B0(T16328_Y),     .A1(T7670_Y), .A0(T739_Y));
KC_AOI22_X1 T7690 ( .Y(T7690_Y), .B1(T7669_Y), .B0(T9381_Y),     .A1(T7564_Y), .A0(T16331_Y));
KC_AOI22_X1 T7689 ( .Y(T7689_Y), .B1(T16334_Y), .B0(T9381_Y),     .A1(T9375_Y), .A0(T7574_Y));
KC_AOI22_X1 T7674 ( .Y(T7674_Y), .B1(T9149_Y), .B0(T8777_Y),     .A1(T9333_Y), .A0(T350_Y));
KC_AOI22_X1 T7673 ( .Y(T7673_Y), .B1(T8143_Y), .B0(T8777_Y),     .A1(T9511_Y), .A0(T350_Y));
KC_AOI22_X1 T7672 ( .Y(T7672_Y), .B1(T8108_Y), .B0(T8777_Y),     .A1(T8649_Y), .A0(T350_Y));
KC_AOI22_X1 T7667 ( .Y(T7667_Y), .B1(T11186_Y), .B0(T8697_Y),     .A1(T11185_Y), .A0(T8741_Y));
KC_AOI22_X1 T7666 ( .Y(T7666_Y), .B1(T8742_Y), .B0(T8136_Y),     .A1(T11207_Y), .A0(T8741_Y));
KC_AOI22_X1 T7665 ( .Y(T7665_Y), .B1(T11213_Y), .B0(T8697_Y),     .A1(T11206_Y), .A0(T8741_Y));
KC_AOI22_X1 T7664 ( .Y(T7664_Y), .B1(T11185_Y), .B0(T8697_Y),     .A1(T11213_Y), .A0(T8741_Y));
KC_AOI22_X1 T7663 ( .Y(T7663_Y), .B1(T8704_Y), .B0(T8697_Y),     .A1(T11186_Y), .A0(T8741_Y));
KC_AOI22_X1 T7628 ( .Y(T7628_Y), .B1(T8107_Y), .B0(T8777_Y),     .A1(T8607_Y), .A0(T350_Y));
KC_AOI22_X1 T7572 ( .Y(T7572_Y), .B1(T7578_Y), .B0(T16328_Y),     .A1(T8753_Y), .A0(T9384_Y));
KC_AOI22_X1 T7571 ( .Y(T7571_Y), .B1(T12607_Y), .B0(T9384_Y),     .A1(T642_Y), .A0(T739_Y));
KC_AOI22_X1 T7570 ( .Y(T7570_Y), .B1(T9143_Y), .B0(T8777_Y),     .A1(T9344_Y), .A0(T382_Y));
KC_AOI22_X1 T7569 ( .Y(T7569_Y), .B1(T9020_Y), .B0(T8777_Y),     .A1(T8606_Y), .A0(T382_Y));
KC_AOI22_X1 T7568 ( .Y(T7568_Y), .B1(T9389_Y), .B0(T642_Y),     .A1(T7669_Y), .A0(T739_Y));
KC_AOI22_X1 T16361 ( .Y(T16361_Y), .B1(T7910_Y), .B0(T8950_Y),     .A1(T7905_Y), .A0(T1334_Y));
KC_AOI22_X1 T16360 ( .Y(T16360_Y), .B1(T970_Y), .B0(T8950_Y),     .A1(T8948_Y), .A0(T16390_Y));
KC_AOI22_X1 T16321 ( .Y(T16321_Y), .B1(T7628_Y), .B0(T16325_Y),     .A1(T7673_Y), .A0(T16331_Y));
KC_AOI22_X1 T12450 ( .Y(T12450_Y), .B1(T9019_Y), .B0(T8865_Y),     .A1(T8669_Y), .A0(T371_Y));
KC_AOI22_X1 T7906 ( .Y(T7906_Y), .B1(T231_Y), .B0(T8865_Y),     .A1(T8669_Y), .A0(T371_Y));
KC_AOI22_X1 T7904 ( .Y(T7904_Y), .B1(T9066_Y), .B0(T8865_Y),     .A1(T8710_Y), .A0(T371_Y));
KC_AOI22_X1 T7903 ( .Y(T7903_Y), .B1(T9018_Y), .B0(T8865_Y),     .A1(T8648_Y), .A0(T371_Y));
KC_AOI22_X1 T7902 ( .Y(T7902_Y), .B1(T9148_Y), .B0(T8865_Y),     .A1(T8635_Y), .A0(T371_Y));
KC_AOI22_X1 T7873 ( .Y(T7873_Y), .B1(T11896_Y), .B0(T8812_Y),     .A1(T11897_Y), .A0(T8868_Y));
KC_AOI22_X1 T7872 ( .Y(T7872_Y), .B1(T15452_Y), .B0(T15354_Y),     .A1(T7677_Y), .A0(T8838_Y));
KC_AOI22_X1 T7862 ( .Y(T7862_Y), .B1(T11897_Y), .B0(T8812_Y),     .A1(T11265_Y), .A0(T8868_Y));
KC_AOI22_X1 T7861 ( .Y(T7861_Y), .B1(T8951_Y), .B0(T8812_Y),     .A1(T11895_Y), .A0(T8868_Y));
KC_AOI22_X1 T7858 ( .Y(T7858_Y), .B1(T9101_Y), .B0(T8865_Y),     .A1(T8605_Y), .A0(T350_Y));
KC_AOI22_X1 T7857 ( .Y(T7857_Y), .B1(T9017_Y), .B0(T8865_Y),     .A1(T8666_Y), .A0(T350_Y));
KC_AOI22_X1 T7856 ( .Y(T7856_Y), .B1(T9068_Y), .B0(T8865_Y),     .A1(T8646_Y), .A0(T371_Y));
KC_AOI22_X1 T7855 ( .Y(T7855_Y), .B1(T11895_Y), .B0(T8812_Y),     .A1(T11896_Y), .A0(T8868_Y));
KC_AOI22_X1 T7829 ( .Y(T7829_Y), .B1(T15452_Y), .B0(T7677_Y),     .A1(T15354_Y), .A0(T8782_Y));
KC_AOI22_X1 T8135 ( .Y(T8135_Y), .B1(T9020_Y), .B0(T9441_Y),     .A1(T5244_Y), .A0(T10069_Y));
KC_AOI22_X1 T8132 ( .Y(T8132_Y), .B1(T8108_Y), .B0(T9441_Y),     .A1(T8645_Y), .A0(T10069_Y));
KC_AOI22_X1 T8105 ( .Y(T8105_Y), .B1(T7858_Y), .B0(T1286_Y),     .A1(T7856_Y), .A0(T1334_Y));
KC_AOI22_X1 T8085 ( .Y(T8085_Y), .B1(T1286_Y), .B0(T16390_Y),     .A1(T7902_Y), .A0(T1272_Y));
KC_AOI22_X1 T8084 ( .Y(T8084_Y), .B1(T8099_Y), .B0(T1321_Y),     .A1(T1225_Y), .A0(T1286_Y));
KC_AOI22_X1 T8075 ( .Y(T8075_Y), .B1(T8148_Y), .B0(T8949_Y),     .A1(T7903_Y), .A0(T1266_Y));
KC_AOI22_X1 T8074 ( .Y(T8074_Y), .B1(T1287_Y), .B0(T1278_Y),     .A1(T7918_Y), .A0(T1284_Y));
KC_AOI22_X1 T8054 ( .Y(T8054_Y), .B1(T7918_Y), .B0(T8948_Y),     .A1(T1225_Y), .A0(T1213_Y));
KC_AOI22_X1 T8052 ( .Y(T8052_Y), .B1(T8077_Y), .B0(T1217_Y),     .A1(T7910_Y), .A0(T1284_Y));
KC_AOI22_X1 T8050 ( .Y(T8050_Y), .B1(T7863_Y), .B0(T1278_Y),     .A1(T8866_Y), .A0(T8949_Y));
KC_AOI22_X1 T8049 ( .Y(T8049_Y), .B1(T9421_Y), .B0(T8950_Y),     .A1(T7905_Y), .A0(T1266_Y));
KC_AOI22_X1 T8048 ( .Y(T8048_Y), .B1(T12886_Y), .B0(T8949_Y),     .A1(T1217_Y), .A0(T1284_Y));
KC_AOI22_X1 T8047 ( .Y(T8047_Y), .B1(T7909_Y), .B0(T1266_Y),     .A1(T8949_Y), .A0(T9424_Y));
KC_AOI22_X1 T219 ( .Y(T219_Y), .B1(T6597_Y), .B0(T5196_Q),     .A1(T6829_Y), .A0(T432_Q));
KC_AOI22_X1 T218 ( .Y(T218_Y), .B1(T6597_Y), .B0(T272_Q), .A1(T6829_Y),     .A0(T5193_Q));
KC_AOI22_X1 T6312 ( .Y(T6312_Y), .B1(T12425_Y), .B0(T5200_Q),     .A1(T12406_Y), .A0(T445_Q));
KC_AOI22_X1 T6311 ( .Y(T6311_Y), .B1(T6799_Y), .B0(T440_Q),     .A1(T15310_Y), .A0(T445_Q));
KC_AOI22_X1 T6310 ( .Y(T6310_Y), .B1(T6799_Y), .B0(T276_Q),     .A1(T15310_Y), .A0(T452_Q));
KC_AOI22_X1 T6309 ( .Y(T6309_Y), .B1(T600_Y), .B0(T5194_Q),     .A1(T12435_Y), .A0(T441_Q));
KC_AOI22_X1 T6296 ( .Y(T6296_Y), .B1(T12425_Y), .B0(T443_Q),     .A1(T12406_Y), .A0(T452_Q));
KC_AOI22_X1 T6291 ( .Y(T6291_Y), .B1(T600_Y), .B0(T432_Q),     .A1(T12435_Y), .A0(T435_Q));
KC_AOI22_X1 T6961 ( .Y(T6961_Y), .B1(T6818_Y), .B0(T283_Q),     .A1(T6828_Y), .A0(T5226_Q));
KC_AOI22_X1 T6956 ( .Y(T6956_Y), .B1(T15311_Y), .B0(T443_Q),     .A1(T15737_Y), .A0(T456_Q));
KC_AOI22_X1 T6925 ( .Y(T6925_Y), .B1(T12409_Y), .B0(T450_Q),     .A1(T12407_Y), .A0(T5204_Q));
KC_AOI22_X1 T6924 ( .Y(T6924_Y), .B1(T6801_Y), .B0(T439_Q),     .A1(T6821_Y), .A0(T450_Q));
KC_AOI22_X1 T6923 ( .Y(T6923_Y), .B1(T600_Y), .B0(T5193_Q),     .A1(T12435_Y), .A0(T274_Q));
KC_AOI22_X1 T6904 ( .Y(T6904_Y), .B1(T6597_Y), .B0(T438_Q),     .A1(T6829_Y), .A0(T5194_Q));
KC_AOI22_X1 T6903 ( .Y(T6903_Y), .B1(T6818_Y), .B0(T5204_Q),     .A1(T6828_Y), .A0(T446_Q));
KC_AOI22_X1 T6338 ( .Y(T6338_Y), .B1(T922_Y), .B0(T274_Q),     .A1(T16116_Y), .A0(T459_Q));
KC_AOI22_X1 T7118 ( .Y(T7118_Y), .B1(T12429_Y), .B0(T5241_Q),     .A1(T12427_Y), .A0(T459_Q));
KC_AOI22_X1 T7064 ( .Y(T7064_Y), .B1(T12405_Y), .B0(T281_Q),     .A1(T12406_Y), .A0(T460_Q));
KC_AOI22_X1 T7063 ( .Y(T7063_Y), .B1(T12399_Y), .B0(T277_Q),     .A1(T12405_Y), .A0(T272_Q));
KC_AOI22_X1 T7059 ( .Y(T7059_Y), .B1(T6799_Y), .B0(T160_Q),     .A1(T15310_Y), .A0(T460_Q));
KC_AOI22_X1 T7058 ( .Y(T7058_Y), .B1(T15734_Y), .B0(T434_Q),     .A1(T15735_Y), .A0(T440_Q));
KC_AOI22_X1 T7057 ( .Y(T7057_Y), .B1(T15734_Y), .B0(T294_Q),     .A1(T15735_Y), .A0(T273_Q));
KC_AOI22_X1 T6644 ( .Y(T6644_Y), .B1(T7650_Y), .B0(T714_Q),     .A1(T12429_Y), .A0(T326_Q));
KC_AOI22_X1 T6643 ( .Y(T6643_Y), .B1(T7650_Y), .B0(T517_Q),     .A1(T12429_Y), .A0(T4823_Q));
KC_AOI22_X1 T6642 ( .Y(T6642_Y), .B1(T7651_Y), .B0(T550_Q),     .A1(T15735_Y), .A0(T160_Q));
KC_AOI22_X1 T6641 ( .Y(T6641_Y), .B1(T922_Y), .B0(T5253_Q),     .A1(T16116_Y), .A0(T5254_Q));
KC_AOI22_X1 T6640 ( .Y(T6640_Y), .B1(T7651_Y), .B0(T741_Q),     .A1(T15735_Y), .A0(T170_Q));
KC_AOI22_X1 T6639 ( .Y(T6639_Y), .B1(T7651_Y), .B0(T4840_Q),     .A1(T15735_Y), .A0(T155_Q));
KC_AOI22_X1 T6617 ( .Y(T6617_Y), .B1(T7650_Y), .B0(T528_Q),     .A1(T12429_Y), .A0(T306_Q));
KC_AOI22_X1 T6616 ( .Y(T6616_Y), .B1(T15734_Y), .B0(T177_Q),     .A1(T12427_Y), .A0(T5254_Q));
KC_AOI22_X1 T6615 ( .Y(T6615_Y), .B1(T12405_Y), .B0(T664_Q),     .A1(T12406_Y), .A0(T5276_Q));
KC_AOI22_X1 T7304 ( .Y(T7304_Y), .B1(T15734_Y), .B0(T282_Q),     .A1(T12427_Y), .A0(T5265_Q));
KC_AOI22_X1 T7303 ( .Y(T7303_Y), .B1(T922_Y), .B0(T4810_Q),     .A1(T16116_Y), .A0(T5257_Q));
KC_AOI22_X1 T7302 ( .Y(T7302_Y), .B1(T6597_Y), .B0(T179_Q),     .A1(T6829_Y), .A0(T672_Q));
KC_AOI22_X1 T7301 ( .Y(T7301_Y), .B1(T600_Y), .B0(T672_Q),     .A1(T12435_Y), .A0(T4810_Q));
KC_AOI22_X1 T7285 ( .Y(T7285_Y), .B1(T12405_Y), .B0(T330_Q),     .A1(T12406_Y), .A0(T489_Q));
KC_AOI22_X1 T7284 ( .Y(T7284_Y), .B1(T6799_Y), .B0(T155_Q),     .A1(T15310_Y), .A0(T5260_Q));
KC_AOI22_X1 T7283 ( .Y(T7283_Y), .B1(T15734_Y), .B0(T154_Q),     .A1(T12427_Y), .A0(T5257_Q));
KC_AOI22_X1 T7266 ( .Y(T7266_Y), .B1(T6799_Y), .B0(T170_Q),     .A1(T15310_Y), .A0(T489_Q));
KC_AOI22_X1 T7265 ( .Y(T7265_Y), .B1(T600_Y), .B0(T5261_Q),     .A1(T12435_Y), .A0(T5253_Q));
KC_AOI22_X1 T7264 ( .Y(T7264_Y), .B1(T6597_Y), .B0(T330_Q),     .A1(T6829_Y), .A0(T5261_Q));
KC_AOI22_X1 T7247 ( .Y(T7247_Y), .B1(T12405_Y), .B0(T179_Q),     .A1(T12406_Y), .A0(T5260_Q));
KC_AOI22_X1 T7246 ( .Y(T7246_Y), .B1(T922_Y), .B0(T7085_Q),     .A1(T16116_Y), .A0(T5265_Q));
KC_AOI22_X1 T7245 ( .Y(T7245_Y), .B1(T6597_Y), .B0(T281_Q),     .A1(T6829_Y), .A0(T4835_Q));
KC_AOI22_X1 T6711 ( .Y(T6711_Y), .B1(T7650_Y), .B0(T713_Q),     .A1(T12429_Y), .A0(T319_Q));
KC_AOI22_X1 T6710 ( .Y(T6710_Y), .B1(T600_Y), .B0(T5560_Q),     .A1(T12435_Y), .A0(T4837_Q));
KC_AOI22_X1 T6666 ( .Y(T6666_Y), .B1(T15734_Y), .B0(T9355_Q),     .A1(T12427_Y), .A0(T519_Q));
KC_AOI22_X1 T6665 ( .Y(T6665_Y), .B1(T15734_Y), .B0(T189_Q),     .A1(T12427_Y), .A0(T525_Q));
KC_AOI22_X1 T6664 ( .Y(T6664_Y), .B1(T12426_Y), .B0(T9350_Q),     .A1(T12424_Y), .A0(T521_Q));
KC_AOI22_X1 T12410 ( .Y(T12410_Y), .B1(T15311_Y), .B0(T522_Q),     .A1(T15737_Y), .A0(T521_Q));
KC_AOI22_X1 T7448 ( .Y(T7448_Y), .B1(T6597_Y), .B0(T9339_Q),     .A1(T6829_Y), .A0(T5283_Q));
KC_AOI22_X1 T7447 ( .Y(T7447_Y), .B1(T12405_Y), .B0(T9339_Q),     .A1(T12406_Y), .A0(T699_Q));
KC_AOI22_X1 T7446 ( .Y(T7446_Y), .B1(T6799_Y), .B0(T9351_Q),     .A1(T15310_Y), .A0(T699_Q));
KC_AOI22_X1 T7445 ( .Y(T7445_Y), .B1(T600_Y), .B0(T5282_Q),     .A1(T12435_Y), .A0(T523_Q));
KC_AOI22_X1 T7420 ( .Y(T7420_Y), .B1(T15310_Y), .B0(T500_Q),     .A1(T6799_Y), .A0(T526_Q));
KC_AOI22_X1 T7419 ( .Y(T7419_Y), .B1(T12405_Y), .B0(T181_Q),     .A1(T12406_Y), .A0(T500_Q));
KC_AOI22_X1 T7395 ( .Y(T7395_Y), .B1(T7651_Y), .B0(T716_Q),     .A1(T15735_Y), .A0(T4799_Q));
KC_AOI22_X1 T7394 ( .Y(T7394_Y), .B1(T15734_Y), .B0(T165_Q),     .A1(T12427_Y), .A0(T681_Q));
KC_AOI22_X1 T7391 ( .Y(T7391_Y), .B1(T16116_Y), .B0(T681_Q),     .A1(T922_Y), .A0(T4837_Q));
KC_AOI22_X1 T7378 ( .Y(T7378_Y), .B1(T12399_Y), .B0(T9353_Q),     .A1(T12425_Y), .A0(T522_Q));
KC_AOI22_X1 T7373 ( .Y(T7373_Y), .B1(T12405_Y), .B0(T9338_Q),     .A1(T12406_Y), .A0(T501_Q));
KC_AOI22_X1 T7372 ( .Y(T7372_Y), .B1(T6597_Y), .B0(T9338_Q),     .A1(T6829_Y), .A0(T5282_Q));
KC_AOI22_X1 T7371 ( .Y(T7371_Y), .B1(T6799_Y), .B0(T360_Q),     .A1(T15310_Y), .A0(T501_Q));
KC_AOI22_X1 T7370 ( .Y(T7370_Y), .B1(T600_Y), .B0(T5279_Q),     .A1(T12435_Y), .A0(T341_Q));
KC_AOI22_X1 T7369 ( .Y(T7369_Y), .B1(T6829_Y), .B0(T5279_Q),     .A1(T6597_Y), .A0(T181_Q));
KC_AOI22_X1 T7659 ( .Y(T7659_Y), .B1(T7640_Y), .B0(T544_Q),     .A1(T7652_Y), .A0(T541_Q));
KC_AOI22_X1 T7658 ( .Y(T7658_Y), .B1(T9016_Y), .B0(T8777_Y),     .A1(T8663_Y), .A0(T382_Y));
KC_AOI22_X1 T7657 ( .Y(T7657_Y), .B1(T7652_Y), .B0(T5342_Q),     .A1(T7640_Y), .A0(T722_Q));
KC_AOI22_X1 T7656 ( .Y(T7656_Y), .B1(T7652_Y), .B0(T5350_Q),     .A1(T7640_Y), .A0(T5357_Q));
KC_AOI22_X1 T7655 ( .Y(T7655_Y), .B1(T7640_Y), .B0(T543_Q),     .A1(T7652_Y), .A0(T5346_Q));
KC_AOI22_X1 T7654 ( .Y(T7654_Y), .B1(T7640_Y), .B0(T5356_Q),     .A1(T7652_Y), .A0(T551_Q));
KC_AOI22_X1 T7622 ( .Y(T7622_Y), .B1(T7650_Y), .B0(T4827_Q),     .A1(T12429_Y), .A0(T344_Q));
KC_AOI22_X1 T7621 ( .Y(T7621_Y), .B1(T7650_Y), .B0(T701_Q),     .A1(T12429_Y), .A0(T524_Q));
KC_AOI22_X1 T7620 ( .Y(T7620_Y), .B1(T7650_Y), .B0(T512_Q),     .A1(T12429_Y), .A0(T362_Q));
KC_AOI22_X1 T7619 ( .Y(T7619_Y), .B1(T7651_Y), .B0(T529_Q),     .A1(T15735_Y), .A0(T526_Q));
KC_AOI22_X1 T7602 ( .Y(T7602_Y), .B1(T7651_Y), .B0(T530_Q),     .A1(T15735_Y), .A0(T360_Q));
KC_AOI22_X1 T7601 ( .Y(T7601_Y), .B1(T16116_Y), .B0(T525_Q),     .A1(T922_Y), .A0(T341_Q));
KC_AOI22_X1 T7600 ( .Y(T7600_Y), .B1(T7651_Y), .B0(T717_Q),     .A1(T15735_Y), .A0(T9351_Q));
KC_AOI22_X1 T7567 ( .Y(T7567_Y), .B1(T8087_Y), .B0(T8777_Y),     .A1(T8663_Y), .A0(T382_Y));
KC_AOI22_X1 T7564 ( .Y(T7564_Y), .B1(T8098_Y), .B0(T8777_Y),     .A1(T1143_Y), .A0(T382_Y));
KC_AOI22_X1 T16359 ( .Y(T16359_Y), .B1(T8087_Y), .B0(T9441_Y),     .A1(T482_Y), .A0(T10069_Y));
KC_AOI22_X1 T16358 ( .Y(T16358_Y), .B1(T554_Y), .B0(T8769_Y),     .A1(T16375_Y), .A0(T15660_Y));
KC_AOI22_X1 T16343 ( .Y(T16343_Y), .B1(T9371_Y), .B0(T554_Y),     .A1(T904_Y), .A0(T4840_Q));
KC_AOI22_X1 T16339 ( .Y(T16339_Y), .B1(T904_Y), .B0(T529_Q),     .A1(T9371_Y), .A0(T5537_Y));
KC_AOI22_X1 T16338 ( .Y(T16338_Y), .B1(T9371_Y), .B0(T2130_Y),     .A1(T904_Y), .A0(T530_Q));
KC_AOI22_X1 T16337 ( .Y(T16337_Y), .B1(T8735_Y), .B0(T776_Y),     .A1(T641_Y), .A0(T528_Q));
KC_AOI22_X1 T7905 ( .Y(T7905_Y), .B1(T240_Y), .B0(T8865_Y),     .A1(T8631_Y), .A0(T371_Y));
KC_AOI22_X1 T7898 ( .Y(T7898_Y), .B1(T9143_Y), .B0(T9441_Y),     .A1(T15733_Y), .A0(T10069_Y));
KC_AOI22_X1 T7897 ( .Y(T7897_Y), .B1(T5537_Y), .B0(T8769_Y),     .A1(T16375_Y), .A0(T975_Y));
KC_AOI22_X1 T7896 ( .Y(T7896_Y), .B1(T776_Y), .B0(T8769_Y),     .A1(T16375_Y), .A0(T15463_Y));
KC_AOI22_X1 T7895 ( .Y(T7895_Y), .B1(T9149_Y), .B0(T9441_Y),     .A1(T4833_Y), .A0(T10069_Y));
KC_AOI22_X1 T7894 ( .Y(T7894_Y), .B1(T8143_Y), .B0(T9441_Y),     .A1(T9347_Y), .A0(T10069_Y));
KC_AOI22_X1 T7890 ( .Y(T7890_Y), .B1(T2130_Y), .B0(T8769_Y),     .A1(T16375_Y), .A0(T1597_Y));
KC_AOI22_X1 T7871 ( .Y(T7871_Y), .B1(T8766_Y), .B0(T2130_Y),     .A1(T944_Y), .A0(T5357_Q));
KC_AOI22_X1 T7852 ( .Y(T7852_Y), .B1(T8766_Y), .B0(T776_Y),     .A1(T944_Y), .A0(T544_Q));
KC_AOI22_X1 T7849 ( .Y(T7849_Y), .B1(T8766_Y), .B0(T554_Y),     .A1(T944_Y), .A0(T543_Q));
KC_AOI22_X1 T7808 ( .Y(T7808_Y), .B1(T9371_Y), .B0(T776_Y),     .A1(T904_Y), .A0(T550_Q));
KC_AOI22_X1 T7807 ( .Y(T7807_Y), .B1(T8766_Y), .B0(T5537_Y),     .A1(T944_Y), .A0(T5356_Q));
KC_AOI22_X1 T1426 ( .Y(T1426_Y), .B1(T9012_Y), .B0(T1422_Y),     .A1(T390_Y), .A0(T1422_Y));
KC_AOI22_X1 T1425 ( .Y(T1425_Y), .B1(T9067_Y), .B0(T9441_Y),     .A1(T8681_Y), .A0(T10069_Y));
KC_AOI22_X1 T1420 ( .Y(T1420_Y), .B1(T9054_S), .B0(T1421_Y),     .A1(T8979_Y), .A0(T8864_Y));
KC_AOI22_X1 T8134 ( .Y(T8134_Y), .B1(T8136_Y), .B0(T9441_Y),     .A1(T8653_Y), .A0(T10069_Y));
KC_AOI22_X1 T8122 ( .Y(T8122_Y), .B1(T9016_Y), .B0(T9441_Y),     .A1(T8674_Y), .A0(T10069_Y));
KC_AOI22_X1 T8096 ( .Y(T8096_Y), .B1(T9116_Y), .B0(T9441_Y),     .A1(T9323_Y), .A0(T10069_Y));
KC_AOI22_X1 T8042 ( .Y(T8042_Y), .B1(T8038_Y), .B0(T8059_Y),     .A1(T8070_Y), .A0(T1205_Y));
KC_AOI22_X1 T4811 ( .Y(T4811_Y), .B1(T16515_Y), .B0(T1421_Y),     .A1(T592_Y), .A0(T9472_Q));
KC_AOI22_X1 T4809 ( .Y(T4809_Y), .B1(T9159_S), .B0(T1421_Y),     .A1(T597_Y), .A0(T1270_Q));
KC_AOI22_X1 T1840 ( .Y(T1840_Y), .B1(T9141_S), .B0(T1421_Y),     .A1(T12447_Y), .A0(T1264_Q));
KC_AOI22_X1 T1837 ( .Y(T1837_Y), .B1(T9142_S), .B0(T1421_Y),     .A1(T12447_Y), .A0(T1265_Q));
KC_AOI22_X1 T1836 ( .Y(T1836_Y), .B1(T9047_S), .B0(T1421_Y),     .A1(T12447_Y), .A0(T1271_Q));
KC_AOI22_X1 T1587 ( .Y(T1587_Y), .B1(T598_Y), .B0(T9061_Y),     .A1(T597_Y), .A0(T1250_Q));
KC_AOI22_X1 T1579 ( .Y(T1579_Y), .B1(T597_Y), .B0(T5404_Q),     .A1(T603_Y), .A0(T4842_Y));
KC_AOI22_X1 T6860 ( .Y(T6860_Y), .B1(T15352_Y), .B0(T5196_Q),     .A1(T13217_Y), .A0(T12374_Y));
KC_AOI22_X1 T6299 ( .Y(T6299_Y), .B1(T6304_Y), .B0(T276_Q),     .A1(T13269_Y), .A0(T6270_Y));
KC_AOI22_X1 T6294 ( .Y(T6294_Y), .B1(T12409_Y), .B0(T453_Q),     .A1(T12407_Y), .A0(T628_Q));
KC_AOI22_X1 T6292 ( .Y(T6292_Y), .B1(T12423_Y), .B0(T626_Q),     .A1(T12408_Y), .A0(T436_Q));
KC_AOI22_X1 T6285 ( .Y(T6285_Y), .B1(T12425_Y), .B0(T624_Q),     .A1(T12406_Y), .A0(T847_Q));
KC_AOI22_X1 T6282 ( .Y(T6282_Y), .B1(T12409_Y), .B0(T824_Q),     .A1(T12407_Y), .A0(T625_Q));
KC_AOI22_X1 T6281 ( .Y(T6281_Y), .B1(T12423_Y), .B0(T814_Q),     .A1(T12408_Y), .A0(T5229_Q));
KC_AOI22_X1 T6276 ( .Y(T6276_Y), .B1(T600_Y), .B0(T621_Q),     .A1(T12435_Y), .A0(T5206_Q));
KC_AOI22_X1 T6275 ( .Y(T6275_Y), .B1(T12409_Y), .B0(T812_Q),     .A1(T12407_Y), .A0(T630_Q));
KC_AOI22_X1 T6954 ( .Y(T6954_Y), .B1(T237_Y), .B0(T443_Q),     .A1(T13220_Y), .A0(T12385_Y));
KC_AOI22_X1 T6953 ( .Y(T6953_Y), .B1(T15311_Y), .B0(T5200_Q),     .A1(T15737_Y), .A0(T5223_Q));
KC_AOI22_X1 T6948 ( .Y(T6948_Y), .B1(T6818_Y), .B0(T625_Q),     .A1(T6828_Y), .A0(T815_Q));
KC_AOI22_X1 T6947 ( .Y(T6947_Y), .B1(T15311_Y), .B0(T624_Q),     .A1(T15737_Y), .A0(T649_Q));
KC_AOI22_X1 T6946 ( .Y(T6946_Y), .B1(T6818_Y), .B0(T630_Q),     .A1(T6828_Y), .A0(T5229_Q));
KC_AOI22_X1 T6940 ( .Y(T6940_Y), .B1(T7364_Y), .B0(T626_Q),     .A1(T8384_Y), .A0(T449_Q));
KC_AOI22_X1 T6938 ( .Y(T6938_Y), .B1(T7364_Y), .B0(T814_Q),     .A1(T8384_Y), .A0(T817_Q));
KC_AOI22_X1 T6920 ( .Y(T6920_Y), .B1(T6801_Y), .B0(T5205_Q),     .A1(T6821_Y), .A0(T453_Q));
KC_AOI22_X1 T6916 ( .Y(T6916_Y), .B1(T246_Y), .B0(T626_Q),     .A1(T13219_Y), .A0(T12381_Y));
KC_AOI22_X1 T6902 ( .Y(T6902_Y), .B1(T6818_Y), .B0(T628_Q),     .A1(T6828_Y), .A0(T436_Q));
KC_AOI22_X1 T6901 ( .Y(T6901_Y), .B1(T15351_Y), .B0(T628_Q),     .A1(T13218_Y), .A0(T12378_Y));
KC_AOI22_X1 T6899 ( .Y(T6899_Y), .B1(T6597_Y), .B0(T5199_Q),     .A1(T6829_Y), .A0(T826_Q));
KC_AOI22_X1 T6898 ( .Y(T6898_Y), .B1(T6597_Y), .B0(T627_Q),     .A1(T6829_Y), .A0(T621_Q));
KC_AOI22_X1 T6337 ( .Y(T6337_Y), .B1(T922_Y), .B0(T435_Q),     .A1(T16116_Y), .A0(T4846_Q));
KC_AOI22_X1 T6336 ( .Y(T6336_Y), .B1(T922_Y), .B0(T441_Q),     .A1(T16116_Y), .A0(T4845_Q));
KC_AOI22_X1 T6329 ( .Y(T6329_Y), .B1(T6331_Y), .B0(T435_Q),     .A1(T13226_Y), .A0(T12392_Y));
KC_AOI22_X1 T7114 ( .Y(T7114_Y), .B1(T12429_Y), .B0(T657_Q),     .A1(T12427_Y), .A0(T4846_Q));
KC_AOI22_X1 T7110 ( .Y(T7110_Y), .B1(T600_Y), .B0(T826_Q),     .A1(T12435_Y), .A0(T811_Q));
KC_AOI22_X1 T7089 ( .Y(T7089_Y), .B1(T12429_Y), .B0(T834_Q),     .A1(T12427_Y), .A0(T838_Q));
KC_AOI22_X1 T7081 ( .Y(T7081_Y), .B1(T12429_Y), .B0(T5240_Q),     .A1(T12427_Y), .A0(T4845_Q));
KC_AOI22_X1 T7080 ( .Y(T7080_Y), .B1(T324_Y), .B0(T5198_Q),     .A1(T13221_Y), .A0(T12394_Y));
KC_AOI22_X1 T7079 ( .Y(T7079_Y), .B1(T15739_Y), .B0(T5198_Q),     .A1(T8389_Y), .A0(T657_Q));
KC_AOI22_X1 T7076 ( .Y(T7076_Y), .B1(T12429_Y), .B0(T843_Q),     .A1(T12427_Y), .A0(T653_Q));
KC_AOI22_X1 T7055 ( .Y(T7055_Y), .B1(T15734_Y), .B0(T5198_Q),     .A1(T15735_Y), .A0(T276_Q));
KC_AOI22_X1 T7054 ( .Y(T7054_Y), .B1(T12426_Y), .B0(T5227_Q),     .A1(T12424_Y), .A0(T5223_Q));
KC_AOI22_X1 T7053 ( .Y(T7053_Y), .B1(T12426_Y), .B0(T449_Q),     .A1(T12424_Y), .A0(T456_Q));
KC_AOI22_X1 T7048 ( .Y(T7048_Y), .B1(T12426_Y), .B0(T823_Q),     .A1(T12424_Y), .A0(T820_Q));
KC_AOI22_X1 T7047 ( .Y(T7047_Y), .B1(T12426_Y), .B0(T817_Q),     .A1(T12424_Y), .A0(T649_Q));
KC_AOI22_X1 T7046 ( .Y(T7046_Y), .B1(T12423_Y), .B0(T816_Q),     .A1(T12408_Y), .A0(T815_Q));
KC_AOI22_X1 T7044 ( .Y(T7044_Y), .B1(T12425_Y), .B0(T793_Q),     .A1(T12406_Y), .A0(T848_Q));
KC_AOI22_X1 T6624 ( .Y(T6624_Y), .B1(T12425_Y), .B0(T665_Q),     .A1(T12406_Y), .A0(T6486_Q));
KC_AOI22_X1 T6623 ( .Y(T6623_Y), .B1(T12423_Y), .B0(T668_Q),     .A1(T12408_Y), .A0(T5264_Q));
KC_AOI22_X1 T6622 ( .Y(T6622_Y), .B1(T12399_Y), .B0(T666_Q),     .A1(T12405_Y), .A0(T663_Q));
KC_AOI22_X1 T7296 ( .Y(T7296_Y), .B1(T12429_Y), .B0(T5258_Q),     .A1(T12427_Y), .A0(T828_Q));
KC_AOI22_X1 T7294 ( .Y(T7294_Y), .B1(T15734_Y), .B0(T676_Q),     .A1(T15735_Y), .A0(T671_Q));
KC_AOI22_X1 T7293 ( .Y(T7293_Y), .B1(T12425_Y), .B0(T670_Q),     .A1(T12406_Y), .A0(T4854_Q));
KC_AOI22_X1 T7277 ( .Y(T7277_Y), .B1(T12426_Y), .B0(T861_Q),     .A1(T12424_Y), .A0(T5259_Q));
KC_AOI22_X1 T7239 ( .Y(T7239_Y), .B1(T12409_Y), .B0(T5565_Q),     .A1(T12407_Y), .A0(T677_Q));
KC_AOI22_X1 T6702 ( .Y(T6702_Y), .B1(T15734_Y), .B0(T694_Q),     .A1(T15735_Y), .A0(T680_Q));
KC_AOI22_X1 T6698 ( .Y(T6698_Y), .B1(T12426_Y), .B0(T863_Q),     .A1(T12424_Y), .A0(T865_Q));
KC_AOI22_X1 T6655 ( .Y(T6655_Y), .B1(T600_Y), .B0(T1040_Q),     .A1(T12435_Y), .A0(T711_Q));
KC_AOI22_X1 T6654 ( .Y(T6654_Y), .B1(T15734_Y), .B0(T710_Q),     .A1(T15735_Y), .A0(T695_Q));
KC_AOI22_X1 T6653 ( .Y(T6653_Y), .B1(T12423_Y), .B0(T5300_Q),     .A1(T12408_Y), .A0(T1041_Q));
KC_AOI22_X1 T7440 ( .Y(T7440_Y), .B1(T12409_Y), .B0(T1045_Q),     .A1(T12407_Y), .A0(T9340_Q));
KC_AOI22_X1 T7439 ( .Y(T7439_Y), .B1(T12407_Y), .B0(T697_Q),     .A1(T12409_Y), .A0(T1048_Q));
KC_AOI22_X1 T7438 ( .Y(T7438_Y), .B1(T12435_Y), .B0(T690_Q),     .A1(T600_Y), .A0(T1037_Q));
KC_AOI22_X1 T7368 ( .Y(T7368_Y), .B1(T12399_Y), .B0(T689_Q),     .A1(T12405_Y), .A0(T7367_Q));
KC_AOI22_X1 T7362 ( .Y(T7362_Y), .B1(T12399_Y), .B0(T712_Q),     .A1(T12405_Y), .A0(T687_Q));
KC_AOI22_X1 T7361 ( .Y(T7361_Y), .B1(T12425_Y), .B0(T688_Q),     .A1(T12406_Y), .A0(T1044_Q));
KC_AOI22_X1 T7360 ( .Y(T7360_Y), .B1(T15734_Y), .B0(T683_Q),     .A1(T15735_Y), .A0(T5280_Q));
KC_AOI22_X1 T7687 ( .Y(T7687_Y), .B1(T8735_Y), .B0(T2242_Y),     .A1(T641_Y), .A0(T713_Q));
KC_AOI22_X1 T7686 ( .Y(T7686_Y), .B1(T8735_Y), .B0(T841_Y),     .A1(T641_Y), .A0(T714_Q));
KC_AOI22_X1 T7649 ( .Y(T7649_Y), .B1(T7652_Y), .B0(T729_Q),     .A1(T7640_Y), .A0(T724_Q));
KC_AOI22_X1 T7595 ( .Y(T7595_Y), .B1(T12429_Y), .B0(T5301_Q),     .A1(T12427_Y), .A0(T5308_Q));
KC_AOI22_X1 T7594 ( .Y(T7594_Y), .B1(T12429_Y), .B0(T8714_Q),     .A1(T12427_Y), .A0(T709_Q));
KC_AOI22_X1 T7559 ( .Y(T7559_Y), .B1(T8735_Y), .B0(T2241_Y),     .A1(T641_Y), .A0(T701_Q));
KC_AOI22_X1 T16357 ( .Y(T16357_Y), .B1(T8086_Y), .B0(T9441_Y),     .A1(T661_Y), .A0(T10069_Y));
KC_AOI22_X1 T16356 ( .Y(T16356_Y), .B1(T996_Q), .B0(T8855_Y),     .A1(T1156_Q), .A0(T723_Y));
KC_AOI22_X1 T16355 ( .Y(T16355_Y), .B1(T8098_Y), .B0(T9441_Y),     .A1(T4839_Y), .A0(T10069_Y));
KC_AOI22_X1 T16354 ( .Y(T16354_Y), .B1(T773_Y), .B0(T8855_Y),     .A1(T1153_Q), .A0(T723_Y));
KC_AOI22_X1 T16346 ( .Y(T16346_Y), .B1(T9371_Y), .B0(T2241_Y),     .A1(T904_Y), .A0(T717_Q));
KC_AOI22_X1 T16345 ( .Y(T16345_Y), .B1(T9371_Y), .B0(T841_Y),     .A1(T904_Y), .A0(T741_Q));
KC_AOI22_X1 T7891 ( .Y(T7891_Y), .B1(T2242_Y), .B0(T8769_Y),     .A1(T16375_Y), .A0(T1709_Y));
KC_AOI22_X1 T7888 ( .Y(T7888_Y), .B1(T9458_Q), .B0(T8855_Y),     .A1(T1159_Q), .A0(T723_Y));
KC_AOI22_X1 T7886 ( .Y(T7886_Y), .B1(T723_Y), .B0(T963_Q),     .A1(T8855_Y), .A0(T759_Y));
KC_AOI22_X1 T7885 ( .Y(T7885_Y), .B1(T1152_Q), .B0(T8855_Y),     .A1(T16232_Q), .A0(T723_Y));
KC_AOI22_X1 T7884 ( .Y(T7884_Y), .B1(T9459_Q), .B0(T8855_Y),     .A1(T1160_Q), .A0(T723_Y));
KC_AOI22_X1 T7882 ( .Y(T7882_Y), .B1(T4844_Y), .B0(T8855_Y),     .A1(T999_Q), .A0(T723_Y));
KC_AOI22_X1 T7851 ( .Y(T7851_Y), .B1(T8769_Y), .B0(T2241_Y),     .A1(T16375_Y), .A0(T1578_Y));
KC_AOI22_X1 T7850 ( .Y(T7850_Y), .B1(T841_Y), .B0(T8769_Y),     .A1(T16375_Y), .A0(T1059_Y));
KC_AOI22_X1 T7806 ( .Y(T7806_Y), .B1(T8766_Y), .B0(T841_Y),     .A1(T944_Y), .A0(T722_Q));
KC_AOI22_X1 T7805 ( .Y(T7805_Y), .B1(T8766_Y), .B0(T2242_Y),     .A1(T944_Y), .A0(T725_Q));
KC_AOI22_X1 T7804 ( .Y(T7804_Y), .B1(T8766_Y), .B0(T2241_Y),     .A1(T944_Y), .A0(T724_Q));
KC_AOI22_X1 T1416 ( .Y(T1416_Y), .B1(T9489_Y), .B0(T9439_Y),     .A1(T9029_Y), .A0(T9440_Y));
KC_AOI22_X1 T1402 ( .Y(T1402_Y), .B1(T5379_Q), .B0(T9433_Y),     .A1(T963_Q), .A0(T9434_Y));
KC_AOI22_X1 T1400 ( .Y(T1400_Y), .B1(T752_Q), .B0(T9433_Y),     .A1(T765_Q), .A0(T9434_Y));
KC_AOI22_X1 T1399 ( .Y(T1399_Y), .B1(T8871_Y), .B0(T9442_Y),     .A1(T768_Q), .A0(T9434_Y));
KC_AOI22_X1 T12454 ( .Y(T12454_Y), .B1(T8107_Y), .B0(T9441_Y),     .A1(T678_Y), .A0(T10069_Y));
KC_AOI22_X1 T8114 ( .Y(T8114_Y), .B1(T5383_Q), .B0(T9433_Y),     .A1(T978_Q), .A0(T9434_Y));
KC_AOI22_X1 T8113 ( .Y(T8113_Y), .B1(T758_Y), .B0(T8996_Y),     .A1(T983_Q), .A0(T9002_Y));
KC_AOI22_X1 T8094 ( .Y(T8094_Y), .B1(T754_Q), .B0(T8996_Y),     .A1(T760_Q), .A0(T9002_Y));
KC_AOI22_X1 T8034 ( .Y(T8034_Y), .B1(T8944_Y), .B0(T1198_Y),     .A1(T8902_Y), .A0(T16388_Y));
KC_AOI22_X1 T8033 ( .Y(T8033_Y), .B1(T15084_Y), .B0(T9441_Y),     .A1(T655_Y), .A0(T10069_Y));
KC_AOI22_X1 T1838 ( .Y(T1838_Y), .B1(T7853_Y), .B0(T9011_Y),     .A1(T9471_Q), .A0(T9034_Y));
KC_AOI22_X1 T1741 ( .Y(T1741_Y), .B1(T7815_Y), .B0(T9011_Y),     .A1(T771_Q), .A0(T9034_Y));
KC_AOI22_X1 T1676 ( .Y(T1676_Y), .B1(T9460_Q), .B0(T9433_Y),     .A1(T1160_Q), .A0(T9434_Y));
KC_AOI22_X1 T1666 ( .Y(T1666_Y), .B1(T9461_Q), .B0(T9433_Y),     .A1(T1159_Q), .A0(T9434_Y));
KC_AOI22_X1 T1636 ( .Y(T1636_Y), .B1(T770_Q), .B0(T9433_Y),     .A1(T1153_Q), .A0(T9434_Y));
KC_AOI22_X1 T1635 ( .Y(T1635_Y), .B1(T780_Q), .B0(T9433_Y),     .A1(T16232_Q), .A0(T9434_Y));
KC_AOI22_X1 T1574 ( .Y(T1574_Y), .B1(T7854_Y), .B0(T9011_Y),     .A1(T769_Q), .A0(T9034_Y));
KC_AOI22_X1 T1568 ( .Y(T1568_Y), .B1(T7899_Y), .B0(T9011_Y),     .A1(T9470_Q), .A0(T9034_Y));
KC_AOI22_X1 T1562 ( .Y(T1562_Y), .B1(T4409_Y), .B0(T8996_Y),     .A1(T9457_Q), .A0(T9002_Y));
KC_AOI22_X1 T1561 ( .Y(T1561_Y), .B1(T4843_Q), .B0(T9433_Y),     .A1(T997_Q), .A0(T9434_Y));
KC_AOI22_X1 T1554 ( .Y(T1554_Y), .B1(T9178_Y), .B0(T10297_Y),     .A1(T1003_Q), .A0(T9033_Y));
KC_AOI22_X1 T6286 ( .Y(T6286_Y), .B1(T6801_Y), .B0(T790_Q),     .A1(T11864_Y), .A0(T812_Q));
KC_AOI22_X1 T6939 ( .Y(T6939_Y), .B1(T15311_Y), .B0(T793_Q),     .A1(T15737_Y), .A0(T820_Q));
KC_AOI22_X1 T6917 ( .Y(T6917_Y), .B1(T6801_Y), .B0(T822_Q),     .A1(T6821_Y), .A0(T824_Q));
KC_AOI22_X1 T6915 ( .Y(T6915_Y), .B1(T7364_Y), .B0(T816_Q),     .A1(T8384_Y), .A0(T823_Q));
KC_AOI22_X1 T7090 ( .Y(T7090_Y), .B1(T922_Y), .B0(T811_Q),     .A1(T16116_Y), .A0(T838_Q));
KC_AOI22_X1 T7078 ( .Y(T7078_Y), .B1(T15739_Y), .B0(T813_Q),     .A1(T8389_Y), .A0(T834_Q));
KC_AOI22_X1 T7077 ( .Y(T7077_Y), .B1(T6172_Y), .B0(T679_Q),     .A1(T315_Y), .A0(T5199_Q));
KC_AOI22_X1 T7075 ( .Y(T7075_Y), .B1(T15739_Y), .B0(T831_Q),     .A1(T8389_Y), .A0(T843_Q));
KC_AOI22_X1 T7045 ( .Y(T7045_Y), .B1(T6799_Y), .B0(T5195_Q),     .A1(T15310_Y), .A0(T847_Q));
KC_AOI22_X1 T7043 ( .Y(T7043_Y), .B1(T6799_Y), .B0(T825_Q),     .A1(T15310_Y), .A0(T848_Q));
KC_AOI22_X1 T6621 ( .Y(T6621_Y), .B1(T9299_Y), .B0(T668_Q),     .A1(T15772_Y), .A0(T715_Y));
KC_AOI22_X1 T6620 ( .Y(T6620_Y), .B1(T9302_Y), .B0(T694_Q),     .A1(T15780_Y), .A0(T715_Y));
KC_AOI22_X1 T6619 ( .Y(T6619_Y), .B1(T9502_Y), .B0(T666_Q),     .A1(T12904_Y), .A0(T715_Y));
KC_AOI22_X1 T7297 ( .Y(T7297_Y), .B1(T7364_Y), .B0(T4855_Q),     .A1(T8384_Y), .A0(T861_Q));
KC_AOI22_X1 T7292 ( .Y(T7292_Y), .B1(T6799_Y), .B0(T671_Q),     .A1(T15310_Y), .A0(T4854_Q));
KC_AOI22_X1 T7291 ( .Y(T7291_Y), .B1(T15739_Y), .B0(T676_Q),     .A1(T8389_Y), .A0(T5258_Q));
KC_AOI22_X1 T7276 ( .Y(T7276_Y), .B1(T15311_Y), .B0(T670_Q),     .A1(T15737_Y), .A0(T5259_Q));
KC_AOI22_X1 T7238 ( .Y(T7238_Y), .B1(T6801_Y), .B0(T829_Q),     .A1(T6821_Y), .A0(T5565_Q));
KC_AOI22_X1 T6648 ( .Y(T6648_Y), .B1(T9506_Y), .B0(T715_Y),     .A1(T9332_Y), .A0(T15223_Y));
KC_AOI22_X1 T6647 ( .Y(T6647_Y), .B1(T9328_Y), .B0(T6691_Y),     .A1(T542_Y), .A0(T1041_Q));
KC_AOI22_X1 T6646 ( .Y(T6646_Y), .B1(T16440_Y), .B0(T547_Y),     .A1(T15722_Y), .A0(T9334_Y));
KC_AOI22_X1 T7407 ( .Y(T7407_Y), .B1(T9507_Y), .B0(T715_Y),     .A1(T10345_Y), .A0(T15223_Y));
KC_AOI22_X1 T7355 ( .Y(T7355_Y), .B1(T9714_Y), .B0(T715_Y),     .A1(T7551_Y), .A0(T15223_Y));
KC_AOI22_X1 T7639 ( .Y(T7639_Y), .B1(T8731_Y), .B0(T727_Y),     .A1(T726_Y), .A0(T709_Q));
KC_AOI22_X1 T7629 ( .Y(T7629_Y), .B1(T7635_Y), .B0(T15223_Y),     .A1(T715_Y), .A0(T8719_Y));
KC_AOI22_X1 T7611 ( .Y(T7611_Y), .B1(T8718_Y), .B0(T669_Q),     .A1(T16090_Y), .A0(T715_Y));
KC_AOI22_X1 T7610 ( .Y(T7610_Y), .B1(T9505_Y), .B0(T715_Y),     .A1(T639_Y), .A0(T15223_Y));
KC_AOI22_X1 T7586 ( .Y(T7586_Y), .B1(T8709_Y), .B0(T9373_Y),     .A1(T700_Y), .A0(T8714_Q));
KC_AOI22_X1 T7585 ( .Y(T7585_Y), .B1(T9504_Y), .B0(T715_Y),     .A1(T15428_Y), .A0(T15223_Y));
KC_AOI22_X1 T7552 ( .Y(T7552_Y), .B1(T8687_Y), .B0(T9374_Y),     .A1(T15432_Y), .A0(T935_Q));
KC_AOI22_X1 T16353 ( .Y(T16353_Y), .B1(T8765_Y), .B0(T8764_Y),     .A1(T8756_Y), .A0(T902_Y));
KC_AOI22_X1 T16352 ( .Y(T16352_Y), .B1(T956_Y), .B0(T8765_Y),     .A1(T8756_Y), .A0(T8829_Y));
KC_AOI22_X1 T16351 ( .Y(T16351_Y), .B1(T8768_Y), .B0(T8764_Y),     .A1(T9365_Y), .A0(T902_Y));
KC_AOI22_X1 T7883 ( .Y(T7883_Y), .B1(T766_Y), .B0(T8855_Y),     .A1(T1158_Q), .A0(T723_Y));
KC_AOI22_X1 T7803 ( .Y(T7803_Y), .B1(T8768_Y), .B0(T956_Y),     .A1(T9365_Y), .A0(T8829_Y));
KC_AOI22_X1 T1415 ( .Y(T1415_Y), .B1(T5386_Q), .B0(T8996_Y),     .A1(T761_Q), .A0(T9002_Y));
KC_AOI22_X1 T1405 ( .Y(T1405_Y), .B1(T750_Q), .B0(T9433_Y),     .A1(T767_Q), .A0(T9434_Y));
KC_AOI22_X1 T1391 ( .Y(T1391_Y), .B1(T976_Q), .B0(T9433_Y),     .A1(T1151_Q), .A0(T9434_Y));
KC_AOI22_X1 T1653 ( .Y(T1653_Y), .B1(T5407_Q), .B0(T9433_Y),     .A1(T1156_Q), .A0(T9434_Y));
KC_AOI22_X1 T1631 ( .Y(T1631_Y), .B1(T1002_Q), .B0(T9433_Y),     .A1(T995_Q), .A0(T9434_Y));
KC_AOI22_X1 T1566 ( .Y(T1566_Y), .B1(T998_Q), .B0(T9433_Y),     .A1(T999_Q), .A0(T9434_Y));
KC_AOI22_X1 T1565 ( .Y(T1565_Y), .B1(T1004_Q), .B0(T9433_Y),     .A1(T5387_Q), .A0(T9434_Y));
KC_AOI22_X1 T1550 ( .Y(T1550_Y), .B1(T1013_Q), .B0(T8996_Y),     .A1(T5385_Q), .A0(T9002_Y));
KC_AOI22_X1 T10846 ( .Y(T10846_Y), .B1(T9579_Y), .B0(T13433_Q),     .A1(T14980_Y), .A0(T13334_Q));
KC_AOI22_X1 T10845 ( .Y(T10845_Y), .B1(T9579_Y), .B0(T13336_Q),     .A1(T14980_Y), .A0(T13333_Q));
KC_AOI22_X1 T10844 ( .Y(T10844_Y), .B1(T9579_Y), .B0(T13386_Q),     .A1(T14980_Y), .A0(T13382_Q));
KC_AOI22_X1 T10843 ( .Y(T10843_Y), .B1(T13357_Q), .B0(T9577_Y),     .A1(T13369_Q), .A0(T7337_Y));
KC_AOI22_X1 T10842 ( .Y(T10842_Y), .B1(T13338_Q), .B0(T9577_Y),     .A1(T13335_Q), .A0(T7337_Y));
KC_AOI22_X1 T6897 ( .Y(T6897_Y), .B1(T9579_Y), .B0(T13357_Q),     .A1(T14980_Y), .A0(T13369_Q));
KC_AOI22_X1 T6896 ( .Y(T6896_Y), .B1(T13386_Q), .B0(T9577_Y),     .A1(T13382_Q), .A0(T7337_Y));
KC_AOI22_X1 T6888 ( .Y(T6888_Y), .B1(T13354_Q), .B0(T9577_Y),     .A1(T13368_Q), .A0(T7337_Y));
KC_AOI22_X1 T6885 ( .Y(T6885_Y), .B1(T9579_Y), .B0(T13338_Q),     .A1(T14980_Y), .A0(T13335_Q));
KC_AOI22_X1 T6884 ( .Y(T6884_Y), .B1(T9579_Y), .B0(T13354_Q),     .A1(T14980_Y), .A0(T13368_Q));
KC_AOI22_X1 T10865 ( .Y(T10865_Y), .B1(T14717_Q), .B0(T9576_Y),     .A1(T14584_Q), .A0(T15237_Y));
KC_AOI22_X1 T10864 ( .Y(T10864_Y), .B1(T14586_Q), .B0(T9576_Y),     .A1(T13569_Q), .A0(T15237_Y));
KC_AOI22_X1 T10862 ( .Y(T10862_Y), .B1(T9585_Y), .B0(T13439_Q),     .A1(T15197_Y), .A0(T14713_Q));
KC_AOI22_X1 T10861 ( .Y(T10861_Y), .B1(T13441_Q), .B0(T9576_Y),     .A1(T14716_Q), .A0(T15237_Y));
KC_AOI22_X1 T10860 ( .Y(T10860_Y), .B1(T9585_Y), .B0(T13441_Q),     .A1(T15197_Y), .A0(T14716_Q));
KC_AOI22_X1 T10859 ( .Y(T10859_Y), .B1(T9585_Y), .B0(T14717_Q),     .A1(T15197_Y), .A0(T14584_Q));
KC_AOI22_X1 T10858 ( .Y(T10858_Y), .B1(T9585_Y), .B0(T14586_Q),     .A1(T15197_Y), .A0(T13569_Q));
KC_AOI22_X1 T7042 ( .Y(T7042_Y), .B1(T13433_Q), .B0(T9577_Y),     .A1(T13334_Q), .A0(T7337_Y));
KC_AOI22_X1 T7041 ( .Y(T7041_Y), .B1(T13336_Q), .B0(T9577_Y),     .A1(T13333_Q), .A0(T7337_Y));
KC_AOI22_X1 T7031 ( .Y(T7031_Y), .B1(T9573_Y), .B0(T14701_Q),     .A1(T9574_Y), .A0(T13437_Q));
KC_AOI22_X1 T7029 ( .Y(T7029_Y), .B1(T14701_Q), .B0(T6450_Y),     .A1(T13437_Q), .A0(T1336_Y));
KC_AOI22_X1 T7028 ( .Y(T7028_Y), .B1(T9573_Y), .B0(T13458_Q),     .A1(T9574_Y), .A0(T13472_Q));
KC_AOI22_X1 T7003 ( .Y(T7003_Y), .B1(T13458_Q), .B0(T6450_Y),     .A1(T13472_Q), .A0(T1336_Y));
KC_AOI22_X1 T10879 ( .Y(T10879_Y), .B1(T9573_Y), .B0(T13567_Q),     .A1(T9574_Y), .A0(T5753_Q));
KC_AOI22_X1 T10648 ( .Y(T10648_Y), .B1(T13436_Q), .B0(T9576_Y),     .A1(T13565_Q), .A0(T15237_Y));
KC_AOI22_X1 T7237 ( .Y(T7237_Y), .B1(T13568_Q), .B0(T6450_Y),     .A1(T1262_Q), .A0(T1336_Y));
KC_AOI22_X1 T7230 ( .Y(T7230_Y), .B1(T9575_Y), .B0(T13564_Q),     .A1(T9586_Y), .A0(T13616_Q));
KC_AOI22_X1 T7229 ( .Y(T7229_Y), .B1(T13564_Q), .B0(T9578_Y),     .A1(T13616_Q), .A0(T12073_Y));
KC_AOI22_X1 T7228 ( .Y(T7228_Y), .B1(T9585_Y), .B0(T13436_Q),     .A1(T15197_Y), .A0(T13565_Q));
KC_AOI22_X1 T7205 ( .Y(T7205_Y), .B1(T9573_Y), .B0(T13566_Q),     .A1(T9574_Y), .A0(T13594_Q));
KC_AOI22_X1 T7204 ( .Y(T7204_Y), .B1(T13567_Q), .B0(T6450_Y),     .A1(T5753_Q), .A0(T1336_Y));
KC_AOI22_X1 T7203 ( .Y(T7203_Y), .B1(T13566_Q), .B0(T6450_Y),     .A1(T13594_Q), .A0(T1336_Y));
KC_AOI22_X1 T7202 ( .Y(T7202_Y), .B1(T9575_Y), .B0(T5768_Q),     .A1(T9586_Y), .A0(T13743_Q));
KC_AOI22_X1 T7168 ( .Y(T7168_Y), .B1(T9573_Y), .B0(T13568_Q),     .A1(T9574_Y), .A0(T1262_Q));
KC_AOI22_X1 T7167 ( .Y(T7167_Y), .B1(T9575_Y), .B0(T13593_Q),     .A1(T9586_Y), .A0(T13592_Q));
KC_AOI22_X1 T7166 ( .Y(T7166_Y), .B1(T5768_Q), .B0(T9578_Y),     .A1(T13743_Q), .A0(T12073_Y));
KC_AOI22_X1 T7165 ( .Y(T7165_Y), .B1(T9575_Y), .B0(T14738_Q),     .A1(T9586_Y), .A0(T14736_Q));
KC_AOI22_X1 T7164 ( .Y(T7164_Y), .B1(T13578_Q), .B0(T6450_Y),     .A1(T13744_Q), .A0(T1336_Y));
KC_AOI22_X1 T7163 ( .Y(T7163_Y), .B1(T9573_Y), .B0(T13578_Q),     .A1(T9574_Y), .A0(T13744_Q));
KC_AOI22_X1 T7162 ( .Y(T7162_Y), .B1(T14738_Q), .B0(T9578_Y),     .A1(T14736_Q), .A0(T12073_Y));
KC_AOI22_X1 T7161 ( .Y(T7161_Y), .B1(T13593_Q), .B0(T9578_Y),     .A1(T13592_Q), .A0(T12073_Y));
KC_AOI22_X1 T7352 ( .Y(T7352_Y), .B1(T13706_Q), .B0(T12327_Y),     .A1(T13702_Q), .A0(T10788_Y));
KC_AOI22_X1 T7343 ( .Y(T7343_Y), .B1(T13707_Q), .B0(T12327_Y),     .A1(T13730_Q), .A0(T10788_Y));
KC_AOI22_X1 T7333 ( .Y(T7333_Y), .B1(T10419_Y), .B0(T13707_Q),     .A1(T1338_Y), .A0(T13730_Q));
KC_AOI22_X1 T7332 ( .Y(T7332_Y), .B1(T13708_Q), .B0(T12327_Y),     .A1(T13709_Q), .A0(T10788_Y));
KC_AOI22_X1 T7331 ( .Y(T7331_Y), .B1(T10419_Y), .B0(T13708_Q),     .A1(T1338_Y), .A0(T13709_Q));
KC_AOI22_X1 T5703 ( .Y(T5703_Y), .B1(T11918_Y), .B0(T9501_Y),     .A1(T15774_Y), .A0(T715_Y));
KC_AOI22_X1 T5702 ( .Y(T5702_Y), .B1(T11880_Y), .B0(T9500_Y),     .A1(T15778_Y), .A0(T715_Y));
KC_AOI22_X1 T5700 ( .Y(T5700_Y), .B1(T14753_Q), .B0(T10422_Y),     .A1(T14675_Q), .A0(T10367_Y));
KC_AOI22_X1 T5699 ( .Y(T5699_Y), .B1(T10420_Y), .B0(T14753_Q),     .A1(T10423_Y), .A0(T14675_Q));
KC_AOI22_X1 T5698 ( .Y(T5698_Y), .B1(T10419_Y), .B0(T14755_Q),     .A1(T1338_Y), .A0(T6745_Q));
KC_AOI22_X1 T5697 ( .Y(T5697_Y), .B1(T14755_Q), .B0(T12327_Y),     .A1(T6745_Q), .A0(T10788_Y));
KC_AOI22_X1 T10834 ( .Y(T10834_Y), .B1(T10420_Y), .B0(T14670_Q),     .A1(T10423_Y), .A0(T13842_Q));
KC_AOI22_X1 T10793 ( .Y(T10793_Y), .B1(T10419_Y), .B0(T14649_Q),     .A1(T1338_Y), .A0(T14652_Q));
KC_AOI22_X1 T10792 ( .Y(T10792_Y), .B1(T10419_Y), .B0(T13797_Q),     .A1(T1338_Y), .A0(T13868_Q));
KC_AOI22_X1 T7498 ( .Y(T7498_Y), .B1(T10419_Y), .B0(T13869_Q),     .A1(T1338_Y), .A0(T13826_Q));
KC_AOI22_X1 T7434 ( .Y(T7434_Y), .B1(T8677_Y), .B0(T497_Y),     .A1(T577_Y), .A0(T1046_Q));
KC_AOI22_X1 T7354 ( .Y(T7354_Y), .B1(T8659_Y), .B0(T549_Y),     .A1(T546_Y), .A0(T1040_Q));
KC_AOI22_X1 T8028 ( .Y(T8028_Y), .B1(T9900_Y), .B0(T15461_Y),     .A1(T9899_Y), .A0(T9891_Y));
KC_AOI22_X1 T8027 ( .Y(T8027_Y), .B1(T9900_Y), .B0(T1050_Y),     .A1(T9897_Y), .A0(T9891_Y));
KC_AOI22_X1 T8026 ( .Y(T8026_Y), .B1(T9900_Y), .B0(T8783_Y),     .A1(T9898_Y), .A0(T9891_Y));
KC_AOI22_X1 T7978 ( .Y(T7978_Y), .B1(T9900_Y), .B0(T8781_Y),     .A1(T9896_Y), .A0(T9891_Y));
KC_AOI22_X1 T10723 ( .Y(T10723_Y), .B1(T1007_Y), .B0(T9998_Y),     .A1(T12087_Y), .A0(T1246_Y));
KC_AOI22_X1 T10698 ( .Y(T10698_Y), .B1(T10028_Y), .B0(T1134_Y),     .A1(T980_Q), .A0(T140_Y));
KC_AOI22_X1 T10841 ( .Y(T10841_Y), .B1(T13356_Q), .B0(T9577_Y),     .A1(T13383_Q), .A0(T7337_Y));
KC_AOI22_X1 T6895 ( .Y(T6895_Y), .B1(T9579_Y), .B0(T13381_Q),     .A1(T14980_Y), .A0(T13363_Q));
KC_AOI22_X1 T6887 ( .Y(T6887_Y), .B1(T9579_Y), .B0(T13385_Q),     .A1(T14980_Y), .A0(T13366_Q));
KC_AOI22_X1 T6883 ( .Y(T6883_Y), .B1(T13385_Q), .B0(T9577_Y),     .A1(T13366_Q), .A0(T7337_Y));
KC_AOI22_X1 T6882 ( .Y(T6882_Y), .B1(T9579_Y), .B0(T13353_Q),     .A1(T14980_Y), .A0(T13384_Q));
KC_AOI22_X1 T6881 ( .Y(T6881_Y), .B1(T9579_Y), .B0(T13351_Q),     .A1(T14980_Y), .A0(T13379_Q));
KC_AOI22_X1 T6880 ( .Y(T6880_Y), .B1(T13353_Q), .B0(T9577_Y),     .A1(T13384_Q), .A0(T7337_Y));
KC_AOI22_X1 T6879 ( .Y(T6879_Y), .B1(T13355_Q), .B0(T9577_Y),     .A1(T13367_Q), .A0(T7337_Y));
KC_AOI22_X1 T6878 ( .Y(T6878_Y), .B1(T9579_Y), .B0(T13355_Q),     .A1(T14980_Y), .A0(T13367_Q));
KC_AOI22_X1 T6877 ( .Y(T6877_Y), .B1(T13381_Q), .B0(T9577_Y),     .A1(T13363_Q), .A0(T7337_Y));
KC_AOI22_X1 T6875 ( .Y(T6875_Y), .B1(T13351_Q), .B0(T9577_Y),     .A1(T13379_Q), .A0(T7337_Y));
KC_AOI22_X1 T10863 ( .Y(T10863_Y), .B1(T13439_Q), .B0(T9576_Y),     .A1(T14713_Q), .A0(T15237_Y));
KC_AOI22_X1 T10857 ( .Y(T10857_Y), .B1(T14711_Q), .B0(T9576_Y),     .A1(T13611_Q), .A0(T15237_Y));
KC_AOI22_X1 T10856 ( .Y(T10856_Y), .B1(T9585_Y), .B0(T14711_Q),     .A1(T15197_Y), .A0(T13611_Q));
KC_AOI22_X1 T10855 ( .Y(T10855_Y), .B1(T9585_Y), .B0(T13459_Q),     .A1(T15197_Y), .A0(T14700_Q));
KC_AOI22_X1 T10854 ( .Y(T10854_Y), .B1(T13459_Q), .B0(T9576_Y),     .A1(T14700_Q), .A0(T15237_Y));
KC_AOI22_X1 T7033 ( .Y(T7033_Y), .B1(T13469_Q), .B0(T9578_Y),     .A1(T13462_Q), .A0(T12073_Y));
KC_AOI22_X1 T7024 ( .Y(T7024_Y), .B1(T9573_Y), .B0(T13470_Q),     .A1(T9574_Y), .A0(T13471_Q));
KC_AOI22_X1 T7023 ( .Y(T7023_Y), .B1(T9573_Y), .B0(T14699_Q),     .A1(T9574_Y), .A0(T13483_Q));
KC_AOI22_X1 T7022 ( .Y(T7022_Y), .B1(T13460_Q), .B0(T9578_Y),     .A1(T13461_Q), .A0(T12073_Y));
KC_AOI22_X1 T7021 ( .Y(T7021_Y), .B1(T9575_Y), .B0(T13469_Q),     .A1(T9586_Y), .A0(T13462_Q));
KC_AOI22_X1 T7020 ( .Y(T7020_Y), .B1(T14699_Q), .B0(T6450_Y),     .A1(T13483_Q), .A0(T1336_Y));
KC_AOI22_X1 T7019 ( .Y(T7019_Y), .B1(T9575_Y), .B0(T13460_Q),     .A1(T9586_Y), .A0(T13461_Q));
KC_AOI22_X1 T7018 ( .Y(T7018_Y), .B1(T13470_Q), .B0(T6450_Y),     .A1(T13471_Q), .A0(T1336_Y));
KC_AOI22_X1 T7002 ( .Y(T7002_Y), .B1(T9575_Y), .B0(T13468_Q),     .A1(T9586_Y), .A0(T13457_Q));
KC_AOI22_X1 T7001 ( .Y(T7001_Y), .B1(T13468_Q), .B0(T9578_Y),     .A1(T13457_Q), .A0(T12073_Y));
KC_AOI22_X1 T7226 ( .Y(T7226_Y), .B1(T9573_Y), .B0(T14715_Q),     .A1(T9574_Y), .A0(T13589_Q));
KC_AOI22_X1 T7225 ( .Y(T7225_Y), .B1(T14715_Q), .B0(T6450_Y),     .A1(T13589_Q), .A0(T1336_Y));
KC_AOI22_X1 T7224 ( .Y(T7224_Y), .B1(T9573_Y), .B0(T14714_Q),     .A1(T9574_Y), .A0(T14735_Q));
KC_AOI22_X1 T7223 ( .Y(T7223_Y), .B1(T14714_Q), .B0(T6450_Y),     .A1(T14735_Q), .A0(T1336_Y));
KC_AOI22_X1 T7222 ( .Y(T7222_Y), .B1(T9573_Y), .B0(T14710_Q),     .A1(T9574_Y), .A0(T13588_Q));
KC_AOI22_X1 T7220 ( .Y(T7220_Y), .B1(T14710_Q), .B0(T6450_Y),     .A1(T13588_Q), .A0(T1336_Y));
KC_AOI22_X1 T7199 ( .Y(T7199_Y), .B1(T9575_Y), .B0(T13576_Q),     .A1(T9586_Y), .A0(T14737_Q));
KC_AOI22_X1 T7198 ( .Y(T7198_Y), .B1(T9575_Y), .B0(T13615_Q),     .A1(T9586_Y), .A0(T14731_Q));
KC_AOI22_X1 T7196 ( .Y(T7196_Y), .B1(T9585_Y), .B0(T13741_Q),     .A1(T15197_Y), .A0(T13742_Q));
KC_AOI22_X1 T7157 ( .Y(T7157_Y), .B1(T9575_Y), .B0(T13612_Q),     .A1(T9586_Y), .A0(T14732_Q));
KC_AOI22_X1 T7156 ( .Y(T7156_Y), .B1(T9573_Y), .B0(T13613_Q),     .A1(T9574_Y), .A0(T13577_Q));
KC_AOI22_X1 T7155 ( .Y(T7155_Y), .B1(T13615_Q), .B0(T9578_Y),     .A1(T14731_Q), .A0(T12073_Y));
KC_AOI22_X1 T7154 ( .Y(T7154_Y), .B1(T13613_Q), .B0(T6450_Y),     .A1(T13577_Q), .A0(T1336_Y));
KC_AOI22_X1 T7153 ( .Y(T7153_Y), .B1(T13612_Q), .B0(T9578_Y),     .A1(T14732_Q), .A0(T12073_Y));
KC_AOI22_X1 T7152 ( .Y(T7152_Y), .B1(T13576_Q), .B0(T9578_Y),     .A1(T14737_Q), .A0(T12073_Y));
KC_AOI22_X1 T7149 ( .Y(T7149_Y), .B1(T13741_Q), .B0(T9576_Y),     .A1(T13742_Q), .A0(T15237_Y));
KC_AOI22_X1 T7145 ( .Y(T7145_Y), .B1(T9575_Y), .B0(T13614_Q),     .A1(T9586_Y), .A0(T13590_Q));
KC_AOI22_X1 T7144 ( .Y(T7144_Y), .B1(T13614_Q), .B0(T9578_Y),     .A1(T13590_Q), .A0(T12073_Y));
KC_AOI22_X1 T7342 ( .Y(T7342_Y), .B1(T10368_Y), .B0(T13705_Q),     .A1(T10366_Y), .A0(T13726_Q));
KC_AOI22_X1 T7341 ( .Y(T7341_Y), .B1(T10368_Y), .B0(T13737_Q),     .A1(T10366_Y), .A0(T14751_Q));
KC_AOI22_X1 T7330 ( .Y(T7330_Y), .B1(T10419_Y), .B0(T13701_Q),     .A1(T1338_Y), .A0(T13699_Q));
KC_AOI22_X1 T7321 ( .Y(T7321_Y), .B1(T13701_Q), .B0(T12327_Y),     .A1(T13699_Q), .A0(T10788_Y));
KC_AOI22_X1 T5692 ( .Y(T5692_Y), .B1(T14674_Q), .B0(T10421_Y),     .A1(T13725_Q), .A0(T15194_Y));
KC_AOI22_X1 T5691 ( .Y(T5691_Y), .B1(T10420_Y), .B0(T13821_Q),     .A1(T10423_Y), .A0(T13839_Q));
KC_AOI22_X1 T5690 ( .Y(T5690_Y), .B1(T10418_Y), .B0(T14674_Q),     .A1(T15248_Y), .A0(T13725_Q));
KC_AOI22_X1 T5689 ( .Y(T5689_Y), .B1(T14754_Q), .B0(T1344_Y),     .A1(T13739_Q), .A0(T1343_Y));
KC_AOI22_X1 T5688 ( .Y(T5688_Y), .B1(T13737_Q), .B0(T1344_Y),     .A1(T14751_Q), .A0(T1343_Y));
KC_AOI22_X1 T5687 ( .Y(T5687_Y), .B1(T13705_Q), .B0(T1344_Y),     .A1(T13726_Q), .A0(T1343_Y));
KC_AOI22_X1 T5686 ( .Y(T5686_Y), .B1(T10368_Y), .B0(T13703_Q),     .A1(T10366_Y), .A0(T13704_Q));
KC_AOI22_X1 T5685 ( .Y(T5685_Y), .B1(T14671_Q), .B0(T10421_Y),     .A1(T13728_Q), .A0(T15194_Y));
KC_AOI22_X1 T5684 ( .Y(T5684_Y), .B1(T10418_Y), .B0(T14671_Q),     .A1(T15248_Y), .A0(T13728_Q));
KC_AOI22_X1 T5683 ( .Y(T5683_Y), .B1(T13703_Q), .B0(T1344_Y),     .A1(T13704_Q), .A0(T1343_Y));
KC_AOI22_X1 T5682 ( .Y(T5682_Y), .B1(T10368_Y), .B0(T14754_Q),     .A1(T10366_Y), .A0(T13739_Q));
KC_AOI22_X1 T5677 ( .Y(T5677_Y), .B1(T10420_Y), .B0(T13825_Q),     .A1(T10423_Y), .A0(T13823_Q));
KC_AOI22_X1 T10833 ( .Y(T10833_Y), .B1(T7234_Y), .B0(T15220_Y),     .A1(T5693_Y), .A0(T12086_Y));
KC_AOI22_X1 T10829 ( .Y(T10829_Y), .B1(T7207_Y), .B0(T15220_Y),     .A1(T5694_Y), .A0(T12086_Y));
KC_AOI22_X1 T7546 ( .Y(T7546_Y), .B1(T10418_Y), .B0(T13860_Q),     .A1(T15248_Y), .A0(T13861_Q));
KC_AOI22_X1 T7543 ( .Y(T7543_Y), .B1(T13860_Q), .B0(T10421_Y),     .A1(T13861_Q), .A0(T15194_Y));
KC_AOI22_X1 T7519 ( .Y(T7519_Y), .B1(T13830_Q), .B0(T10422_Y),     .A1(T13843_Q), .A0(T10367_Y));
KC_AOI22_X1 T7517 ( .Y(T7517_Y), .B1(T10418_Y), .B0(T13828_Q),     .A1(T15248_Y), .A0(T13829_Q));
KC_AOI22_X1 T7516 ( .Y(T7516_Y), .B1(T7034_Y), .B0(T15220_Y),     .A1(T7518_Y), .A0(T12086_Y));
KC_AOI22_X1 T7513 ( .Y(T7513_Y), .B1(T10418_Y), .B0(T14749_Q),     .A1(T15248_Y), .A0(T14667_Q));
KC_AOI22_X1 T7512 ( .Y(T7512_Y), .B1(T14749_Q), .B0(T10421_Y),     .A1(T14667_Q), .A0(T15194_Y));
KC_AOI22_X1 T7497 ( .Y(T7497_Y), .B1(T13869_Q), .B0(T12327_Y),     .A1(T13826_Q), .A0(T10788_Y));
KC_AOI22_X1 T7495 ( .Y(T7495_Y), .B1(T10368_Y), .B0(T13827_Q),     .A1(T10366_Y), .A0(T13863_Q));
KC_AOI22_X1 T7494 ( .Y(T7494_Y), .B1(T13827_Q), .B0(T1344_Y),     .A1(T13863_Q), .A0(T1343_Y));
KC_AOI22_X1 T7493 ( .Y(T7493_Y), .B1(T13828_Q), .B0(T10421_Y),     .A1(T13829_Q), .A0(T15194_Y));
KC_AOI22_X1 T7471 ( .Y(T7471_Y), .B1(T10420_Y), .B0(T13871_Q),     .A1(T10423_Y), .A0(T13867_Q));
KC_AOI22_X1 T7470 ( .Y(T7470_Y), .B1(T13871_Q), .B0(T10422_Y),     .A1(T13867_Q), .A0(T10367_Y));
KC_AOI22_X1 T7469 ( .Y(T7469_Y), .B1(T10420_Y), .B0(T13795_Q),     .A1(T10423_Y), .A0(T13796_Q));
KC_AOI22_X1 T7468 ( .Y(T7468_Y), .B1(T13795_Q), .B0(T10422_Y),     .A1(T13796_Q), .A0(T10367_Y));
KC_AOI22_X1 T7466 ( .Y(T7466_Y), .B1(T7201_Y), .B0(T15220_Y),     .A1(T7472_Y), .A0(T12086_Y));
KC_AOI22_X1 T7774 ( .Y(T7774_Y), .B1(T10418_Y), .B0(T14021_Q),     .A1(T15248_Y), .A0(T14020_Q));
KC_AOI22_X1 T7773 ( .Y(T7773_Y), .B1(T10418_Y), .B0(T13963_Q),     .A1(T15248_Y), .A0(T13964_Q));
KC_AOI22_X1 T7772 ( .Y(T7772_Y), .B1(T10368_Y), .B0(T14022_Q),     .A1(T10366_Y), .A0(T14018_Q));
KC_AOI22_X1 T7771 ( .Y(T7771_Y), .B1(T14651_Q), .B0(T1344_Y),     .A1(T14647_Q), .A0(T1343_Y));
KC_AOI22_X1 T7770 ( .Y(T7770_Y), .B1(T10368_Y), .B0(T14650_Q),     .A1(T10366_Y), .A0(T14644_Q));
KC_AOI22_X1 T7769 ( .Y(T7769_Y), .B1(T10420_Y), .B0(T13983_Q),     .A1(T10423_Y), .A0(T13971_Q));
KC_AOI22_X1 T7768 ( .Y(T7768_Y), .B1(T14003_Q), .B0(T12327_Y),     .A1(T14006_Q), .A0(T10788_Y));
KC_AOI22_X1 T7766 ( .Y(T7766_Y), .B1(T10418_Y), .B0(T13967_Q),     .A1(T15248_Y), .A0(T13968_Q));
KC_AOI22_X1 T7765 ( .Y(T7765_Y), .B1(T13963_Q), .B0(T10421_Y),     .A1(T13964_Q), .A0(T15194_Y));
KC_AOI22_X1 T7761 ( .Y(T7761_Y), .B1(T7158_Y), .B0(T15220_Y),     .A1(T7547_Y), .A0(T12086_Y));
KC_AOI22_X1 T7760 ( .Y(T7760_Y), .B1(T7200_Y), .B0(T15220_Y),     .A1(T7775_Y), .A0(T12086_Y));
KC_AOI22_X1 T7737 ( .Y(T7737_Y), .B1(T13967_Q), .B0(T10421_Y),     .A1(T13968_Q), .A0(T15194_Y));
KC_AOI22_X1 T7736 ( .Y(T7736_Y), .B1(T14005_Q), .B0(T10422_Y),     .A1(T14000_Q), .A0(T10367_Y));
KC_AOI22_X1 T7735 ( .Y(T7735_Y), .B1(T14022_Q), .B0(T1344_Y),     .A1(T14018_Q), .A0(T1343_Y));
KC_AOI22_X1 T7734 ( .Y(T7734_Y), .B1(T10420_Y), .B0(T14005_Q),     .A1(T10423_Y), .A0(T14000_Q));
KC_AOI22_X1 T7728 ( .Y(T7728_Y), .B1(T14021_Q), .B0(T10421_Y),     .A1(T14020_Q), .A0(T15194_Y));
KC_AOI22_X1 T7718 ( .Y(T7718_Y), .B1(T13983_Q), .B0(T10422_Y),     .A1(T13971_Q), .A0(T10367_Y));
KC_AOI22_X1 T10840 ( .Y(T10840_Y), .B1(T9577_Y), .B0(T13364_Q),     .A1(T13380_Q), .A0(T7337_Y));
KC_AOI22_X1 T10839 ( .Y(T10839_Y), .B1(T9579_Y), .B0(T13349_Q),     .A1(T14980_Y), .A0(T13348_Q));
KC_AOI22_X1 T10838 ( .Y(T10838_Y), .B1(T13378_Q), .B0(T9577_Y),     .A1(T13365_Q), .A0(T7337_Y));
KC_AOI22_X1 T10837 ( .Y(T10837_Y), .B1(T13362_Q), .B0(T9577_Y),     .A1(T13377_Q), .A0(T7337_Y));
KC_AOI22_X1 T6876 ( .Y(T6876_Y), .B1(T9579_Y), .B0(T13364_Q),     .A1(T14980_Y), .A0(T13380_Q));
KC_AOI22_X1 T6874 ( .Y(T6874_Y), .B1(T9579_Y), .B0(T13378_Q),     .A1(T14980_Y), .A0(T13365_Q));
KC_AOI22_X1 T6872 ( .Y(T6872_Y), .B1(T9579_Y), .B0(T13362_Q),     .A1(T14980_Y), .A0(T13377_Q));
KC_AOI22_X1 T10853 ( .Y(T10853_Y), .B1(T9585_Y), .B0(T14712_Q),     .A1(T15197_Y), .A0(T14709_Q));
KC_AOI22_X1 T10852 ( .Y(T10852_Y), .B1(T14712_Q), .B0(T9576_Y),     .A1(T14709_Q), .A0(T15237_Y));
KC_AOI22_X1 T10851 ( .Y(T10851_Y), .B1(T9573_Y), .B0(T14698_Q),     .A1(T9574_Y), .A0(T13484_Q));
KC_AOI22_X1 T10850 ( .Y(T10850_Y), .B1(T9585_Y), .B0(T14696_Q),     .A1(T15197_Y), .A0(T14692_Q));
KC_AOI22_X1 T10849 ( .Y(T10849_Y), .B1(T14696_Q), .B0(T9576_Y),     .A1(T14692_Q), .A0(T15237_Y));
KC_AOI22_X1 T7040 ( .Y(T7040_Y), .B1(T13349_Q), .B0(T9577_Y),     .A1(T13348_Q), .A0(T7337_Y));
KC_AOI22_X1 T7015 ( .Y(T7015_Y), .B1(T9573_Y), .B0(T14695_Q),     .A1(T9574_Y), .A0(T13482_Q));
KC_AOI22_X1 T7014 ( .Y(T7014_Y), .B1(T9573_Y), .B0(T13450_Q),     .A1(T9574_Y), .A0(T13449_Q));
KC_AOI22_X1 T7013 ( .Y(T7013_Y), .B1(T14698_Q), .B0(T6450_Y),     .A1(T13484_Q), .A0(T1336_Y));
KC_AOI22_X1 T7012 ( .Y(T7012_Y), .B1(T13450_Q), .B0(T6450_Y),     .A1(T13449_Q), .A0(T1336_Y));
KC_AOI22_X1 T7009 ( .Y(T7009_Y), .B1(T13454_Q), .B0(T9576_Y),     .A1(T13451_Q), .A0(T15237_Y));
KC_AOI22_X1 T7008 ( .Y(T7008_Y), .B1(T9585_Y), .B0(T13454_Q),     .A1(T15197_Y), .A0(T13451_Q));
KC_AOI22_X1 T7007 ( .Y(T7007_Y), .B1(T14695_Q), .B0(T6450_Y),     .A1(T13482_Q), .A0(T1336_Y));
KC_AOI22_X1 T7000 ( .Y(T7000_Y), .B1(T9575_Y), .B0(T13455_Q),     .A1(T9586_Y), .A0(T13500_Q));
KC_AOI22_X1 T6999 ( .Y(T6999_Y), .B1(T9575_Y), .B0(T13453_Q),     .A1(T9586_Y), .A0(T13456_Q));
KC_AOI22_X1 T6998 ( .Y(T6998_Y), .B1(T13455_Q), .B0(T9578_Y),     .A1(T13500_Q), .A0(T12073_Y));
KC_AOI22_X1 T6996 ( .Y(T6996_Y), .B1(T9575_Y), .B0(T13452_Q),     .A1(T9586_Y), .A0(T13481_Q));
KC_AOI22_X1 T6994 ( .Y(T6994_Y), .B1(T13453_Q), .B0(T9578_Y),     .A1(T13456_Q), .A0(T12073_Y));
KC_AOI22_X1 T10647 ( .Y(T10647_Y), .B1(T14734_Q), .B0(T9576_Y),     .A1(T14729_Q), .A0(T15237_Y));
KC_AOI22_X1 T7221 ( .Y(T7221_Y), .B1(T9573_Y), .B0(T13610_Q),     .A1(T9574_Y), .A0(T14697_Q));
KC_AOI22_X1 T7216 ( .Y(T7216_Y), .B1(T9575_Y), .B0(T14694_Q),     .A1(T9586_Y), .A0(T14706_Q));
KC_AOI22_X1 T7214 ( .Y(T7214_Y), .B1(T9576_Y), .B0(T14707_Q),     .A1(T15237_Y), .A0(T14708_Q));
KC_AOI22_X1 T7213 ( .Y(T7213_Y), .B1(T6450_Y), .B0(T13610_Q),     .A1(T1336_Y), .A0(T14697_Q));
KC_AOI22_X1 T7212 ( .Y(T7212_Y), .B1(T9585_Y), .B0(T14707_Q),     .A1(T15197_Y), .A0(T14708_Q));
KC_AOI22_X1 T7211 ( .Y(T7211_Y), .B1(T9578_Y), .B0(T14694_Q),     .A1(T12073_Y), .A0(T14706_Q));
KC_AOI22_X1 T7195 ( .Y(T7195_Y), .B1(T9585_Y), .B0(T13591_Q),     .A1(T15197_Y), .A0(T13587_Q));
KC_AOI22_X1 T7148 ( .Y(T7148_Y), .B1(T9585_Y), .B0(T14734_Q),     .A1(T15197_Y), .A0(T14729_Q));
KC_AOI22_X1 T7147 ( .Y(T7147_Y), .B1(T13591_Q), .B0(T9576_Y),     .A1(T13587_Q), .A0(T15237_Y));
KC_AOI22_X1 T7329 ( .Y(T7329_Y), .B1(T10419_Y), .B0(T13700_Q),     .A1(T1338_Y), .A0(T13698_Q));
KC_AOI22_X1 T7328 ( .Y(T7328_Y), .B1(T13700_Q), .B0(T12327_Y),     .A1(T13698_Q), .A0(T10788_Y));
KC_AOI22_X1 T7327 ( .Y(T7327_Y), .B1(T13694_Q), .B0(T12327_Y),     .A1(T13696_Q), .A0(T10788_Y));
KC_AOI22_X1 T7326 ( .Y(T7326_Y), .B1(T10419_Y), .B0(T13694_Q),     .A1(T1338_Y), .A0(T13696_Q));
KC_AOI22_X1 T7325 ( .Y(T7325_Y), .B1(T13697_Q), .B0(T12327_Y),     .A1(T13722_Q), .A0(T10788_Y));
KC_AOI22_X1 T7324 ( .Y(T7324_Y), .B1(T10419_Y), .B0(T13697_Q),     .A1(T1338_Y), .A0(T13722_Q));
KC_AOI22_X1 T5676 ( .Y(T5676_Y), .B1(T10368_Y), .B0(T13738_Q),     .A1(T10366_Y), .A0(T14752_Q));
KC_AOI22_X1 T5675 ( .Y(T5675_Y), .B1(T13738_Q), .B0(T1344_Y),     .A1(T14752_Q), .A0(T1343_Y));
KC_AOI22_X1 T6792 ( .Y(T6792_Y), .B1(T10368_Y), .B0(T14746_Q),     .A1(T10366_Y), .A0(T14747_Q));
KC_AOI22_X1 T10823 ( .Y(T10823_Y), .B1(T10420_Y), .B0(T13820_Q),     .A1(T10423_Y), .A0(T13817_Q));
KC_AOI22_X1 T10822 ( .Y(T10822_Y), .B1(T10418_Y), .B0(T13838_Q),     .A1(T15248_Y), .A0(T14668_Q));
KC_AOI22_X1 T10821 ( .Y(T10821_Y), .B1(T13820_Q), .B0(T10422_Y),     .A1(T13817_Q), .A0(T10367_Y));
KC_AOI22_X1 T10820 ( .Y(T10820_Y), .B1(T13824_Q), .B0(T10422_Y),     .A1(T13816_Q), .A0(T10367_Y));
KC_AOI22_X1 T10819 ( .Y(T10819_Y), .B1(T10420_Y), .B0(T13824_Q),     .A1(T10423_Y), .A0(T13816_Q));
KC_AOI22_X1 T10818 ( .Y(T10818_Y), .B1(T13838_Q), .B0(T10421_Y),     .A1(T14668_Q), .A0(T15194_Y));
KC_AOI22_X1 T10810 ( .Y(T10810_Y), .B1(T14746_Q), .B0(T1344_Y),     .A1(T14747_Q), .A0(T1343_Y));
KC_AOI22_X1 T10785 ( .Y(T10785_Y), .B1(T13998_Q), .B0(T12327_Y),     .A1(T14640_Q), .A0(T10788_Y));
KC_AOI22_X1 T10784 ( .Y(T10784_Y), .B1(T10419_Y), .B0(T14641_Q),     .A1(T1338_Y), .A0(T13999_Q));
KC_AOI22_X1 T7545 ( .Y(T7545_Y), .B1(T13859_Q), .B0(T10421_Y),     .A1(T13865_Q), .A0(T15194_Y));
KC_AOI22_X1 T7544 ( .Y(T7544_Y), .B1(T10418_Y), .B0(T13859_Q),     .A1(T15248_Y), .A0(T13865_Q));
KC_AOI22_X1 T7515 ( .Y(T7515_Y), .B1(T10418_Y), .B0(T13819_Q),     .A1(T15248_Y), .A0(T13836_Q));
KC_AOI22_X1 T7514 ( .Y(T7514_Y), .B1(T10418_Y), .B0(T13818_Q),     .A1(T15248_Y), .A0(T13837_Q));
KC_AOI22_X1 T7511 ( .Y(T7511_Y), .B1(T13818_Q), .B0(T10421_Y),     .A1(T13837_Q), .A0(T15194_Y));
KC_AOI22_X1 T7510 ( .Y(T7510_Y), .B1(T13819_Q), .B0(T10421_Y),     .A1(T13836_Q), .A0(T15194_Y));
KC_AOI22_X1 T7492 ( .Y(T7492_Y), .B1(T13864_Q), .B0(T1344_Y),     .A1(T13822_Q), .A0(T1343_Y));
KC_AOI22_X1 T7491 ( .Y(T7491_Y), .B1(T10368_Y), .B0(T13864_Q),     .A1(T10366_Y), .A0(T13822_Q));
KC_AOI22_X1 T7465 ( .Y(T7465_Y), .B1(T10420_Y), .B0(T13794_Q),     .A1(T10423_Y), .A0(T13862_Q));
KC_AOI22_X1 T7464 ( .Y(T7464_Y), .B1(T13794_Q), .B0(T10422_Y),     .A1(T13862_Q), .A0(T10367_Y));
KC_AOI22_X1 T7796 ( .Y(T7796_Y), .B1(T14014_Q), .B0(T10421_Y),     .A1(T13947_Q), .A0(T15194_Y));
KC_AOI22_X1 T7795 ( .Y(T7795_Y), .B1(T13948_Q), .B0(T10421_Y),     .A1(T13949_Q), .A0(T15194_Y));
KC_AOI22_X1 T7794 ( .Y(T7794_Y), .B1(T10418_Y), .B0(T13948_Q),     .A1(T15248_Y), .A0(T13949_Q));
KC_AOI22_X1 T7791 ( .Y(T7791_Y), .B1(T10421_Y), .B0(T14015_Q),     .A1(T15194_Y), .A0(T14017_Q));
KC_AOI22_X1 T7767 ( .Y(T7767_Y), .B1(T8022_Y), .B0(T15221_Y),     .A1(T10390_Y), .A0(T15220_Y));
KC_AOI22_X1 T7764 ( .Y(T7764_Y), .B1(T10419_Y), .B0(T14002_Q),     .A1(T1338_Y), .A0(T14645_Q));
KC_AOI22_X1 T7763 ( .Y(T7763_Y), .B1(T14002_Q), .B0(T12327_Y),     .A1(T14645_Q), .A0(T10788_Y));
KC_AOI22_X1 T7759 ( .Y(T7759_Y), .B1(T10419_Y), .B0(T13998_Q),     .A1(T1338_Y), .A0(T14640_Q));
KC_AOI22_X1 T7758 ( .Y(T7758_Y), .B1(T10419_Y), .B0(T14646_Q),     .A1(T1338_Y), .A0(T14639_Q));
KC_AOI22_X1 T7731 ( .Y(T7731_Y), .B1(T10420_Y), .B0(T13966_Q),     .A1(T10423_Y), .A0(T13969_Q));
KC_AOI22_X1 T7730 ( .Y(T7730_Y), .B1(T10420_Y), .B0(T13965_Q),     .A1(T10423_Y), .A0(T13970_Q));
KC_AOI22_X1 T7729 ( .Y(T7729_Y), .B1(T10368_Y), .B0(T14023_Q),     .A1(T10366_Y), .A0(T14019_Q));
KC_AOI22_X1 T7727 ( .Y(T7727_Y), .B1(T10368_Y), .B0(T14024_Q),     .A1(T10366_Y), .A0(T13944_Q));
KC_AOI22_X1 T7726 ( .Y(T7726_Y), .B1(T7989_Y), .B0(T15221_Y),     .A1(T7218_Y), .A0(T15220_Y));
KC_AOI22_X1 T7725 ( .Y(T7725_Y), .B1(T7943_Y), .B0(T15221_Y),     .A1(T7011_Y), .A0(T15220_Y));
KC_AOI22_X1 T7724 ( .Y(T7724_Y), .B1(T1344_Y), .B0(T14016_Q),     .A1(T1343_Y), .A0(T13945_Q));
KC_AOI22_X1 T7723 ( .Y(T7723_Y), .B1(T10368_Y), .B0(T14016_Q),     .A1(T10366_Y), .A0(T13945_Q));
KC_AOI22_X1 T7722 ( .Y(T7722_Y), .B1(T10420_Y), .B0(T13962_Q),     .A1(T10423_Y), .A0(T13961_Q));
KC_AOI22_X1 T7716 ( .Y(T7716_Y), .B1(T10418_Y), .B0(T14014_Q),     .A1(T15248_Y), .A0(T13947_Q));
KC_AOI22_X1 T7715 ( .Y(T7715_Y), .B1(T14023_Q), .B0(T1344_Y),     .A1(T14019_Q), .A0(T1343_Y));
KC_AOI22_X1 T7714 ( .Y(T7714_Y), .B1(T13966_Q), .B0(T10422_Y),     .A1(T13969_Q), .A0(T10367_Y));
KC_AOI22_X1 T7713 ( .Y(T7713_Y), .B1(T14024_Q), .B0(T1344_Y),     .A1(T13944_Q), .A0(T1343_Y));
KC_AOI22_X1 T7712 ( .Y(T7712_Y), .B1(T13965_Q), .B0(T10422_Y),     .A1(T13970_Q), .A0(T10367_Y));
KC_AOI22_X1 T7710 ( .Y(T7710_Y), .B1(T10418_Y), .B0(T14015_Q),     .A1(T15248_Y), .A0(T14017_Q));
KC_AOI22_X1 T7709 ( .Y(T7709_Y), .B1(T10422_Y), .B0(T13962_Q),     .A1(T10367_Y), .A0(T13961_Q));
KC_AOI22_X1 T7708 ( .Y(T7708_Y), .B1(T7996_Y), .B0(T15221_Y),     .A1(T7027_Y), .A0(T15220_Y));
KC_AOI22_X1 T10754 ( .Y(T10754_Y), .B1(T10306_Y), .B0(T14281_Q),     .A1(T10009_Y), .A0(T14605_Q));
KC_AOI22_X1 T10753 ( .Y(T10753_Y), .B1(T12094_Y), .B0(T14606_Q),     .A1(T8000_Y), .A0(T14109_Q));
KC_AOI22_X1 T10751 ( .Y(T10751_Y), .B1(T14606_Q), .B0(T12088_Y),     .A1(T14109_Q), .A0(T8011_Y));
KC_AOI22_X1 T8021 ( .Y(T8021_Y), .B1(T1584_Y), .B0(T14135_Q),     .A1(T1585_Y), .A0(T14619_Q));
KC_AOI22_X1 T8020 ( .Y(T8020_Y), .B1(T10306_Y), .B0(T14133_Q),     .A1(T10009_Y), .A0(T14111_Q));
KC_AOI22_X1 T8019 ( .Y(T8019_Y), .B1(T14623_Q), .B0(T1584_Y),     .A1(T14621_Q), .A0(T1585_Y));
KC_AOI22_X1 T8018 ( .Y(T8018_Y), .B1(T8862_Y), .B0(T14623_Q),     .A1(T9883_Y), .A0(T14621_Q));
KC_AOI22_X1 T8016 ( .Y(T8016_Y), .B1(T10033_Y), .B0(T14624_Q),     .A1(T15228_Y), .A0(T14618_Q));
KC_AOI22_X1 T8015 ( .Y(T8015_Y), .B1(T8017_Y), .B0(T14615_Q),     .A1(T10037_Y), .A0(T1484_Y));
KC_AOI22_X1 T7995 ( .Y(T7995_Y), .B1(T10306_Y), .B0(T14136_Q),     .A1(T10009_Y), .A0(T14112_Q));
KC_AOI22_X1 T7994 ( .Y(T7994_Y), .B1(T9892_Y), .B0(T14123_Q),     .A1(T9902_Y), .A0(T14134_Q));
KC_AOI22_X1 T7993 ( .Y(T7993_Y), .B1(T14136_Q), .B0(T9892_Y),     .A1(T14112_Q), .A0(T9902_Y));
KC_AOI22_X1 T7992 ( .Y(T7992_Y), .B1(T10306_Y), .B0(T14123_Q),     .A1(T10009_Y), .A0(T14134_Q));
KC_AOI22_X1 T7988 ( .Y(T7988_Y), .B1(T8862_Y), .B0(T14622_Q),     .A1(T9883_Y), .A0(T14132_Q));
KC_AOI22_X1 T7974 ( .Y(T7974_Y), .B1(T8862_Y), .B0(T14135_Q),     .A1(T9883_Y), .A0(T14619_Q));
KC_AOI22_X1 T7973 ( .Y(T7973_Y), .B1(T14622_Q), .B0(T1584_Y),     .A1(T14132_Q), .A0(T1585_Y));
KC_AOI22_X1 T7972 ( .Y(T7972_Y), .B1(T14133_Q), .B0(T9892_Y),     .A1(T14111_Q), .A0(T9902_Y));
KC_AOI22_X1 T7969 ( .Y(T7969_Y), .B1(T10033_Y), .B0(T14130_Q),     .A1(T15228_Y), .A0(T14131_Q));
KC_AOI22_X1 T7968 ( .Y(T7968_Y), .B1(T14624_Q), .B0(T9893_Y),     .A1(T14618_Q), .A0(T15229_Y));
KC_AOI22_X1 T7966 ( .Y(T7966_Y), .B1(T14130_Q), .B0(T9893_Y),     .A1(T14131_Q), .A0(T15229_Y));
KC_AOI22_X1 T7965 ( .Y(T7965_Y), .B1(T9893_Y), .B0(T14617_Q),     .A1(T15229_Y), .A0(T14620_Q));
KC_AOI22_X1 T7964 ( .Y(T7964_Y), .B1(T10033_Y), .B0(T14617_Q),     .A1(T15228_Y), .A0(T14620_Q));
KC_AOI22_X1 T7947 ( .Y(T7947_Y), .B1(T12094_Y), .B0(T15068_Q),     .A1(T8000_Y), .A0(T14121_Q));
KC_AOI22_X1 T7946 ( .Y(T7946_Y), .B1(T15068_Q), .B0(T12088_Y),     .A1(T14121_Q), .A0(T8011_Y));
KC_AOI22_X1 T7941 ( .Y(T7941_Y), .B1(T14108_Q), .B0(T9893_Y),     .A1(T14118_Q), .A0(T15229_Y));
KC_AOI22_X1 T7938 ( .Y(T7938_Y), .B1(T10033_Y), .B0(T14108_Q),     .A1(T15228_Y), .A0(T14118_Q));
KC_AOI22_X1 T7937 ( .Y(T7937_Y), .B1(T8862_Y), .B0(T14106_Q),     .A1(T9883_Y), .A0(T14120_Q));
KC_AOI22_X1 T7936 ( .Y(T7936_Y), .B1(T14106_Q), .B0(T1584_Y),     .A1(T14120_Q), .A0(T1585_Y));
KC_AOI22_X1 T10721 ( .Y(T10721_Y), .B1(T14281_Q), .B0(T9892_Y),     .A1(T14605_Q), .A0(T9902_Y));
KC_AOI22_X1 T10720 ( .Y(T10720_Y), .B1(T8862_Y), .B0(T14263_Q),     .A1(T9883_Y), .A0(T14279_Q));
KC_AOI22_X1 T10719 ( .Y(T10719_Y), .B1(T14263_Q), .B0(T1584_Y),     .A1(T14279_Q), .A0(T1585_Y));
KC_AOI22_X1 T10718 ( .Y(T10718_Y), .B1(T10033_Y), .B0(T14278_Q),     .A1(T15228_Y), .A0(T14603_Q));
KC_AOI22_X1 T10717 ( .Y(T10717_Y), .B1(T14278_Q), .B0(T9893_Y),     .A1(T14603_Q), .A0(T15229_Y));
KC_AOI22_X1 T10716 ( .Y(T10716_Y), .B1(T14280_Q), .B0(T12088_Y),     .A1(T14283_Q), .A0(T8011_Y));
KC_AOI22_X1 T10696 ( .Y(T10696_Y), .B1(T14262_Q), .B0(T9892_Y),     .A1(T14256_Q), .A0(T9902_Y));
KC_AOI22_X1 T10695 ( .Y(T10695_Y), .B1(T12094_Y), .B0(T14260_Q),     .A1(T8000_Y), .A0(T14240_Q));
KC_AOI22_X1 T10694 ( .Y(T10694_Y), .B1(T14257_Q), .B0(T9893_Y),     .A1(T14259_Q), .A0(T15229_Y));
KC_AOI22_X1 T10693 ( .Y(T10693_Y), .B1(T10033_Y), .B0(T14239_Q),     .A1(T15228_Y), .A0(T14238_Q));
KC_AOI22_X1 T10692 ( .Y(T10692_Y), .B1(T14260_Q), .B0(T12088_Y),     .A1(T14240_Q), .A0(T8011_Y));
KC_AOI22_X1 T10691 ( .Y(T10691_Y), .B1(T10306_Y), .B0(T14262_Q),     .A1(T10009_Y), .A0(T14256_Q));
KC_AOI22_X1 T10690 ( .Y(T10690_Y), .B1(T10033_Y), .B0(T14257_Q),     .A1(T15228_Y), .A0(T14259_Q));
KC_AOI22_X1 T10689 ( .Y(T10689_Y), .B1(T12094_Y), .B0(T14280_Q),     .A1(T8000_Y), .A0(T14283_Q));
KC_AOI22_X1 T10682 ( .Y(T10682_Y), .B1(T14261_Q), .B0(T9892_Y),     .A1(T14241_Q), .A0(T9902_Y));
KC_AOI22_X1 T10681 ( .Y(T10681_Y), .B1(T14239_Q), .B0(T9893_Y),     .A1(T14238_Q), .A0(T15229_Y));
KC_AOI22_X1 T10675 ( .Y(T10675_Y), .B1(T14231_Q), .B0(T9892_Y),     .A1(T14230_Q), .A0(T9902_Y));
KC_AOI22_X1 T10674 ( .Y(T10674_Y), .B1(T10306_Y), .B0(T14261_Q),     .A1(T10009_Y), .A0(T14241_Q));
KC_AOI22_X1 T10673 ( .Y(T10673_Y), .B1(T8862_Y), .B0(T14215_Q),     .A1(T9883_Y), .A0(T14214_Q));
KC_AOI22_X1 T10672 ( .Y(T10672_Y), .B1(T14229_Q), .B0(T1584_Y),     .A1(T14228_Q), .A0(T1585_Y));
KC_AOI22_X1 T10671 ( .Y(T10671_Y), .B1(T14215_Q), .B0(T1584_Y),     .A1(T14214_Q), .A0(T1585_Y));
KC_AOI22_X1 T10658 ( .Y(T10658_Y), .B1(T10306_Y), .B0(T14231_Q),     .A1(T10009_Y), .A0(T14230_Q));
KC_AOI22_X1 T10657 ( .Y(T10657_Y), .B1(T14597_Q), .B0(T12088_Y),     .A1(T14213_Q), .A0(T8011_Y));
KC_AOI22_X1 T10656 ( .Y(T10656_Y), .B1(T8862_Y), .B0(T14229_Q),     .A1(T9883_Y), .A0(T14228_Q));
KC_AOI22_X1 T10736 ( .Y(T10736_Y), .B1(T12094_Y), .B0(T14382_Q),     .A1(T8000_Y), .A0(T14387_Q));
KC_AOI22_X1 T10735 ( .Y(T10735_Y), .B1(T12088_Y), .B0(T14382_Q),     .A1(T14387_Q), .A0(T8011_Y));
KC_AOI22_X1 T10732 ( .Y(T10732_Y), .B1(T12094_Y), .B0(T14375_Q),     .A1(T8000_Y), .A0(T14381_Q));
KC_AOI22_X1 T1360 ( .Y(T1360_Y), .B1(T10122_Y), .B0(T10724_Y),     .A1(T1359_Y), .A0(T10122_Y));
KC_AOI22_X1 T7215 ( .Y(T7215_Y), .B1(T7217_Y), .B0(T13609_Q),     .A1(T7232_Y), .A0(T9642_Y));
KC_AOI22_X1 T7190 ( .Y(T7190_Y), .B1(T7133_Y), .B0(T13607_Q),     .A1(T10391_Y), .A0(T4937_Y));
KC_AOI22_X1 T7189 ( .Y(T7189_Y), .B1(T7134_Y), .B0(T13585_Q),     .A1(T7010_Y), .A0(T4937_Y));
KC_AOI22_X1 T7179 ( .Y(T7179_Y), .B1(T7180_Y), .B0(T14726_Q),     .A1(T7151_Y), .A0(T9642_Y));
KC_AOI22_X1 T7178 ( .Y(T7178_Y), .B1(T7181_Y), .B0(T14727_Q),     .A1(T7160_Y), .A0(T9642_Y));
KC_AOI22_X1 T7140 ( .Y(T7140_Y), .B1(T7193_Y), .B0(T14725_Q),     .A1(T7235_Y), .A0(T4937_Y));
KC_AOI22_X1 T7132 ( .Y(T7132_Y), .B1(T7138_Y), .B0(T13584_Q),     .A1(T7026_Y), .A0(T9642_Y));
KC_AOI22_X1 T7131 ( .Y(T7131_Y), .B1(T7135_Y), .B0(T13573_Q),     .A1(T7159_Y), .A0(T9642_Y));
KC_AOI22_X1 T7130 ( .Y(T7130_Y), .B1(T7137_Y), .B0(T13606_Q),     .A1(T7227_Y), .A0(T9642_Y));
KC_AOI22_X1 T7127 ( .Y(T7127_Y), .B1(T7136_Y), .B0(T14728_Q),     .A1(T6997_Y), .A0(T9642_Y));
KC_AOI22_X1 T7336 ( .Y(T7336_Y), .B1(T5672_Y), .B0(T13717_Q),     .A1(T7496_Y), .A0(T1484_Y));
KC_AOI22_X1 T7335 ( .Y(T7335_Y), .B1(T5670_Y), .B0(T13692_Q),     .A1(T5681_Y), .A0(T1484_Y));
KC_AOI22_X1 T5668 ( .Y(T5668_Y), .B1(T5669_Y), .B0(T13691_Q),     .A1(T5680_Y), .A0(T2565_Y));
KC_AOI22_X1 T5667 ( .Y(T5667_Y), .B1(T10807_Y), .B0(T14662_Q),     .A1(T5701_Y), .A0(T1484_Y));
KC_AOI22_X1 T5666 ( .Y(T5666_Y), .B1(T10373_Y), .B0(T1484_Y),     .A1(T5671_Y), .A0(T13716_Q));
KC_AOI22_X1 T5665 ( .Y(T5665_Y), .B1(T10362_Y), .B0(T13693_Q),     .A1(T10360_Y), .A0(T13736_Q));
KC_AOI22_X1 T10783 ( .Y(T10783_Y), .B1(T9706_Y), .B0(T14636_Q),     .A1(T1545_Y), .A0(T14634_Q));
KC_AOI22_X1 T10771 ( .Y(T10771_Y), .B1(T14636_Q), .B0(T10359_Y),     .A1(T14634_Q), .A0(T4889_Y));
KC_AOI22_X1 T7538 ( .Y(T7538_Y), .B1(T9706_Y), .B0(T13789_Q),     .A1(T1545_Y), .A0(T13854_Q));
KC_AOI22_X1 T7537 ( .Y(T7537_Y), .B1(T13855_Q), .B0(T10359_Y),     .A1(T13811_Q), .A0(T4889_Y));
KC_AOI22_X1 T7536 ( .Y(T7536_Y), .B1(T9706_Y), .B0(T13855_Q),     .A1(T1545_Y), .A0(T13811_Q));
KC_AOI22_X1 T7535 ( .Y(T7535_Y), .B1(T10359_Y), .B0(T13810_Q),     .A1(T13813_Q), .A0(T4889_Y));
KC_AOI22_X1 T7531 ( .Y(T7531_Y), .B1(T9706_Y), .B0(T13790_Q),     .A1(T1545_Y), .A0(T13788_Q));
KC_AOI22_X1 T7529 ( .Y(T7529_Y), .B1(T13789_Q), .B0(T10359_Y),     .A1(T13854_Q), .A0(T4889_Y));
KC_AOI22_X1 T7508 ( .Y(T7508_Y), .B1(T7509_Y), .B0(T13812_Q),     .A1(T5696_Y), .A0(T1484_Y));
KC_AOI22_X1 T7488 ( .Y(T7488_Y), .B1(T7540_Y), .B0(T13978_Q),     .A1(T5695_Y), .A0(T1484_Y));
KC_AOI22_X1 T7487 ( .Y(T7487_Y), .B1(T9706_Y), .B0(T13810_Q),     .A1(T1545_Y), .A0(T13813_Q));
KC_AOI22_X1 T7790 ( .Y(T7790_Y), .B1(T7776_Y), .B0(T1484_Y),     .A1(T7788_Y), .A0(T13960_Q));
KC_AOI22_X1 T7785 ( .Y(T7785_Y), .B1(T7786_Y), .B0(T14013_Q),     .A1(T7717_Y), .A0(T1484_Y));
KC_AOI22_X1 T7784 ( .Y(T7784_Y), .B1(T7789_Y), .B0(T13943_Q),     .A1(T7739_Y), .A0(T1484_Y));
KC_AOI22_X1 T7783 ( .Y(T7783_Y), .B1(T7701_Y), .B0(T13958_Q),     .A1(T9790_Y), .A0(T1484_Y));
KC_AOI22_X1 T7756 ( .Y(T7756_Y), .B1(T13980_Q), .B0(T10359_Y),     .A1(T13979_Q), .A0(T4889_Y));
KC_AOI22_X1 T7755 ( .Y(T7755_Y), .B1(T9706_Y), .B0(T13981_Q),     .A1(T1545_Y), .A0(T13995_Q));
KC_AOI22_X1 T7743 ( .Y(T7743_Y), .B1(T13981_Q), .B0(T10359_Y),     .A1(T13995_Q), .A0(T4889_Y));
KC_AOI22_X1 T7720 ( .Y(T7720_Y), .B1(T9706_Y), .B0(T13980_Q),     .A1(T1545_Y), .A0(T13979_Q));
KC_AOI22_X1 T7706 ( .Y(T7706_Y), .B1(T7787_Y), .B0(T13959_Q),     .A1(T7548_Y), .A0(T1484_Y));
KC_AOI22_X1 T7699 ( .Y(T7699_Y), .B1(T7700_Y), .B0(T13942_Q),     .A1(T10338_Y), .A0(T1484_Y));
KC_AOI22_X1 T10761 ( .Y(T10761_Y), .B1(T10760_Y), .B0(T14610_Q),     .A1(T1484_Y), .A0(T7990_Y));
KC_AOI22_X1 T10752 ( .Y(T10752_Y), .B1(T10306_Y), .B0(T14274_Q),     .A1(T10009_Y), .A0(T14119_Q));
KC_AOI22_X1 T10750 ( .Y(T10750_Y), .B1(T14601_Q), .B0(T9893_Y),     .A1(T14117_Q), .A0(T15229_Y));
KC_AOI22_X1 T10749 ( .Y(T10749_Y), .B1(T14602_Q), .B0(T9893_Y),     .A1(T14116_Q), .A0(T15229_Y));
KC_AOI22_X1 T10748 ( .Y(T10748_Y), .B1(T10033_Y), .B0(T14602_Q),     .A1(T15228_Y), .A0(T14116_Q));
KC_AOI22_X1 T10747 ( .Y(T10747_Y), .B1(T12094_Y), .B0(T14277_Q),     .A1(T8000_Y), .A0(T14273_Q));
KC_AOI22_X1 T8014 ( .Y(T8014_Y), .B1(T7970_Y), .B0(T14616_Q),     .A1(T7945_Y), .A0(T1484_Y));
KC_AOI22_X1 T8012 ( .Y(T8012_Y), .B1(T7963_Y), .B0(T14129_Q),     .A1(T7928_Y), .A0(T2565_Y));
KC_AOI22_X1 T7987 ( .Y(T7987_Y), .B1(T14604_Q), .B0(T1584_Y),     .A1(T14115_Q), .A0(T1585_Y));
KC_AOI22_X1 T7967 ( .Y(T7967_Y), .B1(T7971_Y), .B0(T14614_Q),     .A1(T9999_Y), .A0(T1484_Y));
KC_AOI22_X1 T7959 ( .Y(T7959_Y), .B1(T7962_Y), .B0(T14126_Q),     .A1(T10012_Y), .A0(T2565_Y));
KC_AOI22_X1 T7958 ( .Y(T7958_Y), .B1(T7960_Y), .B0(T14128_Q),     .A1(T7934_Y), .A0(T2565_Y));
KC_AOI22_X1 T7957 ( .Y(T7957_Y), .B1(T7961_Y), .B0(T14127_Q),     .A1(T9997_Y), .A0(T1484_Y));
KC_AOI22_X1 T7940 ( .Y(T7940_Y), .B1(T10033_Y), .B0(T14107_Q),     .A1(T15228_Y), .A0(T14254_Q));
KC_AOI22_X1 T7933 ( .Y(T7933_Y), .B1(T8862_Y), .B0(T14103_Q),     .A1(T9883_Y), .A0(T14104_Q));
KC_AOI22_X1 T7932 ( .Y(T7932_Y), .B1(T8862_Y), .B0(T14102_Q),     .A1(T9883_Y), .A0(T14105_Q));
KC_AOI22_X1 T7931 ( .Y(T7931_Y), .B1(T14103_Q), .B0(T1584_Y),     .A1(T14104_Q), .A0(T1585_Y));
KC_AOI22_X1 T7930 ( .Y(T7930_Y), .B1(T14102_Q), .B0(T1584_Y),     .A1(T14105_Q), .A0(T1585_Y));
KC_AOI22_X1 T7929 ( .Y(T7929_Y), .B1(T8862_Y), .B0(T14604_Q),     .A1(T9883_Y), .A0(T14115_Q));
KC_AOI22_X1 T1480 ( .Y(T1480_Y), .B1(T14274_Q), .B0(T9892_Y),     .A1(T14119_Q), .A0(T9902_Y));
KC_AOI22_X1 T10715 ( .Y(T10715_Y), .B1(T10306_Y), .B0(T14272_Q),     .A1(T10009_Y), .A0(T14275_Q));
KC_AOI22_X1 T10714 ( .Y(T10714_Y), .B1(T14272_Q), .B0(T9892_Y),     .A1(T14275_Q), .A0(T9902_Y));
KC_AOI22_X1 T10713 ( .Y(T10713_Y), .B1(T10033_Y), .B0(T14601_Q),     .A1(T15228_Y), .A0(T14117_Q));
KC_AOI22_X1 T10712 ( .Y(T10712_Y), .B1(T14277_Q), .B0(T12088_Y),     .A1(T14273_Q), .A0(T8011_Y));
KC_AOI22_X1 T10731 ( .Y(T10731_Y), .B1(T12094_Y), .B0(T14379_Q),     .A1(T8000_Y), .A0(T14373_Q));
KC_AOI22_X1 T10730 ( .Y(T10730_Y), .B1(T14379_Q), .B0(T12088_Y),     .A1(T14373_Q), .A0(T8011_Y));
KC_AOI22_X1 T1511 ( .Y(T1511_Y), .B1(T12094_Y), .B0(T14596_Q),     .A1(T8000_Y), .A0(T14595_Q));
KC_AOI22_X1 T1512 ( .Y(T1512_Y), .B1(T14596_Q), .B0(T12088_Y),     .A1(T14595_Q), .A0(T8011_Y));
KC_AOI22_X1 T1513 ( .Y(T1513_Y), .B1(T12094_Y), .B0(T14456_Q),     .A1(T8000_Y), .A0(T14455_Q));
KC_AOI22_X1 T10836 ( .Y(T10836_Y), .B1(T12325_Y), .B0(T13493_Q),     .A1(T12324_Y), .A0(T16505_Y));
KC_AOI22_X1 T10835 ( .Y(T10835_Y), .B1(T9580_Y), .B0(T13374_Q),     .A1(T2027_Y), .A0(T13341_Q));
KC_AOI22_X1 T6869 ( .Y(T6869_Y), .B1(T13374_Q), .B0(T12075_Y),     .A1(T13341_Q), .A0(T7323_Y));
KC_AOI22_X1 T6865 ( .Y(T6865_Y), .B1(T9580_Y), .B0(T13373_Q),     .A1(T2027_Y), .A0(T13370_Q));
KC_AOI22_X1 T6864 ( .Y(T6864_Y), .B1(T13343_Q), .B0(T12075_Y),     .A1(T13375_Q), .A0(T7323_Y));
KC_AOI22_X1 T6863 ( .Y(T6863_Y), .B1(T9580_Y), .B0(T13343_Q),     .A1(T2027_Y), .A0(T13375_Q));
KC_AOI22_X1 T10848 ( .Y(T10848_Y), .B1(T9580_Y), .B0(T14705_Q),     .A1(T2027_Y), .A0(T14704_Q));
KC_AOI22_X1 T6988 ( .Y(T6988_Y), .B1(T6452_Y), .B0(T13473_Q),     .A1(T1632_Y), .A0(T13463_Q));
KC_AOI22_X1 T6974 ( .Y(T6974_Y), .B1(T6452_Y), .B0(T13465_Q),     .A1(T1632_Y), .A0(T13494_Q));
KC_AOI22_X1 T10871 ( .Y(T10871_Y), .B1(T12075_Y), .B0(T14724_Q),     .A1(T13574_Q), .A0(T7323_Y));
KC_AOI22_X1 T10870 ( .Y(T10870_Y), .B1(T14721_Q), .B0(T12075_Y),     .A1(T14723_Q), .A0(T7323_Y));
KC_AOI22_X1 T7208 ( .Y(T7208_Y), .B1(T13604_Q), .B0(T12075_Y),     .A1(T13605_Q), .A0(T7323_Y));
KC_AOI22_X1 T7188 ( .Y(T7188_Y), .B1(T7177_Y), .B0(T13657_Q),     .A1(T6984_Y), .A0(T4937_Y));
KC_AOI22_X1 T7187 ( .Y(T7187_Y), .B1(T7191_Y), .B0(T13603_Q),     .A1(T7017_Y), .A0(T9642_Y));
KC_AOI22_X1 T7175 ( .Y(T7175_Y), .B1(T9580_Y), .B0(T14724_Q),     .A1(T3640_Y), .A0(T13574_Q));
KC_AOI22_X1 T7170 ( .Y(T7170_Y), .B1(T9580_Y), .B0(T13596_Q),     .A1(T3640_Y), .A0(T13582_Q));
KC_AOI22_X1 T7169 ( .Y(T7169_Y), .B1(T13596_Q), .B0(T12075_Y),     .A1(T13582_Q), .A0(T7323_Y));
KC_AOI22_X1 T7348 ( .Y(T7348_Y), .B1(T7349_Y), .B0(T14720_Q),     .A1(T4937_Y), .A0(T5661_Y));
KC_AOI22_X1 T5660 ( .Y(T5660_Y), .B1(T13714_Q), .B0(T10361_Y),     .A1(T13734_Q), .A0(T15247_Y));
KC_AOI22_X1 T5659 ( .Y(T5659_Y), .B1(T10346_Y), .B0(T13714_Q),     .A1(T15245_Y), .A0(T13734_Q));
KC_AOI22_X1 T5658 ( .Y(T5658_Y), .B1(T10346_Y), .B0(T13688_Q),     .A1(T15245_Y), .A0(T13690_Q));
KC_AOI22_X1 T5657 ( .Y(T5657_Y), .B1(T9707_Y), .B0(T13718_Q),     .A1(T10347_Y), .A0(T13712_Q));
KC_AOI22_X1 T5654 ( .Y(T5654_Y), .B1(T13715_Q), .B0(T10361_Y),     .A1(T13733_Q), .A0(T15247_Y));
KC_AOI22_X1 T5653 ( .Y(T5653_Y), .B1(T10361_Y), .B0(T13688_Q),     .A1(T15247_Y), .A0(T13690_Q));
KC_AOI22_X1 T5652 ( .Y(T5652_Y), .B1(T13718_Q), .B0(T10362_Y),     .A1(T13712_Q), .A0(T10360_Y));
KC_AOI22_X1 T10806 ( .Y(T10806_Y), .B1(T13713_Q), .B0(T10362_Y),     .A1(T14740_Q), .A0(T10360_Y));
KC_AOI22_X1 T10805 ( .Y(T10805_Y), .B1(T9707_Y), .B0(T13713_Q),     .A1(T10347_Y), .A0(T14740_Q));
KC_AOI22_X1 T10800 ( .Y(T10800_Y), .B1(T14655_Q), .B0(T10362_Y),     .A1(T14742_Q), .A0(T10360_Y));
KC_AOI22_X1 T10798 ( .Y(T10798_Y), .B1(T9707_Y), .B0(T14655_Q),     .A1(T10347_Y), .A0(T14742_Q));
KC_AOI22_X1 T10775 ( .Y(T10775_Y), .B1(T13996_Q), .B0(T10358_Y),     .A1(T13976_Q), .A0(T9712_Y));
KC_AOI22_X1 T10774 ( .Y(T10774_Y), .B1(T13975_Q), .B0(T10361_Y),     .A1(T15049_Q), .A0(T15247_Y));
KC_AOI22_X1 T10773 ( .Y(T10773_Y), .B1(T9784_Q), .B0(T10362_Y),     .A1(T13977_Q), .A0(T10360_Y));
KC_AOI22_X1 T10772 ( .Y(T10772_Y), .B1(T13785_Q), .B0(T10358_Y),     .A1(T13851_Q), .A0(T9712_Y));
KC_AOI22_X1 T10765 ( .Y(T10765_Y), .B1(T13974_Q), .B0(T10361_Y),     .A1(T13993_Q), .A0(T15247_Y));
KC_AOI22_X1 T7532 ( .Y(T7532_Y), .B1(T13790_Q), .B0(T10359_Y),     .A1(T13788_Q), .A0(T4889_Y));
KC_AOI22_X1 T7530 ( .Y(T7530_Y), .B1(T10346_Y), .B0(T13803_Q),     .A1(T15245_Y), .A0(T13850_Q));
KC_AOI22_X1 T7527 ( .Y(T7527_Y), .B1(T13803_Q), .B0(T10361_Y),     .A1(T13850_Q), .A0(T15247_Y));
KC_AOI22_X1 T7524 ( .Y(T7524_Y), .B1(T13786_Q), .B0(T10359_Y),     .A1(T13852_Q), .A0(T4889_Y));
KC_AOI22_X1 T7521 ( .Y(T7521_Y), .B1(T9706_Y), .B0(T13786_Q),     .A1(T1545_Y), .A0(T13852_Q));
KC_AOI22_X1 T7506 ( .Y(T7506_Y), .B1(T14657_Q), .B0(T10358_Y),     .A1(T14658_Q), .A0(T9712_Y));
KC_AOI22_X1 T7505 ( .Y(T7505_Y), .B1(T9704_Y), .B0(T14657_Q),     .A1(T9705_Y), .A0(T14658_Q));
KC_AOI22_X1 T7501 ( .Y(T7501_Y), .B1(T9704_Y), .B0(T13809_Q),     .A1(T9705_Y), .A0(T13833_Q));
KC_AOI22_X1 T7500 ( .Y(T7500_Y), .B1(T13809_Q), .B0(T10358_Y),     .A1(T13833_Q), .A0(T9712_Y));
KC_AOI22_X1 T7486 ( .Y(T7486_Y), .B1(T9707_Y), .B0(T13808_Q),     .A1(T10347_Y), .A0(T13787_Q));
KC_AOI22_X1 T7485 ( .Y(T7485_Y), .B1(T13807_Q), .B0(T10358_Y),     .A1(T13853_Q), .A0(T9712_Y));
KC_AOI22_X1 T7484 ( .Y(T7484_Y), .B1(T13808_Q), .B0(T10362_Y),     .A1(T13787_Q), .A0(T10360_Y));
KC_AOI22_X1 T7483 ( .Y(T7483_Y), .B1(T9704_Y), .B0(T13807_Q),     .A1(T9705_Y), .A0(T13853_Q));
KC_AOI22_X1 T7476 ( .Y(T7476_Y), .B1(T13846_Q), .B0(T10358_Y),     .A1(T13798_Q), .A0(T9712_Y));
KC_AOI22_X1 T7752 ( .Y(T7752_Y), .B1(T10346_Y), .B0(T13974_Q),     .A1(T15245_Y), .A0(T13993_Q));
KC_AOI22_X1 T7751 ( .Y(T7751_Y), .B1(T7732_Y), .B0(T12086_Y),     .A1(T7463_Y), .A0(T2531_Y));
KC_AOI22_X1 T7750 ( .Y(T7750_Y), .B1(T7733_Y), .B0(T12086_Y),     .A1(T7507_Y), .A0(T2531_Y));
KC_AOI22_X1 T7749 ( .Y(T7749_Y), .B1(T9704_Y), .B0(T14633_Q),     .A1(T9705_Y), .A0(T14632_Q));
KC_AOI22_X1 T7748 ( .Y(T7748_Y), .B1(T7467_Y), .B0(T12086_Y),     .A1(T10365_Y), .A0(T2531_Y));
KC_AOI22_X1 T7747 ( .Y(T7747_Y), .B1(T10346_Y), .B0(T14011_Q),     .A1(T15245_Y), .A0(T13955_Q));
KC_AOI22_X1 T7746 ( .Y(T7746_Y), .B1(T9707_Y), .B0(T13992_Q),     .A1(T10347_Y), .A0(T13991_Q));
KC_AOI22_X1 T7745 ( .Y(T7745_Y), .B1(T9707_Y), .B0(T13954_Q),     .A1(T10347_Y), .A0(T16178_Q));
KC_AOI22_X1 T7744 ( .Y(T7744_Y), .B1(T9707_Y), .B0(T9784_Q),     .A1(T10347_Y), .A0(T13977_Q));
KC_AOI22_X1 T7742 ( .Y(T7742_Y), .B1(T10346_Y), .B0(T13975_Q),     .A1(T15245_Y), .A0(T15049_Q));
KC_AOI22_X1 T10746 ( .Y(T10746_Y), .B1(T14599_Q), .B0(T9893_Y),     .A1(T14099_Q), .A0(T15229_Y));
KC_AOI22_X1 T10745 ( .Y(T10745_Y), .B1(T8862_Y), .B0(T14101_Q),     .A1(T9883_Y), .A0(T14114_Q));
KC_AOI22_X1 T10744 ( .Y(T10744_Y), .B1(T14600_Q), .B0(T9893_Y),     .A1(T14267_Q), .A0(T15229_Y));
KC_AOI22_X1 T8009 ( .Y(T8009_Y), .B1(T7954_Y), .B0(T14611_Q),     .A1(T7935_Y), .A0(T2565_Y));
KC_AOI22_X1 T8008 ( .Y(T8008_Y), .B1(T7955_Y), .B0(T14125_Q),     .A1(T10310_Y), .A0(T2565_Y));
KC_AOI22_X1 T8007 ( .Y(T8007_Y), .B1(T7956_Y), .B0(T14124_Q),     .A1(T9994_Y), .A0(T2565_Y));
KC_AOI22_X1 T8006 ( .Y(T8006_Y), .B1(T8010_Y), .B0(T14609_Q),     .A1(T10010_Y), .A0(T2565_Y));
KC_AOI22_X1 T7926 ( .Y(T7926_Y), .B1(T14100_Q), .B0(T1584_Y),     .A1(T14098_Q), .A0(T1585_Y));
KC_AOI22_X1 T10711 ( .Y(T10711_Y), .B1(T8862_Y), .B0(T14247_Q),     .A1(T9883_Y), .A0(T14268_Q));
KC_AOI22_X1 T10710 ( .Y(T10710_Y), .B1(T8862_Y), .B0(T14100_Q),     .A1(T9883_Y), .A0(T14098_Q));
KC_AOI22_X1 T10709 ( .Y(T10709_Y), .B1(T10033_Y), .B0(T14599_Q),     .A1(T15228_Y), .A0(T14099_Q));
KC_AOI22_X1 T10708 ( .Y(T10708_Y), .B1(T10306_Y), .B0(T14246_Q),     .A1(T10009_Y), .A0(T14266_Q));
KC_AOI22_X1 T10707 ( .Y(T10707_Y), .B1(T14246_Q), .B0(T9892_Y),     .A1(T14266_Q), .A0(T9902_Y));
KC_AOI22_X1 T10706 ( .Y(T10706_Y), .B1(T10306_Y), .B0(T14265_Q),     .A1(T10009_Y), .A0(T14249_Q));
KC_AOI22_X1 T10704 ( .Y(T10704_Y), .B1(T14243_Q), .B0(T9892_Y),     .A1(T14264_Q), .A0(T9902_Y));
KC_AOI22_X1 T10703 ( .Y(T10703_Y), .B1(T10306_Y), .B0(T14243_Q),     .A1(T10009_Y), .A0(T14264_Q));
KC_AOI22_X1 T10699 ( .Y(T10699_Y), .B1(T10033_Y), .B0(T14600_Q),     .A1(T15228_Y), .A0(T14267_Q));
KC_AOI22_X1 T10688 ( .Y(T10688_Y), .B1(T10306_Y), .B0(T14226_Q),     .A1(T10009_Y), .A0(T14235_Q));
KC_AOI22_X1 T10687 ( .Y(T10687_Y), .B1(T14269_Q), .B0(T9893_Y),     .A1(T14248_Q), .A0(T15229_Y));
KC_AOI22_X1 T10686 ( .Y(T10686_Y), .B1(T14247_Q), .B0(T1584_Y),     .A1(T14268_Q), .A0(T1585_Y));
KC_AOI22_X1 T10685 ( .Y(T10685_Y), .B1(T14226_Q), .B0(T9892_Y),     .A1(T14235_Q), .A0(T9902_Y));
KC_AOI22_X1 T10684 ( .Y(T10684_Y), .B1(T14232_Q), .B0(T9892_Y),     .A1(T14242_Q), .A0(T9902_Y));
KC_AOI22_X1 T10683 ( .Y(T10683_Y), .B1(T10033_Y), .B0(T14269_Q),     .A1(T15228_Y), .A0(T14248_Q));
KC_AOI22_X1 T10680 ( .Y(T10680_Y), .B1(T14234_Q), .B0(T9893_Y),     .A1(T14245_Q), .A0(T15229_Y));
KC_AOI22_X1 T10679 ( .Y(T10679_Y), .B1(T14223_Q), .B0(T9893_Y),     .A1(T14244_Q), .A0(T15229_Y));
KC_AOI22_X1 T10678 ( .Y(T10678_Y), .B1(T14222_Q), .B0(T9893_Y),     .A1(T14233_Q), .A0(T15229_Y));
KC_AOI22_X1 T10677 ( .Y(T10677_Y), .B1(T10306_Y), .B0(T14232_Q),     .A1(T10009_Y), .A0(T14242_Q));
KC_AOI22_X1 T10676 ( .Y(T10676_Y), .B1(T10033_Y), .B0(T14222_Q),     .A1(T15228_Y), .A0(T14233_Q));
KC_AOI22_X1 T10670 ( .Y(T10670_Y), .B1(T14220_Q), .B0(T1584_Y),     .A1(T14206_Q), .A0(T1585_Y));
KC_AOI22_X1 T10669 ( .Y(T10669_Y), .B1(T10033_Y), .B0(T14234_Q),     .A1(T15228_Y), .A0(T14245_Q));
KC_AOI22_X1 T10668 ( .Y(T10668_Y), .B1(T8862_Y), .B0(T14220_Q),     .A1(T9883_Y), .A0(T14206_Q));
KC_AOI22_X1 T10666 ( .Y(T10666_Y), .B1(T8862_Y), .B0(T14219_Q),     .A1(T9883_Y), .A0(T14208_Q));
KC_AOI22_X1 T10665 ( .Y(T10665_Y), .B1(T10033_Y), .B0(T14223_Q),     .A1(T15228_Y), .A0(T14244_Q));
KC_AOI22_X1 T10663 ( .Y(T10663_Y), .B1(T10306_Y), .B0(T14204_Q),     .A1(T10009_Y), .A0(T14205_Q));
KC_AOI22_X1 T10662 ( .Y(T10662_Y), .B1(T14204_Q), .B0(T9892_Y),     .A1(T14205_Q), .A0(T9902_Y));
KC_AOI22_X1 T10655 ( .Y(T10655_Y), .B1(T8862_Y), .B0(T14221_Q),     .A1(T9883_Y), .A0(T14207_Q));
KC_AOI22_X1 T10654 ( .Y(T10654_Y), .B1(T14221_Q), .B0(T1584_Y),     .A1(T14207_Q), .A0(T1585_Y));
KC_AOI22_X1 T10653 ( .Y(T10653_Y), .B1(T14217_Q), .B0(T9892_Y),     .A1(T14218_Q), .A0(T9902_Y));
KC_AOI22_X1 T10733 ( .Y(T10733_Y), .B1(T14376_Q), .B0(T12088_Y),     .A1(T14383_Q), .A0(T8011_Y));
KC_AOI22_X1 T10729 ( .Y(T10729_Y), .B1(T12094_Y), .B0(T13328_Q),     .A1(T8000_Y), .A0(T14453_Q));
KC_AOI22_X1 T10726 ( .Y(T10726_Y), .B1(T14371_Q), .B0(T12088_Y),     .A1(T14590_Q), .A0(T8011_Y));
KC_AOI22_X1 T1605 ( .Y(T1605_Y), .B1(T13328_Q), .B0(T12088_Y),     .A1(T14453_Q), .A0(T8011_Y));
KC_AOI22_X1 T1606 ( .Y(T1606_Y), .B1(T14593_Q), .B0(T12088_Y),     .A1(T14454_Q), .A0(T8011_Y));
KC_AOI22_X1 T1607 ( .Y(T1607_Y), .B1(T14458_Q), .B0(T12088_Y),     .A1(T14457_Q), .A0(T8011_Y));
KC_AOI22_X1 T6893 ( .Y(T6893_Y), .B1(T13373_Q), .B0(T12075_Y),     .A1(T13370_Q), .A0(T7323_Y));
KC_AOI22_X1 T6892 ( .Y(T6892_Y), .B1(T13372_Q), .B0(T12075_Y),     .A1(T13359_Q), .A0(T7323_Y));
KC_AOI22_X1 T6868 ( .Y(T6868_Y), .B1(T9580_Y), .B0(T13358_Q),     .A1(T2027_Y), .A0(T13360_Q));
KC_AOI22_X1 T6867 ( .Y(T6867_Y), .B1(T9580_Y), .B0(T13372_Q),     .A1(T2027_Y), .A0(T13359_Q));
KC_AOI22_X1 T6866 ( .Y(T6866_Y), .B1(T13358_Q), .B0(T12075_Y),     .A1(T13360_Q), .A0(T7323_Y));
KC_AOI22_X1 T1618 ( .Y(T1618_Y), .B1(T9580_Y), .B0(T15045_Q),     .A1(T2027_Y), .A0(T13416_Q));
KC_AOI22_X1 T7006 ( .Y(T7006_Y), .B1(T14686_Q), .B0(T12076_Y),     .A1(T14685_Q), .A0(T12074_Y));
KC_AOI22_X1 T7005 ( .Y(T7005_Y), .B1(T13480_Q), .B0(T12077_Y),     .A1(T13479_Q), .A0(T12078_Y));
KC_AOI22_X1 T7004 ( .Y(T7004_Y), .B1(T6452_Y), .B0(T13480_Q),     .A1(T1632_Y), .A0(T13479_Q));
KC_AOI22_X1 T6987 ( .Y(T6987_Y), .B1(T13477_Q), .B0(T12077_Y),     .A1(T13488_Q), .A0(T12078_Y));
KC_AOI22_X1 T6986 ( .Y(T6986_Y), .B1(T13474_Q), .B0(T1547_Y),     .A1(T13476_Q), .A0(T15202_Y));
KC_AOI22_X1 T6985 ( .Y(T6985_Y), .B1(T13473_Q), .B0(T12077_Y),     .A1(T13463_Q), .A0(T12078_Y));
KC_AOI22_X1 T6979 ( .Y(T6979_Y), .B1(T13442_Q), .B0(T1547_Y),     .A1(T13444_Q), .A0(T15202_Y));
KC_AOI22_X1 T6978 ( .Y(T6978_Y), .B1(T6452_Y), .B0(T13477_Q),     .A1(T1632_Y), .A0(T13488_Q));
KC_AOI22_X1 T6977 ( .Y(T6977_Y), .B1(T10397_Y), .B0(T13474_Q),     .A1(T15204_Y), .A0(T13476_Q));
KC_AOI22_X1 T6976 ( .Y(T6976_Y), .B1(T12325_Y), .B0(T13447_Q),     .A1(T12324_Y), .A0(T13487_Q));
KC_AOI22_X1 T6973 ( .Y(T6973_Y), .B1(T10397_Y), .B0(T13442_Q),     .A1(T15204_Y), .A0(T13444_Q));
KC_AOI22_X1 T6972 ( .Y(T6972_Y), .B1(T13447_Q), .B0(T12076_Y),     .A1(T13487_Q), .A0(T12074_Y));
KC_AOI22_X1 T5720 ( .Y(T5720_Y), .B1(T13443_Q), .B0(T1547_Y),     .A1(T13475_Q), .A0(T15202_Y));
KC_AOI22_X1 T5719 ( .Y(T5719_Y), .B1(T10397_Y), .B0(T13563_Q),     .A1(T15204_Y), .A0(T13536_Q));
KC_AOI22_X1 T5718 ( .Y(T5718_Y), .B1(T14809_Q), .B0(T12076_Y),     .A1(T13489_Q), .A0(T12074_Y));
KC_AOI22_X1 T1619 ( .Y(T1619_Y), .B1(T10397_Y), .B0(T13599_Q),     .A1(T15204_Y), .A0(T13601_Q));
KC_AOI22_X1 T1623 ( .Y(T1623_Y), .B1(T12325_Y), .B0(T14809_Q),     .A1(T12324_Y), .A0(T13489_Q));
KC_AOI22_X1 T1624 ( .Y(T1624_Y), .B1(T10397_Y), .B0(T13443_Q),     .A1(T15204_Y), .A0(T13475_Q));
KC_AOI22_X1 T10873 ( .Y(T10873_Y), .B1(T10397_Y), .B0(T13662_Q),     .A1(T15204_Y), .A0(T14774_Q));
KC_AOI22_X1 T10872 ( .Y(T10872_Y), .B1(T1547_Y), .B0(T13662_Q),     .A1(T15202_Y), .A0(T14774_Q));
KC_AOI22_X1 T7210 ( .Y(T7210_Y), .B1(T6452_Y), .B0(T13598_Q),     .A1(T1632_Y), .A0(T13602_Q));
KC_AOI22_X1 T7209 ( .Y(T7209_Y), .B1(T13598_Q), .B0(T12077_Y),     .A1(T13602_Q), .A0(T12078_Y));
KC_AOI22_X1 T7174 ( .Y(T7174_Y), .B1(T14718_Q), .B0(T12077_Y),     .A1(T14719_Q), .A0(T12078_Y));
KC_AOI22_X1 T7173 ( .Y(T7173_Y), .B1(T12077_Y), .B0(T13579_Q),     .A1(T12078_Y), .A0(T13595_Q));
KC_AOI22_X1 T7172 ( .Y(T7172_Y), .B1(T6452_Y), .B0(T13579_Q),     .A1(T1632_Y), .A0(T13595_Q));
KC_AOI22_X1 T7171 ( .Y(T7171_Y), .B1(T6452_Y), .B0(T14718_Q),     .A1(T1632_Y), .A0(T14719_Q));
KC_AOI22_X1 T7125 ( .Y(T7125_Y), .B1(T13572_Q), .B0(T1547_Y),     .A1(T13570_Q), .A0(T15202_Y));
KC_AOI22_X1 T7124 ( .Y(T7124_Y), .B1(T13571_Q), .B0(T12076_Y),     .A1(T13600_Q), .A0(T12074_Y));
KC_AOI22_X1 T7123 ( .Y(T7123_Y), .B1(T12325_Y), .B0(T13571_Q),     .A1(T12324_Y), .A0(T13600_Q));
KC_AOI22_X1 T1625 ( .Y(T1625_Y), .B1(T10397_Y), .B0(T13572_Q),     .A1(T15204_Y), .A0(T13570_Q));
KC_AOI22_X1 T1626 ( .Y(T1626_Y), .B1(T12325_Y), .B0(T14789_Q),     .A1(T12324_Y), .A0(T13683_Q));
KC_AOI22_X1 T1629 ( .Y(T1629_Y), .B1(T13632_Q), .B0(T1547_Y),     .A1(T13684_Q), .A0(T15202_Y));
KC_AOI22_X1 T1630 ( .Y(T1630_Y), .B1(T10397_Y), .B0(T13632_Q),     .A1(T15204_Y), .A0(T13684_Q));
KC_AOI22_X1 T7345 ( .Y(T7345_Y), .B1(T12325_Y), .B0(T13685_Q),     .A1(T12324_Y), .A0(T13687_Q));
KC_AOI22_X1 T7344 ( .Y(T7344_Y), .B1(T13685_Q), .B0(T12076_Y),     .A1(T13687_Q), .A0(T12074_Y));
KC_AOI22_X1 T7319 ( .Y(T7319_Y), .B1(T6461_Q), .B0(T1547_Y),     .A1(T13581_Q), .A0(T15202_Y));
KC_AOI22_X1 T10799 ( .Y(T10799_Y), .B1(T13832_Q), .B0(T10362_Y),     .A1(T14654_Q), .A0(T10360_Y));
KC_AOI22_X1 T10764 ( .Y(T10764_Y), .B1(T13989_Q), .B0(T10359_Y),     .A1(T14626_Q), .A0(T4889_Y));
KC_AOI22_X1 T10763 ( .Y(T10763_Y), .B1(T13972_Q), .B0(T10359_Y),     .A1(T13988_Q), .A0(T4889_Y));
KC_AOI22_X1 T10650 ( .Y(T10650_Y), .B1(T9707_Y), .B0(T13832_Q),     .A1(T10347_Y), .A0(T14654_Q));
KC_AOI22_X1 T7526 ( .Y(T7526_Y), .B1(T9704_Y), .B0(T13987_Q),     .A1(T9705_Y), .A0(T13984_Q));
KC_AOI22_X1 T7525 ( .Y(T7525_Y), .B1(T13844_Q), .B0(T10358_Y),     .A1(T13847_Q), .A0(T9712_Y));
KC_AOI22_X1 T7523 ( .Y(T7523_Y), .B1(T9707_Y), .B0(T13848_Q),     .A1(T10347_Y), .A0(T13845_Q));
KC_AOI22_X1 T7522 ( .Y(T7522_Y), .B1(T9704_Y), .B0(T13844_Q),     .A1(T9705_Y), .A0(T13847_Q));
KC_AOI22_X1 T7503 ( .Y(T7503_Y), .B1(T14653_Q), .B0(T10362_Y),     .A1(T14656_Q), .A0(T10360_Y));
KC_AOI22_X1 T7502 ( .Y(T7502_Y), .B1(T9707_Y), .B0(T14653_Q),     .A1(T10347_Y), .A0(T14656_Q));
KC_AOI22_X1 T7480 ( .Y(T7480_Y), .B1(T9704_Y), .B0(T13846_Q),     .A1(T9705_Y), .A0(T13798_Q));
KC_AOI22_X1 T7479 ( .Y(T7479_Y), .B1(T13800_Q), .B0(T10362_Y),     .A1(T13802_Q), .A0(T10360_Y));
KC_AOI22_X1 T7478 ( .Y(T7478_Y), .B1(T9704_Y), .B0(T13799_Q),     .A1(T9705_Y), .A0(T13801_Q));
KC_AOI22_X1 T7477 ( .Y(T7477_Y), .B1(T13799_Q), .B0(T10358_Y),     .A1(T13801_Q), .A0(T9712_Y));
KC_AOI22_X1 T7475 ( .Y(T7475_Y), .B1(T9707_Y), .B0(T13800_Q),     .A1(T10347_Y), .A0(T13802_Q));
KC_AOI22_X1 T7474 ( .Y(T7474_Y), .B1(T10346_Y), .B0(T14841_Q),     .A1(T15245_Y), .A0(T13923_Q));
KC_AOI22_X1 T7462 ( .Y(T7462_Y), .B1(T9706_Y), .B0(T14630_Q),     .A1(T1545_Y), .A0(T14631_Q));
KC_AOI22_X1 T7461 ( .Y(T7461_Y), .B1(T13987_Q), .B0(T10358_Y),     .A1(T13984_Q), .A0(T9712_Y));
KC_AOI22_X1 T7460 ( .Y(T7460_Y), .B1(T9706_Y), .B0(T13989_Q),     .A1(T1545_Y), .A0(T14626_Q));
KC_AOI22_X1 T1639 ( .Y(T1639_Y), .B1(T9706_Y), .B0(T13985_Q),     .A1(T1545_Y), .A0(T13990_Q));
KC_AOI22_X1 T1641 ( .Y(T1641_Y), .B1(T13848_Q), .B0(T10362_Y),     .A1(T13845_Q), .A0(T10360_Y));
KC_AOI22_X1 T1642 ( .Y(T1642_Y), .B1(T10346_Y), .B0(T13922_Q),     .A1(T15245_Y), .A0(T13921_Q));
KC_AOI22_X1 T1643 ( .Y(T1643_Y), .B1(T13922_Q), .B0(T10361_Y),     .A1(T13921_Q), .A0(T15247_Y));
KC_AOI22_X1 T1644 ( .Y(T1644_Y), .B1(T10346_Y), .B0(T6785_Q),     .A1(T15245_Y), .A0(T13898_Q));
KC_AOI22_X1 T1646 ( .Y(T1646_Y), .B1(T6785_Q), .B0(T10361_Y),     .A1(T13898_Q), .A0(T15247_Y));
KC_AOI22_X1 T1649 ( .Y(T1649_Y), .B1(T13887_Q), .B0(T10361_Y),     .A1(T13886_Q), .A0(T15247_Y));
KC_AOI22_X1 T1652 ( .Y(T1652_Y), .B1(T14058_Q), .B0(T10359_Y),     .A1(T14060_Q), .A0(T4889_Y));
KC_AOI22_X1 T7984 ( .Y(T7984_Y), .B1(T2038_Y), .B0(T1059_Y),     .A1(T4933_Y), .A0(T16413_Q));
KC_AOI22_X1 T7983 ( .Y(T7983_Y), .B1(T2038_Y), .B0(T15463_Y),     .A1(T4933_Y), .A0(T8877_Q));
KC_AOI22_X1 T7982 ( .Y(T7982_Y), .B1(T2038_Y), .B0(T1578_Y),     .A1(T4933_Y), .A0(T1719_Q));
KC_AOI22_X1 T7981 ( .Y(T7981_Y), .B1(T2038_Y), .B0(T1597_Y),     .A1(T4933_Y), .A0(T16433_Q));
KC_AOI22_X1 T7980 ( .Y(T7980_Y), .B1(T2038_Y), .B0(T975_Y),     .A1(T4933_Y), .A0(T1717_Q));
KC_AOI22_X1 T7924 ( .Y(T7924_Y), .B1(T2038_Y), .B0(T15660_Y),     .A1(T4933_Y), .A0(T1691_Q));
KC_AOI22_X1 T7923 ( .Y(T7923_Y), .B1(T2038_Y), .B0(T1456_Y),     .A1(T10525_Y), .A0(T8877_Q));
KC_AOI22_X1 T7922 ( .Y(T7922_Y), .B1(T2038_Y), .B0(T1471_Y),     .A1(T4933_Y), .A0(T1707_Q));
KC_AOI22_X1 T7921 ( .Y(T7921_Y), .B1(T2038_Y), .B0(T1709_Y),     .A1(T4933_Y), .A0(T8880_Q));
KC_AOI22_X1 T1686 ( .Y(T1686_Y), .B1(T2038_Y), .B0(T16440_Y),     .A1(T10525_Y), .A0(T5364_Q));
KC_AOI22_X1 T10702 ( .Y(T10702_Y), .B1(T2038_Y), .B0(T1058_Y),     .A1(T10525_Y), .A0(T8880_Q));
KC_AOI22_X1 T10701 ( .Y(T10701_Y), .B1(T2038_Y), .B0(T15531_Y),     .A1(T10525_Y), .A0(T1691_Q));
KC_AOI22_X1 T10700 ( .Y(T10700_Y), .B1(T2038_Y), .B0(T1472_Y),     .A1(T10525_Y), .A0(T1717_Q));
KC_AOI22_X1 T1749 ( .Y(T1749_Y), .B1(T5794_Y), .B0(T10207_Y),     .A1(T1750_Y), .A0(T15810_Y));
KC_AOI22_X1 T1784 ( .Y(T1784_Y), .B1(T1785_Q), .B0(T12269_Y),     .A1(T1806_Q), .A0(T12270_Y));
KC_AOI22_X1 T1794 ( .Y(T1794_Y), .B1(T1807_Q), .B0(T12269_Y),     .A1(T1790_Q), .A0(T6164_Y));
KC_AOI22_X1 T1795 ( .Y(T1795_Y), .B1(T1823_Q), .B0(T12269_Y),     .A1(T1787_Q), .A0(T6164_Y));
KC_AOI22_X1 T1796 ( .Y(T1796_Y), .B1(T1803_Q), .B0(T4965_Y),     .A1(T3784_Y), .A0(T12268_Y));
KC_AOI22_X1 T1798 ( .Y(T1798_Y), .B1(T1787_Q), .B0(T4965_Y),     .A1(T3304_Y), .A0(T12268_Y));
KC_AOI22_X1 T1799 ( .Y(T1799_Y), .B1(T1806_Q), .B0(T12269_Y),     .A1(T1803_Q), .A0(T12270_Y));
KC_AOI22_X1 T1800 ( .Y(T1800_Y), .B1(T1806_Q), .B0(T4965_Y),     .A1(T8354_Y), .A0(T12268_Y));
KC_AOI22_X1 T1801 ( .Y(T1801_Y), .B1(T1803_Q), .B0(T12269_Y),     .A1(T1787_Q), .A0(T12270_Y));
KC_AOI22_X1 T1802 ( .Y(T1802_Y), .B1(T1789_Q), .B0(T11728_Y),     .A1(T2876_Y), .A0(T5480_Q));
KC_AOI22_X1 T1808 ( .Y(T1808_Y), .B1(T1823_Q), .B0(T6164_Y),     .A1(T1789_Q), .A0(T12270_Y));
KC_AOI22_X1 T1809 ( .Y(T1809_Y), .B1(T4925_Q), .B0(T12269_Y),     .A1(T1806_Q), .A0(T6164_Y));
KC_AOI22_X1 T1811 ( .Y(T1811_Y), .B1(T4925_Q), .B0(T6164_Y),     .A1(T1821_Q), .A0(T12270_Y));
KC_AOI22_X1 T1812 ( .Y(T1812_Y), .B1(T1821_Q), .B0(T12269_Y),     .A1(T1826_Q), .A0(T6164_Y));
KC_AOI22_X1 T1817 ( .Y(T1817_Y), .B1(T5524_Q), .B0(T4965_Y),     .A1(T15990_Q), .A0(T2876_Y));
KC_AOI22_X1 T1819 ( .Y(T1819_Y), .B1(T1830_Q), .B0(T12269_Y),     .A1(T5524_Q), .A0(T12270_Y));
KC_AOI22_X1 T1858 ( .Y(T1858_Y), .B1(T9580_Y), .B0(T13415_Q),     .A1(T2027_Y), .A0(T13401_Q));
KC_AOI22_X1 T1859 ( .Y(T1859_Y), .B1(T9580_Y), .B0(T13414_Q),     .A1(T2027_Y), .A0(T13400_Q));
KC_AOI22_X1 T1860 ( .Y(T1860_Y), .B1(T13414_Q), .B0(T12075_Y),     .A1(T13400_Q), .A0(T7323_Y));
KC_AOI22_X1 T1861 ( .Y(T1861_Y), .B1(T13415_Q), .B0(T12075_Y),     .A1(T13401_Q), .A0(T7323_Y));
KC_AOI22_X1 T5726 ( .Y(T5726_Y), .B1(T6452_Y), .B0(T13538_Q),     .A1(T1632_Y), .A0(T13517_Q));
KC_AOI22_X1 T1872 ( .Y(T1872_Y), .B1(T12325_Y), .B0(T13537_Q),     .A1(T12324_Y), .A0(T13518_Q));
KC_AOI22_X1 T1876 ( .Y(T1876_Y), .B1(T6452_Y), .B0(T13561_Q),     .A1(T1632_Y), .A0(T13559_Q));
KC_AOI22_X1 T1877 ( .Y(T1877_Y), .B1(T13510_Q), .B0(T12077_Y),     .A1(T13544_Q), .A0(T12078_Y));
KC_AOI22_X1 T1878 ( .Y(T1878_Y), .B1(T13516_Q), .B0(T12076_Y),     .A1(T13513_Q), .A0(T12074_Y));
KC_AOI22_X1 T1879 ( .Y(T1879_Y), .B1(T6452_Y), .B0(T13510_Q),     .A1(T1632_Y), .A0(T13544_Q));
KC_AOI22_X1 T1880 ( .Y(T1880_Y), .B1(T6452_Y), .B0(T13512_Q),     .A1(T1632_Y), .A0(T13557_Q));
KC_AOI22_X1 T1881 ( .Y(T1881_Y), .B1(T13427_Q), .B0(T12076_Y),     .A1(T14818_Q), .A0(T12074_Y));
KC_AOI22_X1 T1882 ( .Y(T1882_Y), .B1(T6452_Y), .B0(T13562_Q),     .A1(T1632_Y), .A0(T13560_Q));
KC_AOI22_X1 T1883 ( .Y(T1883_Y), .B1(T12325_Y), .B0(T13516_Q),     .A1(T12324_Y), .A0(T13513_Q));
KC_AOI22_X1 T1884 ( .Y(T1884_Y), .B1(T13563_Q), .B0(T1547_Y),     .A1(T13536_Q), .A0(T15202_Y));
KC_AOI22_X1 T1887 ( .Y(T1887_Y), .B1(T13533_Q), .B0(T1547_Y),     .A1(T14805_Q), .A0(T15202_Y));
KC_AOI22_X1 T1888 ( .Y(T1888_Y), .B1(T13531_Q), .B0(T1547_Y),     .A1(T14803_Q), .A0(T15202_Y));
KC_AOI22_X1 T1889 ( .Y(T1889_Y), .B1(T13534_Q), .B0(T1547_Y),     .A1(T13535_Q), .A0(T15202_Y));
KC_AOI22_X1 T1890 ( .Y(T1890_Y), .B1(T13562_Q), .B0(T12077_Y),     .A1(T13560_Q), .A0(T12078_Y));
KC_AOI22_X1 T1891 ( .Y(T1891_Y), .B1(T13561_Q), .B0(T12077_Y),     .A1(T13559_Q), .A0(T12078_Y));
KC_AOI22_X1 T1893 ( .Y(T1893_Y), .B1(T10397_Y), .B0(T13533_Q),     .A1(T15204_Y), .A0(T14805_Q));
KC_AOI22_X1 T1894 ( .Y(T1894_Y), .B1(T10397_Y), .B0(T13534_Q),     .A1(T15204_Y), .A0(T13535_Q));
KC_AOI22_X1 T1895 ( .Y(T1895_Y), .B1(T12325_Y), .B0(T13427_Q),     .A1(T12324_Y), .A0(T14818_Q));
KC_AOI22_X1 T1896 ( .Y(T1896_Y), .B1(T13515_Q), .B0(T12076_Y),     .A1(T14817_Q), .A0(T12074_Y));
KC_AOI22_X1 T1897 ( .Y(T1897_Y), .B1(T13514_Q), .B0(T12076_Y),     .A1(T14819_Q), .A0(T12074_Y));
KC_AOI22_X1 T1898 ( .Y(T1898_Y), .B1(T12325_Y), .B0(T13514_Q),     .A1(T12324_Y), .A0(T14819_Q));
KC_AOI22_X1 T5739 ( .Y(T5739_Y), .B1(T14772_Q), .B0(T12075_Y),     .A1(T13660_Q), .A0(T7323_Y));
KC_AOI22_X1 T1900 ( .Y(T1900_Y), .B1(T13627_Q), .B0(T1547_Y),     .A1(T13628_Q), .A0(T15202_Y));
KC_AOI22_X1 T1901 ( .Y(T1901_Y), .B1(T14804_Q), .B0(T12076_Y),     .A1(T13678_Q), .A0(T12074_Y));
KC_AOI22_X1 T1902 ( .Y(T1902_Y), .B1(T13679_Q), .B0(T1547_Y),     .A1(T13629_Q), .A0(T15202_Y));
KC_AOI22_X1 T1903 ( .Y(T1903_Y), .B1(T12325_Y), .B0(T14784_Q),     .A1(T12324_Y), .A0(T13640_Q));
KC_AOI22_X1 T1904 ( .Y(T1904_Y), .B1(T12325_Y), .B0(T14804_Q),     .A1(T12324_Y), .A0(T13678_Q));
KC_AOI22_X1 T1905 ( .Y(T1905_Y), .B1(T14785_Q), .B0(T12076_Y),     .A1(T13680_Q), .A0(T12074_Y));
KC_AOI22_X1 T1906 ( .Y(T1906_Y), .B1(T12325_Y), .B0(T14785_Q),     .A1(T12324_Y), .A0(T13680_Q));
KC_AOI22_X1 T1907 ( .Y(T1907_Y), .B1(T13681_Q), .B0(T1547_Y),     .A1(T13631_Q), .A0(T15202_Y));
KC_AOI22_X1 T1908 ( .Y(T1908_Y), .B1(T13661_Q), .B0(T12075_Y),     .A1(T14770_Q), .A0(T7323_Y));
KC_AOI22_X1 T1909 ( .Y(T1909_Y), .B1(T9580_Y), .B0(T14772_Q),     .A1(T3640_Y), .A0(T13660_Q));
KC_AOI22_X1 T1910 ( .Y(T1910_Y), .B1(T14768_Q), .B0(T12075_Y),     .A1(T13658_Q), .A0(T7323_Y));
KC_AOI22_X1 T1911 ( .Y(T1911_Y), .B1(T9580_Y), .B0(T14768_Q),     .A1(T3640_Y), .A0(T13658_Q));
KC_AOI22_X1 T1912 ( .Y(T1912_Y), .B1(T9580_Y), .B0(T13661_Q),     .A1(T3640_Y), .A0(T14770_Q));
KC_AOI22_X1 T1915 ( .Y(T1915_Y), .B1(T14784_Q), .B0(T12076_Y),     .A1(T13640_Q), .A0(T12074_Y));
KC_AOI22_X1 T1919 ( .Y(T1919_Y), .B1(T10397_Y), .B0(T13681_Q),     .A1(T15204_Y), .A0(T13631_Q));
KC_AOI22_X1 T1920 ( .Y(T1920_Y), .B1(T10397_Y), .B0(T13679_Q),     .A1(T15204_Y), .A0(T13629_Q));
KC_AOI22_X1 T1921 ( .Y(T1921_Y), .B1(T10397_Y), .B0(T13627_Q),     .A1(T15204_Y), .A0(T13628_Q));
KC_AOI22_X1 T1922 ( .Y(T1922_Y), .B1(T6452_Y), .B0(T14786_Q),     .A1(T1632_Y), .A0(T14787_Q));
KC_AOI22_X1 T1923 ( .Y(T1923_Y), .B1(T14786_Q), .B0(T12077_Y),     .A1(T14787_Q), .A0(T12078_Y));
KC_AOI22_X1 T1924 ( .Y(T1924_Y), .B1(T6452_Y), .B0(T14806_Q),     .A1(T1632_Y), .A0(T14807_Q));
KC_AOI22_X1 T1925 ( .Y(T1925_Y), .B1(T14806_Q), .B0(T12077_Y),     .A1(T14807_Q), .A0(T12078_Y));
KC_AOI22_X1 T1926 ( .Y(T1926_Y), .B1(T14788_Q), .B0(T12077_Y),     .A1(T14808_Q), .A0(T12078_Y));
KC_AOI22_X1 T1927 ( .Y(T1927_Y), .B1(T6452_Y), .B0(T14788_Q),     .A1(T1632_Y), .A0(T14808_Q));
KC_AOI22_X1 T1928 ( .Y(T1928_Y), .B1(T14810_Q), .B0(T12077_Y),     .A1(T14811_Q), .A0(T12078_Y));
KC_AOI22_X1 T6679 ( .Y(T6679_Y), .B1(T9704_Y), .B0(T14072_Q),     .A1(T9705_Y), .A0(T14070_Q));
KC_AOI22_X1 T6678 ( .Y(T6678_Y), .B1(T14072_Q), .B0(T10358_Y),     .A1(T14070_Q), .A0(T9712_Y));
KC_AOI22_X1 T5797 ( .Y(T5797_Y), .B1(T13884_Q), .B0(T10362_Y),     .A1(T14861_Q), .A0(T10360_Y));
KC_AOI22_X1 T1932 ( .Y(T1932_Y), .B1(T9704_Y), .B0(T14055_Q),     .A1(T9705_Y), .A0(T14057_Q));
KC_AOI22_X1 T1933 ( .Y(T1933_Y), .B1(T14054_Q), .B0(T10358_Y),     .A1(T14056_Q), .A0(T9712_Y));
KC_AOI22_X1 T1934 ( .Y(T1934_Y), .B1(T9704_Y), .B0(T14054_Q),     .A1(T9705_Y), .A0(T14056_Q));
KC_AOI22_X1 T1935 ( .Y(T1935_Y), .B1(T14055_Q), .B0(T10358_Y),     .A1(T14057_Q), .A0(T9712_Y));
KC_AOI22_X1 T1936 ( .Y(T1936_Y), .B1(T9704_Y), .B0(T14073_Q),     .A1(T9705_Y), .A0(T14052_Q));
KC_AOI22_X1 T1942 ( .Y(T1942_Y), .B1(T9707_Y), .B0(T13883_Q),     .A1(T10347_Y), .A0(T13930_Q));
KC_AOI22_X1 T1943 ( .Y(T1943_Y), .B1(T9707_Y), .B0(T13884_Q),     .A1(T10347_Y), .A0(T14861_Q));
KC_AOI22_X1 T1944 ( .Y(T1944_Y), .B1(T9707_Y), .B0(T13882_Q),     .A1(T10347_Y), .A0(T14863_Q));
KC_AOI22_X1 T1945 ( .Y(T1945_Y), .B1(T9707_Y), .B0(T13885_Q),     .A1(T10347_Y), .A0(T14860_Q));
KC_AOI22_X1 T1946 ( .Y(T1946_Y), .B1(T10346_Y), .B0(T13915_Q),     .A1(T15245_Y), .A0(T13914_Q));
KC_AOI22_X1 T1947 ( .Y(T1947_Y), .B1(T13917_Q), .B0(T10361_Y),     .A1(T13918_Q), .A0(T15247_Y));
KC_AOI22_X1 T1948 ( .Y(T1948_Y), .B1(T13915_Q), .B0(T10361_Y),     .A1(T13914_Q), .A0(T15247_Y));
KC_AOI22_X1 T1951 ( .Y(T1951_Y), .B1(T10346_Y), .B0(T13919_Q),     .A1(T15245_Y), .A0(T13897_Q));
KC_AOI22_X1 T1952 ( .Y(T1952_Y), .B1(T13883_Q), .B0(T10362_Y),     .A1(T13930_Q), .A0(T10360_Y));
KC_AOI22_X1 T1953 ( .Y(T1953_Y), .B1(T13885_Q), .B0(T10362_Y),     .A1(T14860_Q), .A0(T10360_Y));
KC_AOI22_X1 T1954 ( .Y(T1954_Y), .B1(T13882_Q), .B0(T10362_Y),     .A1(T14863_Q), .A0(T10360_Y));
KC_AOI22_X1 T1955 ( .Y(T1955_Y), .B1(T13919_Q), .B0(T10361_Y),     .A1(T13897_Q), .A0(T15247_Y));
KC_AOI22_X1 T1956 ( .Y(T1956_Y), .B1(T10346_Y), .B0(T13916_Q),     .A1(T15245_Y), .A0(T13920_Q));
KC_AOI22_X1 T1957 ( .Y(T1957_Y), .B1(T10346_Y), .B0(T13917_Q),     .A1(T15245_Y), .A0(T13918_Q));
KC_AOI22_X1 T1958 ( .Y(T1958_Y), .B1(T13916_Q), .B0(T10361_Y),     .A1(T13920_Q), .A0(T15247_Y));
KC_AOI22_X1 T1967 ( .Y(T1967_Y), .B1(T9706_Y), .B0(T14058_Q),     .A1(T1545_Y), .A0(T14060_Q));
KC_AOI22_X1 T1968 ( .Y(T1968_Y), .B1(T14071_Q), .B0(T10359_Y),     .A1(T14059_Q), .A0(T4889_Y));
KC_AOI22_X1 T1969 ( .Y(T1969_Y), .B1(T14073_Q), .B0(T10358_Y),     .A1(T14052_Q), .A0(T9712_Y));
KC_AOI22_X1 T1989 ( .Y(T1989_Y), .B1(T2038_Y), .B0(T16271_Y),     .A1(T4933_Y), .A0(T5362_Q));
KC_AOI22_X1 T2041 ( .Y(T2041_Y), .B1(T9974_Y), .B0(T10100_Y),     .A1(T1987_Y), .A0(T16411_Y));
KC_AOI22_X1 T2084 ( .Y(T2084_Y), .B1(T2689_Q), .B0(T5848_Y),     .A1(T16482_Q), .A0(T11499_Y));
KC_AOI22_X1 T2085 ( .Y(T2085_Y), .B1(T13065_Q), .B0(T12248_Y),     .A1(T15828_Q), .A0(T11499_Y));
KC_AOI22_X1 T2086 ( .Y(T2086_Y), .B1(T5434_Q), .B0(T5909_Y),     .A1(T2089_Q), .A0(T11499_Y));
KC_AOI22_X1 T2087 ( .Y(T2087_Y), .B1(T16483_Q), .B0(T12248_Y),     .A1(T2095_Q), .A0(T5909_Y));
KC_AOI22_X1 T2101 ( .Y(T2101_Y), .B1(T5848_Y), .B0(T15879_Q),     .A1(T1746_Y), .A0(T11499_Y));
KC_AOI22_X1 T2102 ( .Y(T2102_Y), .B1(T4969_Q), .B0(T5909_Y),     .A1(T5574_Q), .A0(T5848_Y));
KC_AOI22_X1 T2108 ( .Y(T2108_Y), .B1(T15894_Q), .B0(T5848_Y),     .A1(T11480_Y), .A0(T8446_Y));
KC_AOI22_X1 T2135 ( .Y(T2135_Y), .B1(T2151_Q), .B0(T5944_Y),     .A1(T5452_Q), .A0(T11641_Y));
KC_AOI22_X1 T2136 ( .Y(T2136_Y), .B1(T5438_Q), .B0(T5909_Y),     .A1(T13132_Q), .A0(T11604_Y));
KC_AOI22_X1 T2137 ( .Y(T2137_Y), .B1(T14968_Y), .B0(T12248_Y),     .A1(T11480_Y), .A0(T2739_Y));
KC_AOI22_X1 T2138 ( .Y(T2138_Y), .B1(T4924_Q), .B0(T12248_Y),     .A1(T1761_Q), .A0(T5944_Y));
KC_AOI22_X1 T2139 ( .Y(T2139_Y), .B1(T5944_Y), .B0(T2162_Q),     .A1(T2150_Q), .A0(T11641_Y));
KC_AOI22_X1 T2142 ( .Y(T2142_Y), .B1(T1758_Q), .B0(T12248_Y),     .A1(T11480_Y), .A0(T2740_Y));
KC_AOI22_X1 T2143 ( .Y(T2143_Y), .B1(T2160_Q), .B0(T5944_Y),     .A1(T2119_Q), .A0(T11604_Y));
KC_AOI22_X1 T2144 ( .Y(T2144_Y), .B1(T13102_Q), .B0(T12248_Y),     .A1(T1760_Q), .A0(T11641_Y));
KC_AOI22_X1 T2147 ( .Y(T2147_Y), .B1(T5442_Q), .B0(T5909_Y),     .A1(T2152_Q), .A0(T11604_Y));
KC_AOI22_X1 T2174 ( .Y(T2174_Y), .B1(T2118_Q), .B0(T11620_Y),     .A1(T11435_Y), .A0(T11551_Y));
KC_AOI22_X1 T15983 ( .Y(T15983_Y), .B1(T2212_Y), .B0(T5987_Q),     .A1(T2792_Y), .A0(T16098_Y));
KC_AOI22_X1 T6302 ( .Y(T6302_Y), .B1(T4967_Q), .B0(T11586_Y),     .A1(T5480_Q), .A0(T5990_Y));
KC_AOI22_X1 T6301 ( .Y(T6301_Y), .B1(T5474_Q), .B0(T11620_Y),     .A1(T16071_Y), .A0(T15232_Y));
KC_AOI22_X1 T2190 ( .Y(T2190_Y), .B1(T16235_Y), .B0(T15232_Y),     .A1(T2809_Q), .A0(T5990_Y));
KC_AOI22_X1 T2192 ( .Y(T2192_Y), .B1(T2670_Y), .B0(T6015_Y),     .A1(T16075_Y), .A0(T15232_Y));
KC_AOI22_X1 T2193 ( .Y(T2193_Y), .B1(T16076_Y), .B0(T15232_Y),     .A1(T2281_Q), .A0(T5990_Y));
KC_AOI22_X1 T2194 ( .Y(T2194_Y), .B1(T16069_Y), .B0(T6015_Y),     .A1(T16074_Y), .A0(T15232_Y));
KC_AOI22_X1 T2195 ( .Y(T2195_Y), .B1(T1777_Q), .B0(T11620_Y),     .A1(T2249_Q), .A0(T5990_Y));
KC_AOI22_X1 T2196 ( .Y(T2196_Y), .B1(T2236_Q), .B0(T5990_Y),     .A1(T8249_Y), .A0(T11551_Y));
KC_AOI22_X1 T2197 ( .Y(T2197_Y), .B1(T16076_Y), .B0(T6015_Y),     .A1(T2141_Y), .A0(T11551_Y));
KC_AOI22_X1 T2198 ( .Y(T2198_Y), .B1(T2276_Q), .B0(T11586_Y),     .A1(T16069_Y), .A0(T15232_Y));
KC_AOI22_X1 T2201 ( .Y(T2201_Y), .B1(T5473_Q), .B0(T11620_Y),     .A1(T2670_Y), .A0(T15232_Y));
KC_AOI22_X1 T2202 ( .Y(T2202_Y), .B1(T6071_Q), .B0(T11620_Y),     .A1(T9162_Y), .A0(T15232_Y));
KC_AOI22_X1 T2203 ( .Y(T2203_Y), .B1(T1778_Q), .B0(T11620_Y),     .A1(T16070_Y), .A0(T15232_Y));
KC_AOI22_X1 T2204 ( .Y(T2204_Y), .B1(T1775_Q), .B0(T11586_Y),     .A1(T2835_Q), .A0(T5990_Y));
KC_AOI22_X1 T2208 ( .Y(T2208_Y), .B1(T16235_Y), .B0(T6015_Y),     .A1(T12028_Y), .A0(T13129_Q));
KC_AOI22_X1 T2209 ( .Y(T2209_Y), .B1(T5471_Y), .B0(T16097_Y),     .A1(T2851_Y), .A0(T12102_Y));
KC_AOI22_X1 T2210 ( .Y(T2210_Y), .B1(T1774_Q), .B0(T11620_Y),     .A1(T1779_Q), .A0(T11586_Y));
KC_AOI22_X1 T2211 ( .Y(T2211_Y), .B1(T16098_Y), .B0(T15232_Y),     .A1(T12028_Y), .A0(T13136_Q));
KC_AOI22_X1 T2221 ( .Y(T2221_Y), .B1(T4960_Y), .B0(T6070_Y),     .A1(T11613_Y), .A0(T2220_Y));
KC_AOI22_X1 T2222 ( .Y(T2222_Y), .B1(T2218_Y), .B0(T6070_Y),     .A1(T11613_Y), .A0(T2207_Y));
KC_AOI22_X1 T2223 ( .Y(T2223_Y), .B1(T2191_Y), .B0(T6070_Y),     .A1(T11613_Y), .A0(T8340_Y));
KC_AOI22_X1 T2224 ( .Y(T2224_Y), .B1(T6003_Y), .B0(T12106_Y),     .A1(T2851_Y), .A0(T12108_Y));
KC_AOI22_X1 T2225 ( .Y(T2225_Y), .B1(T16073_Y), .B0(T6015_Y),     .A1(T16010_Q), .A0(T5990_Y));
KC_AOI22_X1 T2226 ( .Y(T2226_Y), .B1(T16096_Y), .B0(T15232_Y),     .A1(T6073_Y), .A0(T12106_Y));
KC_AOI22_X1 T2232 ( .Y(T2232_Y), .B1(T8471_Y), .B0(T11613_Y),     .A1(T11727_Y), .A0(T5494_Q));
KC_AOI22_X1 T2233 ( .Y(T2233_Y), .B1(T6214_Y), .B0(T5571_Q),     .A1(T6003_Y), .A0(T12102_Y));
KC_AOI22_X1 T2234 ( .Y(T2234_Y), .B1(T6214_Y), .B0(T2311_Q),     .A1(T6003_Y), .A0(T16270_Y));
KC_AOI22_X1 T2235 ( .Y(T2235_Y), .B1(T2200_Y), .B0(T11613_Y),     .A1(T11727_Y), .A0(T8352_Q));
KC_AOI22_X1 T2252 ( .Y(T2252_Y), .B1(T6464_Y), .B0(T2278_Q),     .A1(T12270_Y), .A0(T2345_Q));
KC_AOI22_X1 T2253 ( .Y(T2253_Y), .B1(T6464_Y), .B0(T8352_Q),     .A1(T12270_Y), .A0(T15138_Q));
KC_AOI22_X1 T2254 ( .Y(T2254_Y), .B1(T6464_Y), .B0(T15138_Q),     .A1(T12270_Y), .A0(T2278_Q));
KC_AOI22_X1 T2255 ( .Y(T2255_Y), .B1(T2819_Y), .B0(T16007_Q),     .A1(T6164_Y), .A0(T15138_Q));
KC_AOI22_X1 T2257 ( .Y(T2257_Y), .B1(T8374_Y), .B0(T12268_Y),     .A1(T11728_Y), .A0(T4964_Q));
KC_AOI22_X1 T2258 ( .Y(T2258_Y), .B1(T8363_Y), .B0(T12268_Y),     .A1(T4965_Y), .A0(T2314_Q));
KC_AOI22_X1 T2265 ( .Y(T2265_Y), .B1(T2819_Y), .B0(T16018_Q),     .A1(T6164_Y), .A0(T8352_Q));
KC_AOI22_X1 T2269 ( .Y(T2269_Y), .B1(T2819_Y), .B0(T16010_Q),     .A1(T6164_Y), .A0(T16082_Q));
KC_AOI22_X1 T2270 ( .Y(T2270_Y), .B1(T2819_Y), .B0(T5987_Q),     .A1(T6164_Y), .A0(T2278_Q));
KC_AOI22_X1 T2272 ( .Y(T2272_Y), .B1(T2236_Q), .B0(T2876_Y),     .A1(T11728_Y), .A0(T8352_Q));
KC_AOI22_X1 T2273 ( .Y(T2273_Y), .B1(T5481_Q), .B0(T2876_Y),     .A1(T11728_Y), .A0(T15138_Q));
KC_AOI22_X1 T2285 ( .Y(T2285_Y), .B1(T8402_Y), .B0(T12268_Y),     .A1(T6164_Y), .A0(T2314_Q));
KC_AOI22_X1 T2286 ( .Y(T2286_Y), .B1(T2687_Y), .B0(T12268_Y),     .A1(T4965_Y), .A0(T2315_Q));
KC_AOI22_X1 T2287 ( .Y(T2287_Y), .B1(T2295_Y), .B0(T12268_Y),     .A1(T6164_Y), .A0(T4964_Q));
KC_AOI22_X1 T2288 ( .Y(T2288_Y), .B1(T3079_Y), .B0(T12268_Y),     .A1(T4965_Y), .A0(T5494_Q));
KC_AOI22_X1 T2289 ( .Y(T2289_Y), .B1(T12270_Y), .B0(T6419_Q),     .A1(T12269_Y), .A0(T2313_Q));
KC_AOI22_X1 T2290 ( .Y(T2290_Y), .B1(T12270_Y), .B0(T4964_Q),     .A1(T6464_Y), .A0(T2345_Q));
KC_AOI22_X1 T2291 ( .Y(T2291_Y), .B1(T8400_Y), .B0(T12268_Y),     .A1(T4965_Y), .A0(T6419_Q));
KC_AOI22_X1 T2292 ( .Y(T2292_Y), .B1(T6464_Y), .B0(T2314_Q),     .A1(T12270_Y), .A0(T2315_Q));
KC_AOI22_X1 T2296 ( .Y(T2296_Y), .B1(T2398_Y), .B0(T12268_Y),     .A1(T6164_Y), .A0(T2345_Q));
KC_AOI22_X1 T2297 ( .Y(T2297_Y), .B1(T6070_Y), .B0(T6147_Y),     .A1(T2316_Q), .A0(T6164_Y));
KC_AOI22_X1 T2302 ( .Y(T2302_Y), .B1(T8388_Y), .B0(T12268_Y),     .A1(T4965_Y), .A0(T2311_Q));
KC_AOI22_X1 T2303 ( .Y(T2303_Y), .B1(T6464_Y), .B0(T4964_Q),     .A1(T10593_Y), .A0(T2316_Q));
KC_AOI22_X1 T2305 ( .Y(T2305_Y), .B1(T2574_Y), .B0(T12268_Y),     .A1(T4965_Y), .A0(T2313_Q));
KC_AOI22_X1 T2306 ( .Y(T2306_Y), .B1(T10593_Y), .B0(T2314_Q),     .A1(T6464_Y), .A0(T2316_Q));
KC_AOI22_X1 T2307 ( .Y(T2307_Y), .B1(T5526_Q), .B0(T12269_Y),     .A1(T1829_Q), .A0(T10593_Y));
KC_AOI22_X1 T2308 ( .Y(T2308_Y), .B1(T2353_Q), .B0(T12269_Y),     .A1(T5566_Q), .A0(T10593_Y));
KC_AOI22_X1 T2330 ( .Y(T2330_Y), .B1(T11774_Y), .B0(T2354_Y),     .A1(T2329_Y), .A0(T12101_Y));
KC_AOI22_X1 T2337 ( .Y(T2337_Y), .B1(T2333_Y), .B0(T2335_Y),     .A1(T6523_Y), .A0(T11775_Y));
KC_AOI22_X1 T2402 ( .Y(T2402_Y), .B1(T12325_Y), .B0(T13515_Q),     .A1(T12324_Y), .A0(T14817_Q));
KC_AOI22_X1 T2403 ( .Y(T2403_Y), .B1(T3027_Y), .B0(T14815_Q),     .A1(T9636_Y), .A0(T13395_Q));
KC_AOI22_X1 T2404 ( .Y(T2404_Y), .B1(T3027_Y), .B0(T14816_Q),     .A1(T9636_Y), .A0(T13410_Q));
KC_AOI22_X1 T2405 ( .Y(T2405_Y), .B1(T3027_Y), .B0(T13399_Q),     .A1(T9636_Y), .A0(T13413_Q));
KC_AOI22_X1 T2406 ( .Y(T2406_Y), .B1(T14816_Q), .B0(T3611_Y),     .A1(T13410_Q), .A0(T6482_Y));
KC_AOI22_X1 T2407 ( .Y(T2407_Y), .B1(T13399_Q), .B0(T3611_Y),     .A1(T13413_Q), .A0(T6482_Y));
KC_AOI22_X1 T2410 ( .Y(T2410_Y), .B1(T10387_Y), .B0(T2535_Y),     .A1(T2990_Y), .A0(T2532_Y));
KC_AOI22_X1 T2411 ( .Y(T2411_Y), .B1(T6981_Y), .B0(T2535_Y),     .A1(T2985_Y), .A0(T2532_Y));
KC_AOI22_X1 T2413 ( .Y(T2413_Y), .B1(T13512_Q), .B0(T12077_Y),     .A1(T13557_Q), .A0(T12078_Y));
KC_AOI22_X1 T2414 ( .Y(T2414_Y), .B1(T1875_Y), .B0(T2535_Y),     .A1(T3564_Y), .A0(T2532_Y));
KC_AOI22_X1 T2415 ( .Y(T2415_Y), .B1(T10436_Y), .B0(T13528_Q),     .A1(T10437_Y), .A0(T13543_Q));
KC_AOI22_X1 T2416 ( .Y(T2416_Y), .B1(T13528_Q), .B0(T9637_Y),     .A1(T13543_Q), .A0(T6483_Y));
KC_AOI22_X1 T2417 ( .Y(T2417_Y), .B1(T1873_Y), .B0(T2535_Y),     .A1(T3566_Y), .A0(T2532_Y));
KC_AOI22_X1 T2418 ( .Y(T2418_Y), .B1(T1622_Y), .B0(T2535_Y),     .A1(T2426_Y), .A0(T2532_Y));
KC_AOI22_X1 T2419 ( .Y(T2419_Y), .B1(T10436_Y), .B0(T13558_Q),     .A1(T10437_Y), .A0(T13511_Q));
KC_AOI22_X1 T2420 ( .Y(T2420_Y), .B1(T10436_Y), .B0(T14800_Q),     .A1(T10437_Y), .A0(T13556_Q));
KC_AOI22_X1 T2421 ( .Y(T2421_Y), .B1(T1874_Y), .B0(T2535_Y),     .A1(T3548_Y), .A0(T2532_Y));
KC_AOI22_X1 T2422 ( .Y(T2422_Y), .B1(T10397_Y), .B0(T13531_Q),     .A1(T15204_Y), .A0(T14803_Q));
KC_AOI22_X1 T2423 ( .Y(T2423_Y), .B1(T7038_Y), .B0(T2535_Y),     .A1(T2980_Y), .A0(T2532_Y));
KC_AOI22_X1 T2424 ( .Y(T2424_Y), .B1(T10397_Y), .B0(T13530_Q),     .A1(T15204_Y), .A0(T13532_Q));
KC_AOI22_X1 T2427 ( .Y(T2427_Y), .B1(T13558_Q), .B0(T9637_Y),     .A1(T13511_Q), .A0(T6483_Y));
KC_AOI22_X1 T2428 ( .Y(T2428_Y), .B1(T6633_Y), .B0(T14765_Q),     .A1(T3579_Y), .A0(T4937_Y));
KC_AOI22_X1 T2429 ( .Y(T2429_Y), .B1(T6632_Y), .B0(T13656_Q),     .A1(T7219_Y), .A0(T4937_Y));
KC_AOI22_X1 T2430 ( .Y(T2430_Y), .B1(T1918_Y), .B0(T2535_Y),     .A1(T3000_Y), .A0(T2532_Y));
KC_AOI22_X1 T2431 ( .Y(T2431_Y), .B1(T1917_Y), .B0(T2535_Y),     .A1(T3578_Y), .A0(T2532_Y));
KC_AOI22_X1 T2432 ( .Y(T2432_Y), .B1(T1916_Y), .B0(T2535_Y),     .A1(T2425_Y), .A0(T2532_Y));
KC_AOI22_X1 T2433 ( .Y(T2433_Y), .B1(T1627_Y), .B0(T2535_Y),     .A1(T5034_Y), .A0(T2532_Y));
KC_AOI22_X1 T2456 ( .Y(T2456_Y), .B1(T7482_Y), .B0(T2531_Y),     .A1(T3655_Y), .A0(T16165_Y));
KC_AOI22_X1 T2462 ( .Y(T2462_Y), .B1(T1937_Y), .B0(T2531_Y),     .A1(T3617_Y), .A0(T16165_Y));
KC_AOI22_X1 T2463 ( .Y(T2463_Y), .B1(T1940_Y), .B0(T2531_Y),     .A1(T4232_Y), .A0(T16165_Y));
KC_AOI22_X1 T2471 ( .Y(T2471_Y), .B1(T1647_Y), .B0(T2531_Y),     .A1(T3622_Y), .A0(T16165_Y));
KC_AOI22_X1 T2472 ( .Y(T2472_Y), .B1(T7528_Y), .B0(T2531_Y),     .A1(T5084_Y), .A0(T16165_Y));
KC_AOI22_X1 T2473 ( .Y(T2473_Y), .B1(T1640_Y), .B0(T2531_Y),     .A1(T4240_Y), .A0(T16165_Y));
KC_AOI22_X1 T2479 ( .Y(T2479_Y), .B1(T4937_Y), .B0(T3605_Y),     .A1(T5805_Y), .A0(T13835_Q));
KC_AOI22_X1 T2486 ( .Y(T2486_Y), .B1(T1931_Y), .B0(T2531_Y),     .A1(T4251_Y), .A0(T16165_Y));
KC_AOI22_X1 T2487 ( .Y(T2487_Y), .B1(T1938_Y), .B0(T2531_Y),     .A1(T3628_Y), .A0(T16165_Y));
KC_AOI22_X1 T5850 ( .Y(T5850_Y), .B1(T3656_Y), .B0(T14994_Y),     .A1(T5841_Y), .A0(T14859_Q));
KC_AOI22_X1 T2499 ( .Y(T2499_Y), .B1(T6682_Y), .B0(T14151_Q),     .A1(T5083_Y), .A0(T14994_Y));
KC_AOI22_X1 T2506 ( .Y(T2506_Y), .B1(T5847_Y), .B0(T14081_Q),     .A1(T3627_Y), .A0(T14994_Y));
KC_AOI22_X1 T2510 ( .Y(T2510_Y), .B1(T5839_Y), .B0(T14083_Q),     .A1(T4250_Y), .A0(T14994_Y));
KC_AOI22_X1 T2517 ( .Y(T2517_Y), .B1(T7721_Y), .B0(T2531_Y),     .A1(T3670_Y), .A0(T16165_Y));
KC_AOI22_X1 T2518 ( .Y(T2518_Y), .B1(T7753_Y), .B0(T2531_Y),     .A1(T5327_Y), .A0(T16165_Y));
KC_AOI22_X1 T2519 ( .Y(T2519_Y), .B1(T7754_Y), .B0(T2531_Y),     .A1(T5882_Y), .A0(T16165_Y));
KC_AOI22_X1 T2546 ( .Y(T2546_Y), .B1(T3171_Y), .B0(T15218_Y),     .A1(T10034_Y), .A0(T15221_Y));
KC_AOI22_X1 T2552 ( .Y(T2552_Y), .B1(T5886_Y), .B0(T15072_Q),     .A1(T4291_Y), .A0(T2565_Y));
KC_AOI22_X1 T2553 ( .Y(T2553_Y), .B1(T3138_Y), .B0(T15218_Y),     .A1(T10038_Y), .A0(T15221_Y));
KC_AOI22_X1 T2554 ( .Y(T2554_Y), .B1(T5883_Y), .B0(T14892_Q),     .A1(T5322_Y), .A0(T14994_Y));
KC_AOI22_X1 T2555 ( .Y(T2555_Y), .B1(T3145_Y), .B0(T15218_Y),     .A1(T7944_Y), .A0(T15221_Y));
KC_AOI22_X1 T2556 ( .Y(T2556_Y), .B1(T3692_Y), .B0(T9946_Y),     .A1(T2549_Y), .A0(T2548_Y));
KC_AOI22_X1 T2557 ( .Y(T2557_Y), .B1(T3103_Y), .B0(T9946_Y),     .A1(T2549_Y), .A0(T2559_Y));
KC_AOI22_X1 T2563 ( .Y(T2563_Y), .B1(T5864_Y), .B0(T14882_Q),     .A1(T12089_Y), .A0(T14994_Y));
KC_AOI22_X1 T2568 ( .Y(T2568_Y), .B1(T4307_Y), .B0(T9946_Y),     .A1(T2549_Y), .A0(T2558_Y));
KC_AOI22_X1 T2569 ( .Y(T2569_Y), .B1(T5856_Y), .B0(T14152_Q),     .A1(T14994_Y), .A0(T4307_Y));
KC_AOI22_X1 T2594 ( .Y(T2594_Y), .B1(T3130_Y), .B0(T15218_Y),     .A1(T9980_Y), .A0(T15221_Y));
KC_AOI22_X1 T2595 ( .Y(T2595_Y), .B1(T5935_Y), .B0(T14345_Q),     .A1(T3741_Y), .A0(T2565_Y));
KC_AOI22_X1 T2600 ( .Y(T2600_Y), .B1(T3176_Y), .B0(T15218_Y),     .A1(T9989_Y), .A0(T15221_Y));
KC_AOI22_X1 T2601 ( .Y(T2601_Y), .B1(T16258_Y), .B0(T15218_Y),     .A1(T9996_Y), .A0(T15221_Y));
KC_AOI22_X1 T2602 ( .Y(T2602_Y), .B1(T3738_Y), .B0(T15218_Y),     .A1(T9990_Y), .A0(T15221_Y));
KC_AOI22_X1 T2603 ( .Y(T2603_Y), .B1(T3760_Y), .B0(T15218_Y),     .A1(T9993_Y), .A0(T15221_Y));
KC_AOI22_X1 T2605 ( .Y(T2605_Y), .B1(T3740_Y), .B0(T15218_Y),     .A1(T10035_Y), .A0(T15221_Y));
KC_AOI22_X1 T2606 ( .Y(T2606_Y), .B1(T3167_Y), .B0(T15218_Y),     .A1(T9991_Y), .A0(T15221_Y));
KC_AOI22_X1 T2607 ( .Y(T2607_Y), .B1(T2361_Q), .B0(T15518_Y),     .A1(T2621_Y), .A0(T2957_Y));
KC_AOI22_X1 T2615 ( .Y(T2615_Y), .B1(T2832_Q), .B0(T15518_Y),     .A1(T2628_Q), .A0(T2550_Y));
KC_AOI22_X1 T2616 ( .Y(T2616_Y), .B1(T3762_Y), .B0(T15218_Y),     .A1(T10011_Y), .A0(T15221_Y));
KC_AOI22_X1 T2617 ( .Y(T2617_Y), .B1(T3750_Y), .B0(T15218_Y),     .A1(T10307_Y), .A0(T15221_Y));
KC_AOI22_X1 T2634 ( .Y(T2634_Y), .B1(T5959_Y), .B0(T14425_Q),     .A1(T3166_Y), .A0(T2565_Y));
KC_AOI22_X1 T2635 ( .Y(T2635_Y), .B1(T5960_Y), .B0(T14427_Q),     .A1(T2565_Y), .A0(T3177_Y));
KC_AOI22_X1 T2636 ( .Y(T2636_Y), .B1(T3763_Y), .B0(T2565_Y),     .A1(T5962_Y), .A0(T14403_Q));
KC_AOI22_X1 T2637 ( .Y(T2637_Y), .B1(T5961_Y), .B0(T14426_Q),     .A1(T2565_Y), .A0(T3692_Y));
KC_AOI22_X1 T2638 ( .Y(T2638_Y), .B1(T5950_Y), .B0(T14363_Q),     .A1(T3742_Y), .A0(T2565_Y));
KC_AOI22_X1 T2657 ( .Y(T2657_Y), .B1(T2664_Y), .B0(T10280_Y),     .A1(T10251_Y), .A0(T14522_Q));
KC_AOI22_X1 T2659 ( .Y(T2659_Y), .B1(T10244_Y), .B0(T15815_Q),     .A1(T10251_Y), .A0(T14984_Y));
KC_AOI22_X1 T2730 ( .Y(T2730_Y), .B1(T6133_S), .B0(T6133_S),     .A1(T2750_Y), .A0(T5861_Y));
KC_AOI22_X1 T2733 ( .Y(T2733_Y), .B1(T8238_Y), .B0(T2735_Q),     .A1(T15582_Y), .A0(T11604_Y));
KC_AOI22_X1 T2756 ( .Y(T2756_Y), .B1(T15582_Y), .B0(T5944_Y),     .A1(T8238_Y), .A0(T2746_Q));
KC_AOI22_X1 T2769 ( .Y(T2769_Y), .B1(T8277_Y), .B0(T12009_Y),     .A1(T5069_Y), .A0(T15798_Q));
KC_AOI22_X1 T2771 ( .Y(T2771_Y), .B1(T8489_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T16301_Q));
KC_AOI22_X1 T2772 ( .Y(T2772_Y), .B1(T8491_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T16299_Q));
KC_AOI22_X1 T2773 ( .Y(T2773_Y), .B1(T8293_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T16088_Q));
KC_AOI22_X1 T2774 ( .Y(T2774_Y), .B1(T8260_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T15844_Q));
KC_AOI22_X1 T2775 ( .Y(T2775_Y), .B1(T8285_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T15803_Q));
KC_AOI22_X1 T2776 ( .Y(T2776_Y), .B1(T8294_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T15807_Q));
KC_AOI22_X1 T2780 ( .Y(T2780_Y), .B1(T8295_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T15809_Q));
KC_AOI22_X1 T2781 ( .Y(T2781_Y), .B1(T8276_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T15796_Q));
KC_AOI22_X1 T2795 ( .Y(T2795_Y), .B1(T2814_Q), .B0(T11620_Y),     .A1(T12028_Y), .A0(T13133_Q));
KC_AOI22_X1 T2796 ( .Y(T2796_Y), .B1(T11620_Y), .B0(T2833_Q),     .A1(T2851_Y), .A0(T12106_Y));
KC_AOI22_X1 T2799 ( .Y(T2799_Y), .B1(T8279_Y), .B0(T12009_Y),     .A1(T12008_Y), .A0(T15808_Q));
KC_AOI22_X1 T2801 ( .Y(T2801_Y), .B1(T5072_Y), .B0(T3411_Y),     .A1(T2803_Y), .A0(T15942_Y));
KC_AOI22_X1 T2828 ( .Y(T2828_Y), .B1(T8308_Y), .B0(T11613_Y),     .A1(T11727_Y), .A0(T5497_Q));
KC_AOI22_X1 T2829 ( .Y(T2829_Y), .B1(T6040_Y), .B0(T15942_Y),     .A1(T16156_Y), .A0(T6086_Y));
KC_AOI22_X1 T2853 ( .Y(T2853_Y), .B1(T10592_Y), .B0(T12105_Y),     .A1(T12038_Y), .A0(T10581_Y));
KC_AOI22_X1 T2858 ( .Y(T2858_Y), .B1(T10607_Y), .B0(T16100_Y),     .A1(T12038_Y), .A0(T15621_Y));
KC_AOI22_X1 T2863 ( .Y(T2863_Y), .B1(T2800_Y), .B0(T10607_Y),     .A1(T11598_Y), .A0(T11743_Y));
KC_AOI22_X1 T2864 ( .Y(T2864_Y), .B1(T16121_Y), .B0(T12048_Y),     .A1(T8378_Y), .A0(T6221_Y));
KC_AOI22_X1 T2895 ( .Y(T2895_Y), .B1(T2902_Y), .B0(T11742_Y),     .A1(T16270_Y), .A0(T10553_Y));
KC_AOI22_X1 T2963 ( .Y(T2963_Y), .B1(T13396_Q), .B0(T9665_Y),     .A1(T13397_Q), .A0(T15256_Y));
KC_AOI22_X1 T2964 ( .Y(T2964_Y), .B1(T3024_Y), .B0(T13398_Q),     .A1(T15211_Y), .A0(T13412_Q));
KC_AOI22_X1 T2965 ( .Y(T2965_Y), .B1(T14815_Q), .B0(T3611_Y),     .A1(T13395_Q), .A0(T6482_Y));
KC_AOI22_X1 T2967 ( .Y(T2967_Y), .B1(T13428_Q), .B0(T9665_Y),     .A1(T13425_Q), .A0(T15256_Y));
KC_AOI22_X1 T2968 ( .Y(T2968_Y), .B1(T13506_Q), .B0(T9635_Y),     .A1(T13507_Q), .A0(T5088_Y));
KC_AOI22_X1 T2969 ( .Y(T2969_Y), .B1(T13392_Q), .B0(T9635_Y),     .A1(T13393_Q), .A0(T5088_Y));
KC_AOI22_X1 T2970 ( .Y(T2970_Y), .B1(T3024_Y), .B0(T13428_Q),     .A1(T15211_Y), .A0(T13425_Q));
KC_AOI22_X1 T2971 ( .Y(T2971_Y), .B1(T13394_Q), .B0(T9665_Y),     .A1(T13411_Q), .A0(T15256_Y));
KC_AOI22_X1 T2972 ( .Y(T2972_Y), .B1(T13398_Q), .B0(T9665_Y),     .A1(T13412_Q), .A0(T15256_Y));
KC_AOI22_X1 T2974 ( .Y(T2974_Y), .B1(T3027_Y), .B0(T14799_Q),     .A1(T9636_Y), .A0(T14801_Q));
KC_AOI22_X1 T2975 ( .Y(T2975_Y), .B1(T14799_Q), .B0(T3611_Y),     .A1(T14801_Q), .A0(T6482_Y));
KC_AOI22_X1 T2976 ( .Y(T2976_Y), .B1(T14802_Q), .B0(T3611_Y),     .A1(T13527_Q), .A0(T6482_Y));
KC_AOI22_X1 T2977 ( .Y(T2977_Y), .B1(T14782_Q), .B0(T9637_Y),     .A1(T14783_Q), .A0(T6483_Y));
KC_AOI22_X1 T2978 ( .Y(T2978_Y), .B1(T10436_Y), .B0(T14782_Q),     .A1(T10437_Y), .A0(T14783_Q));
KC_AOI22_X1 T2979 ( .Y(T2979_Y), .B1(T3027_Y), .B0(T13509_Q),     .A1(T9636_Y), .A0(T13426_Q));
KC_AOI22_X1 T2982 ( .Y(T2982_Y), .B1(T13526_Q), .B0(T9635_Y),     .A1(T13551_Q), .A0(T5088_Y));
KC_AOI22_X1 T2983 ( .Y(T2983_Y), .B1(T14798_Q), .B0(T9637_Y),     .A1(T13529_Q), .A0(T6483_Y));
KC_AOI22_X1 T2984 ( .Y(T2984_Y), .B1(T10436_Y), .B0(T14798_Q),     .A1(T10437_Y), .A0(T13529_Q));
KC_AOI22_X1 T2986 ( .Y(T2986_Y), .B1(T13554_Q), .B0(T9665_Y),     .A1(T13555_Q), .A0(T15256_Y));
KC_AOI22_X1 T2987 ( .Y(T2987_Y), .B1(T3027_Y), .B0(T14802_Q),     .A1(T9636_Y), .A0(T13527_Q));
KC_AOI22_X1 T2988 ( .Y(T2988_Y), .B1(T9664_Y), .B0(T13526_Q),     .A1(T3610_Y), .A0(T13551_Q));
KC_AOI22_X1 T2989 ( .Y(T2989_Y), .B1(T3024_Y), .B0(T13554_Q),     .A1(T15211_Y), .A0(T13555_Q));
KC_AOI22_X1 T2992 ( .Y(T2992_Y), .B1(T3024_Y), .B0(T13394_Q),     .A1(T15211_Y), .A0(T13411_Q));
KC_AOI22_X1 T2993 ( .Y(T2993_Y), .B1(T13423_Q), .B0(T9635_Y),     .A1(T14814_Q), .A0(T5088_Y));
KC_AOI22_X1 T2994 ( .Y(T2994_Y), .B1(T13509_Q), .B0(T3611_Y),     .A1(T13426_Q), .A0(T6482_Y));
KC_AOI22_X1 T2995 ( .Y(T2995_Y), .B1(T3024_Y), .B0(T13396_Q),     .A1(T15211_Y), .A0(T13397_Q));
KC_AOI22_X1 T2996 ( .Y(T2996_Y), .B1(T6631_Y), .B0(T14761_Q),     .A1(T3001_Y), .A0(T4937_Y));
KC_AOI22_X1 T2997 ( .Y(T2997_Y), .B1(T6635_Y), .B0(T13653_Q),     .A1(T2981_Y), .A0(T4937_Y));
KC_AOI22_X1 T2998 ( .Y(T2998_Y), .B1(T10436_Y), .B0(T13651_Q),     .A1(T10437_Y), .A0(T13637_Q));
KC_AOI22_X1 T2999 ( .Y(T2999_Y), .B1(T6634_Y), .B0(T13639_Q),     .A1(T4937_Y), .A0(T2966_Y));
KC_AOI22_X1 T3002 ( .Y(T3002_Y), .B1(T3024_Y), .B0(T13672_Q),     .A1(T15211_Y), .A0(T13675_Q));
KC_AOI22_X1 T3003 ( .Y(T3003_Y), .B1(T13674_Q), .B0(T9637_Y),     .A1(T13624_Q), .A0(T6483_Y));
KC_AOI22_X1 T3004 ( .Y(T3004_Y), .B1(T3024_Y), .B0(T13676_Q),     .A1(T15211_Y), .A0(T13677_Q));
KC_AOI22_X1 T3005 ( .Y(T3005_Y), .B1(T13676_Q), .B0(T9665_Y),     .A1(T13677_Q), .A0(T15256_Y));
KC_AOI22_X1 T3006 ( .Y(T3006_Y), .B1(T3027_Y), .B0(T14781_Q),     .A1(T9636_Y), .A0(T14780_Q));
KC_AOI22_X1 T3007 ( .Y(T3007_Y), .B1(T10436_Y), .B0(T13674_Q),     .A1(T10437_Y), .A0(T13624_Q));
KC_AOI22_X1 T3015 ( .Y(T3015_Y), .B1(T3586_Y), .B0(T9655_Y),     .A1(T5080_Y), .A0(T3012_Y));
KC_AOI22_X1 T3016 ( .Y(T3016_Y), .B1(T5752_Y), .B0(T14930_Q),     .A1(T4937_Y), .A0(T3586_Y));
KC_AOI22_X1 T3017 ( .Y(T3017_Y), .B1(T3544_Y), .B0(T9669_Y),     .A1(T3020_Y), .A0(T5037_Y));
KC_AOI22_X1 T3018 ( .Y(T3018_Y), .B1(T2966_Y), .B0(T9669_Y),     .A1(T3020_Y), .A0(T5038_Y));
KC_AOI22_X1 T3019 ( .Y(T3019_Y), .B1(T6636_Y), .B0(T13755_Q),     .A1(T4937_Y), .A0(T3544_Y));
KC_AOI22_X1 T3028 ( .Y(T3028_Y), .B1(T9729_Y), .B0(T14045_Q),     .A1(T14049_Q), .A0(T5134_Y));
KC_AOI22_X1 T3029 ( .Y(T3029_Y), .B1(T14044_Q), .B0(T9729_Y),     .A1(T14068_Q), .A0(T5134_Y));
KC_AOI22_X1 T3030 ( .Y(T3030_Y), .B1(T5810_Y), .B0(T14051_Q),     .A1(T5268_Y), .A0(T14994_Y));
KC_AOI22_X1 T3033 ( .Y(T3033_Y), .B1(T9765_Y), .B0(T14837_Q),     .A1(T9768_Y), .A0(T14929_Q));
KC_AOI22_X1 T3034 ( .Y(T3034_Y), .B1(T9765_Y), .B0(T13893_Q),     .A1(T9768_Y), .A0(T14925_Q));
KC_AOI22_X1 T3040 ( .Y(T3040_Y), .B1(T13913_Q), .B0(T9728_Y),     .A1(T13881_Q), .A0(T9767_Y));
KC_AOI22_X1 T3041 ( .Y(T3041_Y), .B1(T13912_Q), .B0(T9728_Y),     .A1(T13910_Q), .A0(T9767_Y));
KC_AOI22_X1 T3042 ( .Y(T3042_Y), .B1(T631_Y), .B0(T14833_Q),     .A1(T3032_Y), .A0(T14830_Q));
KC_AOI22_X1 T3043 ( .Y(T3043_Y), .B1(T9766_Y), .B0(T13911_Q),     .A1(T9764_Y), .A0(T14829_Q));
KC_AOI22_X1 T3044 ( .Y(T3044_Y), .B1(T9765_Y), .B0(T13911_Q),     .A1(T9768_Y), .A0(T14829_Q));
KC_AOI22_X1 T3046 ( .Y(T3046_Y), .B1(T631_Y), .B0(T14831_Q),     .A1(T3032_Y), .A0(T14834_Q));
KC_AOI22_X1 T3047 ( .Y(T3047_Y), .B1(T631_Y), .B0(T14922_Q),     .A1(T3032_Y), .A0(T14926_Q));
KC_AOI22_X1 T3048 ( .Y(T3048_Y), .B1(T13893_Q), .B0(T9766_Y),     .A1(T14925_Q), .A0(T9764_Y));
KC_AOI22_X1 T3049 ( .Y(T3049_Y), .B1(T14835_Q), .B0(T9766_Y),     .A1(T14832_Q), .A0(T9764_Y));
KC_AOI22_X1 T3050 ( .Y(T3050_Y), .B1(T9765_Y), .B0(T14835_Q),     .A1(T9768_Y), .A0(T14832_Q));
KC_AOI22_X1 T3055 ( .Y(T3055_Y), .B1(T9732_Y), .B0(T13929_Q),     .A1(T9730_Y), .A0(T14858_Q));
KC_AOI22_X1 T3056 ( .Y(T3056_Y), .B1(T5811_Y), .B0(T14856_Q),     .A1(T4252_Y), .A0(T14994_Y));
KC_AOI22_X1 T3057 ( .Y(T3057_Y), .B1(T9732_Y), .B0(T13913_Q),     .A1(T9730_Y), .A0(T13881_Q));
KC_AOI22_X1 T3058 ( .Y(T3058_Y), .B1(T9732_Y), .B0(T13879_Q),     .A1(T9730_Y), .A0(T13880_Q));
KC_AOI22_X1 T3059 ( .Y(T3059_Y), .B1(T9728_Y), .B0(T13879_Q),     .A1(T9767_Y), .A0(T13880_Q));
KC_AOI22_X1 T3060 ( .Y(T3060_Y), .B1(T9732_Y), .B0(T13912_Q),     .A1(T9730_Y), .A0(T13910_Q));
KC_AOI22_X1 T3063 ( .Y(T3063_Y), .B1(T3102_Y), .B0(T15218_Y),     .A1(T3036_Y), .A0(T5021_Y));
KC_AOI22_X1 T3064 ( .Y(T3064_Y), .B1(T3087_Y), .B0(T15218_Y),     .A1(T3053_Y), .A0(T5021_Y));
KC_AOI22_X1 T3065 ( .Y(T3065_Y), .B1(T3109_Y), .B0(T15218_Y),     .A1(T3052_Y), .A0(T5021_Y));
KC_AOI22_X1 T3066 ( .Y(T3066_Y), .B1(T9731_Y), .B0(T14045_Q),     .A1(T3640_Y), .A0(T14049_Q));
KC_AOI22_X1 T3067 ( .Y(T3067_Y), .B1(T3094_Y), .B0(T15218_Y),     .A1(T3035_Y), .A0(T5021_Y));
KC_AOI22_X1 T5863 ( .Y(T5863_Y), .B1(T5866_Y), .B0(T14172_Q),     .A1(T14994_Y), .A0(T3146_Y));
KC_AOI22_X1 T3083 ( .Y(T3083_Y), .B1(T10501_Y), .B0(T14197_Q),     .A1(T10502_Y), .A0(T14299_Q));
KC_AOI22_X1 T3084 ( .Y(T3084_Y), .B1(T14298_Q), .B0(T16442_Y),     .A1(T14891_Q), .A0(T15254_Y));
KC_AOI22_X1 T3085 ( .Y(T3085_Y), .B1(T14197_Q), .B0(T9936_Y),     .A1(T14299_Q), .A0(T9937_Y));
KC_AOI22_X1 T3086 ( .Y(T3086_Y), .B1(T14890_Q), .B0(T3117_Y),     .A1(T14300_Q), .A0(T12329_Y));
KC_AOI22_X1 T3088 ( .Y(T3088_Y), .B1(T5579_Y), .B0(T14150_Q),     .A1(T16443_Y), .A0(T14880_Q));
KC_AOI22_X1 T3089 ( .Y(T3089_Y), .B1(T10504_Y), .B0(T14879_Q),     .A1(T15215_Y), .A0(T14092_Q));
KC_AOI22_X1 T3090 ( .Y(T3090_Y), .B1(T10504_Y), .B0(T14090_Q),     .A1(T15215_Y), .A0(T14030_Q));
KC_AOI22_X1 T3091 ( .Y(T3091_Y), .B1(T5579_Y), .B0(T14883_Q),     .A1(T16443_Y), .A0(T14091_Q));
KC_AOI22_X1 T3092 ( .Y(T3092_Y), .B1(T14883_Q), .B0(T3117_Y),     .A1(T14091_Q), .A0(T12329_Y));
KC_AOI22_X1 T3095 ( .Y(T3095_Y), .B1(T5579_Y), .B0(T14194_Q),     .A1(T16443_Y), .A0(T14192_Q));
KC_AOI22_X1 T3096 ( .Y(T3096_Y), .B1(T5579_Y), .B0(T14890_Q),     .A1(T16443_Y), .A0(T14300_Q));
KC_AOI22_X1 T3097 ( .Y(T3097_Y), .B1(T10504_Y), .B0(T14298_Q),     .A1(T15215_Y), .A0(T14891_Q));
KC_AOI22_X1 T3098 ( .Y(T3098_Y), .B1(T3117_Y), .B0(T14194_Q),     .A1(T12329_Y), .A0(T14192_Q));
KC_AOI22_X1 T3099 ( .Y(T3099_Y), .B1(T3108_Y), .B0(T9946_Y),     .A1(T2549_Y), .A0(T5330_Y));
KC_AOI22_X1 T3100 ( .Y(T3100_Y), .B1(T10501_Y), .B0(T14183_Q),     .A1(T10502_Y), .A0(T14181_Q));
KC_AOI22_X1 T3101 ( .Y(T3101_Y), .B1(T14183_Q), .B0(T9936_Y),     .A1(T14181_Q), .A0(T9937_Y));
KC_AOI22_X1 T3104 ( .Y(T3104_Y), .B1(T16442_Y), .B0(T14193_Q),     .A1(T15254_Y), .A0(T14167_Q));
KC_AOI22_X1 T3105 ( .Y(T3105_Y), .B1(T10504_Y), .B0(T14193_Q),     .A1(T15215_Y), .A0(T14167_Q));
KC_AOI22_X1 T3106 ( .Y(T3106_Y), .B1(T9936_Y), .B0(T14169_Q),     .A1(T9937_Y), .A0(T14168_Q));
KC_AOI22_X1 T3107 ( .Y(T3107_Y), .B1(T10501_Y), .B0(T14169_Q),     .A1(T10502_Y), .A0(T14168_Q));
KC_AOI22_X1 T3111 ( .Y(T3111_Y), .B1(T14147_Q), .B0(T9936_Y),     .A1(T14148_Q), .A0(T9937_Y));
KC_AOI22_X1 T3112 ( .Y(T3112_Y), .B1(T14879_Q), .B0(T16442_Y),     .A1(T14092_Q), .A0(T15254_Y));
KC_AOI22_X1 T3113 ( .Y(T3113_Y), .B1(T14090_Q), .B0(T16442_Y),     .A1(T14030_Q), .A0(T15254_Y));
KC_AOI22_X1 T3114 ( .Y(T3114_Y), .B1(T10501_Y), .B0(T14147_Q),     .A1(T10502_Y), .A0(T14148_Q));
KC_AOI22_X1 T3115 ( .Y(T3115_Y), .B1(T14150_Q), .B0(T3117_Y),     .A1(T14880_Q), .A0(T12329_Y));
KC_AOI22_X1 T3124 ( .Y(T3124_Y), .B1(T14364_Q), .B0(T3117_Y),     .A1(T14359_Q), .A0(T12329_Y));
KC_AOI22_X1 T3125 ( .Y(T3125_Y), .B1(T14365_Q), .B0(T9936_Y),     .A1(T14362_Q), .A0(T9937_Y));
KC_AOI22_X1 T3126 ( .Y(T3126_Y), .B1(T14338_Q), .B0(T9936_Y),     .A1(T14357_Q), .A0(T9937_Y));
KC_AOI22_X1 T3127 ( .Y(T3127_Y), .B1(T10501_Y), .B0(T14338_Q),     .A1(T10502_Y), .A0(T14357_Q));
KC_AOI22_X1 T3128 ( .Y(T3128_Y), .B1(T10501_Y), .B0(T14365_Q),     .A1(T10502_Y), .A0(T14362_Q));
KC_AOI22_X1 T3131 ( .Y(T3131_Y), .B1(T10501_Y), .B0(T14343_Q),     .A1(T10502_Y), .A0(T14341_Q));
KC_AOI22_X1 T3132 ( .Y(T3132_Y), .B1(T14343_Q), .B0(T9936_Y),     .A1(T14341_Q), .A0(T9937_Y));
KC_AOI22_X1 T3133 ( .Y(T3133_Y), .B1(T5579_Y), .B0(T14344_Q),     .A1(T16443_Y), .A0(T14339_Q));
KC_AOI22_X1 T3134 ( .Y(T3134_Y), .B1(T10504_Y), .B0(T14360_Q),     .A1(T15215_Y), .A0(T14340_Q));
KC_AOI22_X1 T3135 ( .Y(T3135_Y), .B1(T14360_Q), .B0(T16442_Y),     .A1(T14340_Q), .A0(T15254_Y));
KC_AOI22_X1 T3136 ( .Y(T3136_Y), .B1(T14344_Q), .B0(T3117_Y),     .A1(T14339_Q), .A0(T12329_Y));
KC_AOI22_X1 T3139 ( .Y(T3139_Y), .B1(T14323_Q), .B0(T16442_Y),     .A1(T14325_Q), .A0(T15254_Y));
KC_AOI22_X1 T3140 ( .Y(T3140_Y), .B1(T10504_Y), .B0(T14323_Q),     .A1(T15215_Y), .A0(T14325_Q));
KC_AOI22_X1 T3141 ( .Y(T3141_Y), .B1(T5579_Y), .B0(T14318_Q),     .A1(T16443_Y), .A0(T14315_Q));
KC_AOI22_X1 T3142 ( .Y(T3142_Y), .B1(T14318_Q), .B0(T3117_Y),     .A1(T14315_Q), .A0(T12329_Y));
KC_AOI22_X1 T3143 ( .Y(T3143_Y), .B1(T10501_Y), .B0(T14316_Q),     .A1(T10502_Y), .A0(T14296_Q));
KC_AOI22_X1 T3144 ( .Y(T3144_Y), .B1(T14316_Q), .B0(T9936_Y),     .A1(T14296_Q), .A0(T9937_Y));
KC_AOI22_X1 T3162 ( .Y(T3162_Y), .B1(T5579_Y), .B0(T14450_Q),     .A1(T16443_Y), .A0(T14446_Q));
KC_AOI22_X1 T3163 ( .Y(T3163_Y), .B1(T14909_Q), .B0(T16442_Y),     .A1(T14908_Q), .A0(T15254_Y));
KC_AOI22_X1 T3164 ( .Y(T3164_Y), .B1(T14450_Q), .B0(T3117_Y),     .A1(T14446_Q), .A0(T12329_Y));
KC_AOI22_X1 T3165 ( .Y(T3165_Y), .B1(T14447_Q), .B0(T16442_Y),     .A1(T14444_Q), .A0(T15254_Y));
KC_AOI22_X1 T3168 ( .Y(T3168_Y), .B1(T14423_Q), .B0(T3117_Y),     .A1(T14433_Q), .A0(T12329_Y));
KC_AOI22_X1 T3169 ( .Y(T3169_Y), .B1(T10501_Y), .B0(T14449_Q),     .A1(T10502_Y), .A0(T14907_Q));
KC_AOI22_X1 T3170 ( .Y(T3170_Y), .B1(T14449_Q), .B0(T9936_Y),     .A1(T14907_Q), .A0(T9937_Y));
KC_AOI22_X1 T3172 ( .Y(T3172_Y), .B1(T14432_Q), .B0(T16442_Y),     .A1(T14419_Q), .A0(T15254_Y));
KC_AOI22_X1 T3173 ( .Y(T3173_Y), .B1(T5579_Y), .B0(T14423_Q),     .A1(T16443_Y), .A0(T14433_Q));
KC_AOI22_X1 T3174 ( .Y(T3174_Y), .B1(T10501_Y), .B0(T14424_Q),     .A1(T10502_Y), .A0(T14420_Q));
KC_AOI22_X1 T3175 ( .Y(T3175_Y), .B1(T14424_Q), .B0(T9936_Y),     .A1(T14420_Q), .A0(T9937_Y));
KC_AOI22_X1 T3178 ( .Y(T3178_Y), .B1(T14402_Q), .B0(T9936_Y),     .A1(T14400_Q), .A0(T9937_Y));
KC_AOI22_X1 T3179 ( .Y(T3179_Y), .B1(T10504_Y), .B0(T14399_Q),     .A1(T15215_Y), .A0(T14421_Q));
KC_AOI22_X1 T3180 ( .Y(T3180_Y), .B1(T14399_Q), .B0(T16442_Y),     .A1(T14421_Q), .A0(T15254_Y));
KC_AOI22_X1 T3181 ( .Y(T3181_Y), .B1(T5579_Y), .B0(T14401_Q),     .A1(T16443_Y), .A0(T14396_Q));
KC_AOI22_X1 T3182 ( .Y(T3182_Y), .B1(T10501_Y), .B0(T14402_Q),     .A1(T10502_Y), .A0(T14400_Q));
KC_AOI22_X1 T3183 ( .Y(T3183_Y), .B1(T14401_Q), .B0(T3117_Y),     .A1(T14396_Q), .A0(T12329_Y));
KC_AOI22_X1 T3247 ( .Y(T3247_Y), .B1(T3226_Q), .B0(T5141_Y),     .A1(T3878_Q), .A0(T11506_Y));
KC_AOI22_X1 T3291 ( .Y(T3291_Y), .B1(T3314_Y), .B0(T3292_Y),     .A1(T12202_Y), .A0(T11485_Y));
KC_AOI22_X1 T3356 ( .Y(T3356_Y), .B1(T16037_Y), .B0(T2806_Y),     .A1(T8278_Y), .A0(T12263_Y));
KC_AOI22_X1 T3357 ( .Y(T3357_Y), .B1(T15598_Y), .B0(T964_Q),     .A1(T8259_Y), .A0(T12263_Y));
KC_AOI22_X1 T3392 ( .Y(T3392_Y), .B1(T3378_Y), .B0(T12876_Y),     .A1(T10968_Y), .A0(T11769_Y));
KC_AOI22_X1 T3422 ( .Y(T3422_Y), .B1(T3416_Y), .B0(T3412_Q),     .A1(T13177_Y), .A0(T6549_Q));
KC_AOI22_X1 T3423 ( .Y(T3423_Y), .B1(T3421_Y), .B0(T6141_Y),     .A1(T11719_Y), .A0(T8510_Y));
KC_AOI22_X1 T3434 ( .Y(T3434_Y), .B1(T6579_Y), .B0(T12104_Y),     .A1(T11702_Y), .A0(T6139_Y));
KC_AOI22_X1 T6584 ( .Y(T6584_Y), .B1(T11805_Y), .B0(T6561_Y),     .A1(T15761_Y), .A0(T6586_Y));
KC_AOI22_X1 T3463 ( .Y(T3463_Y), .B1(T15234_Y), .B0(T15616_Y),     .A1(T5109_Y), .A0(T11816_Y));
KC_AOI22_X1 T3464 ( .Y(T3464_Y), .B1(T12874_Y), .B0(T6561_Y),     .A1(T8503_Y), .A0(T5116_Y));
KC_AOI22_X1 T3471 ( .Y(T3471_Y), .B1(T3475_Y), .B0(T6209_Y),     .A1(T10995_Y), .A0(T16082_Q));
KC_AOI22_X1 T3472 ( .Y(T3472_Y), .B1(T11721_Y), .B0(T6586_Y),     .A1(T3446_Y), .A0(T8503_Y));
KC_AOI22_X1 T3476 ( .Y(T3476_Y), .B1(T10991_Y), .B0(T6568_S),     .A1(T2923_Y), .A0(T6238_Y));
KC_AOI22_X1 T3488 ( .Y(T3488_Y), .B1(T6211_Y), .B0(T4609_Y),     .A1(T2926_Y), .A0(T11742_Y));
KC_AOI22_X1 T3491 ( .Y(T3491_Y), .B1(T6611_S), .B0(T10571_Y),     .A1(T12107_Y), .A0(T10553_Y));
KC_AOI22_X1 T3492 ( .Y(T3492_Y), .B1(T10987_Y), .B0(T11742_Y),     .A1(T6591_S), .A0(T10571_Y));
KC_AOI22_X1 T3493 ( .Y(T3493_Y), .B1(T10987_Y), .B0(T6196_Y),     .A1(T4128_Y), .A0(T8503_Y));
KC_AOI22_X1 T3518 ( .Y(T3518_Y), .B1(T8425_Y), .B0(T11817_Y),     .A1(T10593_Y), .A0(T6610_S));
KC_AOI22_X1 T3537 ( .Y(T3537_Y), .B1(T13388_Q), .B0(T9665_Y),     .A1(T13420_Q), .A0(T15256_Y));
KC_AOI22_X1 T3538 ( .Y(T3538_Y), .B1(T3024_Y), .B0(T13388_Q),     .A1(T15211_Y), .A0(T13420_Q));
KC_AOI22_X1 T3539 ( .Y(T3539_Y), .B1(T13418_Q), .B0(T9635_Y),     .A1(T13417_Q), .A0(T5088_Y));
KC_AOI22_X1 T3540 ( .Y(T3540_Y), .B1(T13403_Q), .B0(T9665_Y),     .A1(T13404_Q), .A0(T15256_Y));
KC_AOI22_X1 T3541 ( .Y(T3541_Y), .B1(T3024_Y), .B0(T13403_Q),     .A1(T15211_Y), .A0(T13404_Q));
KC_AOI22_X1 T3542 ( .Y(T3542_Y), .B1(T9664_Y), .B0(T13405_Q),     .A1(T3610_Y), .A0(T13406_Q));
KC_AOI22_X1 T3543 ( .Y(T3543_Y), .B1(T13405_Q), .B0(T9635_Y),     .A1(T13406_Q), .A0(T5088_Y));
KC_AOI22_X1 T3546 ( .Y(T3546_Y), .B1(T14776_Q), .B0(T9637_Y),     .A1(T13520_Q), .A0(T6483_Y));
KC_AOI22_X1 T3547 ( .Y(T3547_Y), .B1(T10436_Y), .B0(T14776_Q),     .A1(T10437_Y), .A0(T13520_Q));
KC_AOI22_X1 T3550 ( .Y(T3550_Y), .B1(T13550_Q), .B0(T9637_Y),     .A1(T13548_Q), .A0(T6483_Y));
KC_AOI22_X1 T3551 ( .Y(T3551_Y), .B1(T13546_Q), .B0(T3611_Y),     .A1(T13549_Q), .A0(T6482_Y));
KC_AOI22_X1 T3552 ( .Y(T3552_Y), .B1(T3027_Y), .B0(T13546_Q),     .A1(T9636_Y), .A0(T13549_Q));
KC_AOI22_X1 T3553 ( .Y(T3553_Y), .B1(T10436_Y), .B0(T13550_Q),     .A1(T10437_Y), .A0(T13548_Q));
KC_AOI22_X1 T3554 ( .Y(T3554_Y), .B1(T13540_Q), .B0(T9637_Y),     .A1(T13547_Q), .A0(T6483_Y));
KC_AOI22_X1 T3555 ( .Y(T3555_Y), .B1(T10436_Y), .B0(T13540_Q),     .A1(T10437_Y), .A0(T13547_Q));
KC_AOI22_X1 T3556 ( .Y(T3556_Y), .B1(T3027_Y), .B0(T13521_Q),     .A1(T9636_Y), .A0(T14777_Q));
KC_AOI22_X1 T3557 ( .Y(T3557_Y), .B1(T13522_Q), .B0(T9635_Y),     .A1(T14795_Q), .A0(T5088_Y));
KC_AOI22_X1 T3558 ( .Y(T3558_Y), .B1(T13541_Q), .B0(T9637_Y),     .A1(T13523_Q), .A0(T6483_Y));
KC_AOI22_X1 T3559 ( .Y(T3559_Y), .B1(T13539_Q), .B0(T9635_Y),     .A1(T13545_Q), .A0(T5088_Y));
KC_AOI22_X1 T3560 ( .Y(T3560_Y), .B1(T9664_Y), .B0(T13539_Q),     .A1(T3610_Y), .A0(T13545_Q));
KC_AOI22_X1 T3561 ( .Y(T3561_Y), .B1(T10436_Y), .B0(T13541_Q),     .A1(T10437_Y), .A0(T13523_Q));
KC_AOI22_X1 T3562 ( .Y(T3562_Y), .B1(T9664_Y), .B0(T13522_Q),     .A1(T3610_Y), .A0(T14795_Q));
KC_AOI22_X1 T3563 ( .Y(T3563_Y), .B1(T13521_Q), .B0(T3611_Y),     .A1(T14777_Q), .A0(T6482_Y));
KC_AOI22_X1 T3567 ( .Y(T3567_Y), .B1(T3027_Y), .B0(T13422_Q),     .A1(T9636_Y), .A0(T13419_Q));
KC_AOI22_X1 T3568 ( .Y(T3568_Y), .B1(T13505_Q), .B0(T9665_Y),     .A1(T13504_Q), .A0(T15256_Y));
KC_AOI22_X1 T3569 ( .Y(T3569_Y), .B1(T3024_Y), .B0(T13505_Q),     .A1(T15211_Y), .A0(T13504_Q));
KC_AOI22_X1 T3570 ( .Y(T3570_Y), .B1(T3027_Y), .B0(T13390_Q),     .A1(T9636_Y), .A0(T14813_Q));
KC_AOI22_X1 T3571 ( .Y(T3571_Y), .B1(T13422_Q), .B0(T3611_Y),     .A1(T13419_Q), .A0(T6482_Y));
KC_AOI22_X1 T3572 ( .Y(T3572_Y), .B1(T13390_Q), .B0(T3611_Y),     .A1(T14813_Q), .A0(T6482_Y));
KC_AOI22_X1 T5733 ( .Y(T5733_Y), .B1(T13652_Q), .B0(T9637_Y),     .A1(T13638_Q), .A0(T6483_Y));
KC_AOI22_X1 T3573 ( .Y(T3573_Y), .B1(T10436_Y), .B0(T13670_Q),     .A1(T10437_Y), .A0(T13635_Q));
KC_AOI22_X1 T3574 ( .Y(T3574_Y), .B1(T10436_Y), .B0(T13673_Q),     .A1(T10437_Y), .A0(T13636_Q));
KC_AOI22_X1 T3575 ( .Y(T3575_Y), .B1(T9637_Y), .B0(T13673_Q),     .A1(T6483_Y), .A0(T13636_Q));
KC_AOI22_X1 T3576 ( .Y(T3576_Y), .B1(T10436_Y), .B0(T13652_Q),     .A1(T10437_Y), .A0(T13638_Q));
KC_AOI22_X1 T3577 ( .Y(T3577_Y), .B1(T13670_Q), .B0(T9637_Y),     .A1(T13635_Q), .A0(T6483_Y));
KC_AOI22_X1 T3580 ( .Y(T3580_Y), .B1(T13669_Q), .B0(T9637_Y),     .A1(T13623_Q), .A0(T6483_Y));
KC_AOI22_X1 T3581 ( .Y(T3581_Y), .B1(T3024_Y), .B0(T13668_Q),     .A1(T15211_Y), .A0(T13671_Q));
KC_AOI22_X1 T3582 ( .Y(T3582_Y), .B1(T13668_Q), .B0(T9665_Y),     .A1(T13671_Q), .A0(T15256_Y));
KC_AOI22_X1 T3583 ( .Y(T3583_Y), .B1(T10436_Y), .B0(T13669_Q),     .A1(T10437_Y), .A0(T13623_Q));
KC_AOI22_X1 T3590 ( .Y(T3590_Y), .B1(T3024_Y), .B0(T13768_Q),     .A1(T15211_Y), .A0(T13754_Q));
KC_AOI22_X1 T3591 ( .Y(T3591_Y), .B1(T13764_Q), .B0(T9635_Y),     .A1(T13747_Q), .A0(T5088_Y));
KC_AOI22_X1 T3592 ( .Y(T3592_Y), .B1(T13750_Q), .B0(T9635_Y),     .A1(T13759_Q), .A0(T5088_Y));
KC_AOI22_X1 T3593 ( .Y(T3593_Y), .B1(T9664_Y), .B0(T13764_Q),     .A1(T3610_Y), .A0(T13747_Q));
KC_AOI22_X1 T3594 ( .Y(T3594_Y), .B1(T9635_Y), .B0(T13647_Q),     .A1(T13763_Q), .A0(T5088_Y));
KC_AOI22_X1 T3595 ( .Y(T3595_Y), .B1(T9665_Y), .B0(T13768_Q),     .A1(T15256_Y), .A0(T13754_Q));
KC_AOI22_X1 T3596 ( .Y(T3596_Y), .B1(T3024_Y), .B0(T13766_Q),     .A1(T15211_Y), .A0(T13751_Q));
KC_AOI22_X1 T3597 ( .Y(T3597_Y), .B1(T13756_Q), .B0(T9665_Y),     .A1(T13765_Q), .A0(T15256_Y));
KC_AOI22_X1 T3598 ( .Y(T3598_Y), .B1(T13766_Q), .B0(T9665_Y),     .A1(T13751_Q), .A0(T15256_Y));
KC_AOI22_X1 T3599 ( .Y(T3599_Y), .B1(T9664_Y), .B0(T13750_Q),     .A1(T3610_Y), .A0(T13759_Q));
KC_AOI22_X1 T3600 ( .Y(T3600_Y), .B1(T3024_Y), .B0(T14927_Q),     .A1(T15211_Y), .A0(T14918_Q));
KC_AOI22_X1 T3601 ( .Y(T3601_Y), .B1(T14927_Q), .B0(T9665_Y),     .A1(T14918_Q), .A0(T15256_Y));
KC_AOI22_X1 T3602 ( .Y(T3602_Y), .B1(T3024_Y), .B0(T13756_Q),     .A1(T15211_Y), .A0(T13765_Q));
KC_AOI22_X1 T3606 ( .Y(T3606_Y), .B1(T14762_Q), .B0(T3611_Y),     .A1(T14764_Q), .A0(T6482_Y));
KC_AOI22_X1 T3609 ( .Y(T3609_Y), .B1(T14826_Q), .B0(T9866_Y),     .A1(T14920_Q), .A0(T15222_Y));
KC_AOI22_X1 T6847 ( .Y(T6847_Y), .B1(T13909_Q), .B0(T9863_Y),     .A1(T13904_Q), .A0(T9868_Y));
KC_AOI22_X1 T3612 ( .Y(T3612_Y), .B1(T14048_Q), .B0(T9729_Y),     .A1(T14853_Q), .A0(T5134_Y));
KC_AOI22_X1 T3613 ( .Y(T3613_Y), .B1(T14852_Q), .B0(T9866_Y),     .A1(T14850_Q), .A0(T15222_Y));
KC_AOI22_X1 T3615 ( .Y(T3615_Y), .B1(T12084_Y), .B0(T14915_Q),     .A1(T15219_Y), .A0(T14919_Q));
KC_AOI22_X1 T3616 ( .Y(T3616_Y), .B1(T14828_Q), .B0(T9866_Y),     .A1(T14916_Q), .A0(T15222_Y));
KC_AOI22_X1 T3618 ( .Y(T3618_Y), .B1(T9862_Y), .B0(T13925_Q),     .A1(T9824_Y), .A0(T13876_Q));
KC_AOI22_X1 T3619 ( .Y(T3619_Y), .B1(T13925_Q), .B0(T9863_Y),     .A1(T13876_Q), .A0(T9868_Y));
KC_AOI22_X1 T3620 ( .Y(T3620_Y), .B1(T12084_Y), .B0(T14852_Q),     .A1(T15219_Y), .A0(T14850_Q));
KC_AOI22_X1 T3624 ( .Y(T3624_Y), .B1(T9862_Y), .B0(T13903_Q),     .A1(T9824_Y), .A0(T13908_Q));
KC_AOI22_X1 T3625 ( .Y(T3625_Y), .B1(T13903_Q), .B0(T9863_Y),     .A1(T13908_Q), .A0(T9868_Y));
KC_AOI22_X1 T3629 ( .Y(T3629_Y), .B1(T14831_Q), .B0(T9763_Y),     .A1(T14834_Q), .A0(T3623_Y));
KC_AOI22_X1 T3630 ( .Y(T3630_Y), .B1(T631_Y), .B0(T14923_Q),     .A1(T3032_Y), .A0(T14924_Q));
KC_AOI22_X1 T3631 ( .Y(T3631_Y), .B1(T9862_Y), .B0(T14827_Q),     .A1(T9824_Y), .A0(T13892_Q));
KC_AOI22_X1 T3632 ( .Y(T3632_Y), .B1(T9823_Y), .B0(T14917_Q),     .A1(T9825_Y), .A0(T14910_Q));
KC_AOI22_X1 T3633 ( .Y(T3633_Y), .B1(T14915_Q), .B0(T9866_Y),     .A1(T14919_Q), .A0(T15222_Y));
KC_AOI22_X1 T3634 ( .Y(T3634_Y), .B1(T14827_Q), .B0(T9863_Y),     .A1(T13892_Q), .A0(T9868_Y));
KC_AOI22_X1 T3637 ( .Y(T3637_Y), .B1(T9862_Y), .B0(T13909_Q),     .A1(T9824_Y), .A0(T13904_Q));
KC_AOI22_X1 T3652 ( .Y(T3652_Y), .B1(T14029_Q), .B0(T9863_Y),     .A1(T14875_Q), .A0(T9868_Y));
KC_AOI22_X1 T3658 ( .Y(T3658_Y), .B1(T12084_Y), .B0(T14064_Q),     .A1(T15219_Y), .A0(T14041_Q));
KC_AOI22_X1 T3659 ( .Y(T3659_Y), .B1(T14065_Q), .B0(T9863_Y),     .A1(T14066_Q), .A0(T9868_Y));
KC_AOI22_X1 T3660 ( .Y(T3660_Y), .B1(T9862_Y), .B0(T14065_Q),     .A1(T9824_Y), .A0(T14066_Q));
KC_AOI22_X1 T3661 ( .Y(T3661_Y), .B1(T9823_Y), .B0(T14043_Q),     .A1(T9825_Y), .A0(T14042_Q));
KC_AOI22_X1 T3662 ( .Y(T3662_Y), .B1(T14064_Q), .B0(T9866_Y),     .A1(T14041_Q), .A0(T15222_Y));
KC_AOI22_X1 T3663 ( .Y(T3663_Y), .B1(T3708_Y), .B0(T16165_Y),     .A1(T3604_Y), .A0(T2532_Y));
KC_AOI22_X1 T3664 ( .Y(T3664_Y), .B1(T4306_Y), .B0(T16165_Y),     .A1(T3603_Y), .A0(T2532_Y));
KC_AOI22_X1 T3665 ( .Y(T3665_Y), .B1(T3709_Y), .B0(T16165_Y),     .A1(T3588_Y), .A0(T2532_Y));
KC_AOI22_X1 T3671 ( .Y(T3671_Y), .B1(T9862_Y), .B0(T14029_Q),     .A1(T9824_Y), .A0(T14875_Q));
KC_AOI22_X1 T3672 ( .Y(T3672_Y), .B1(T14876_Q), .B0(T9866_Y),     .A1(T14088_Q), .A0(T15222_Y));
KC_AOI22_X1 T3673 ( .Y(T3673_Y), .B1(T12084_Y), .B0(T14876_Q),     .A1(T15219_Y), .A0(T14088_Q));
KC_AOI22_X1 T3674 ( .Y(T3674_Y), .B1(T14087_Q), .B0(T9864_Y),     .A1(T14089_Q), .A0(T9865_Y));
KC_AOI22_X1 T3675 ( .Y(T3675_Y), .B1(T9823_Y), .B0(T14087_Q),     .A1(T9825_Y), .A0(T14089_Q));
KC_AOI22_X1 T6689 ( .Y(T6689_Y), .B1(T12084_Y), .B0(T14295_Q),     .A1(T15219_Y), .A0(T14289_Q));
KC_AOI22_X1 T6688 ( .Y(T6688_Y), .B1(T14888_Q), .B0(T9863_Y),     .A1(T14189_Q), .A0(T9868_Y));
KC_AOI22_X1 T3686 ( .Y(T3686_Y), .B1(T14293_Q), .B0(T9866_Y),     .A1(T14312_Q), .A0(T15222_Y));
KC_AOI22_X1 T3687 ( .Y(T3687_Y), .B1(T14291_Q), .B0(T9863_Y),     .A1(T14309_Q), .A0(T9868_Y));
KC_AOI22_X1 T3689 ( .Y(T3689_Y), .B1(T9862_Y), .B0(T14878_Q),     .A1(T9824_Y), .A0(T14874_Q));
KC_AOI22_X1 T3690 ( .Y(T3690_Y), .B1(T14878_Q), .B0(T9863_Y),     .A1(T14874_Q), .A0(T9868_Y));
KC_AOI22_X1 T3691 ( .Y(T3691_Y), .B1(T12084_Y), .B0(T14146_Q),     .A1(T15219_Y), .A0(T14140_Q));
KC_AOI22_X1 T3693 ( .Y(T3693_Y), .B1(T9866_Y), .B0(T14295_Q),     .A1(T15222_Y), .A0(T14289_Q));
KC_AOI22_X1 T3694 ( .Y(T3694_Y), .B1(T10503_Y), .B0(T14302_Q),     .A1(T3684_Y), .A0(T14889_Q));
KC_AOI22_X1 T3695 ( .Y(T3695_Y), .B1(T9862_Y), .B0(T14291_Q),     .A1(T9824_Y), .A0(T14309_Q));
KC_AOI22_X1 T3696 ( .Y(T3696_Y), .B1(T9862_Y), .B0(T14888_Q),     .A1(T9824_Y), .A0(T14189_Q));
KC_AOI22_X1 T3697 ( .Y(T3697_Y), .B1(T9863_Y), .B0(T14190_Q),     .A1(T9868_Y), .A0(T14191_Q));
KC_AOI22_X1 T3698 ( .Y(T3698_Y), .B1(T9932_Y), .B0(T14196_Q),     .A1(T14160_Q), .A0(T3719_Y));
KC_AOI22_X1 T3699 ( .Y(T3699_Y), .B1(T10503_Y), .B0(T14196_Q),     .A1(T3684_Y), .A0(T14160_Q));
KC_AOI22_X1 T3700 ( .Y(T3700_Y), .B1(T12084_Y), .B0(T14293_Q),     .A1(T15219_Y), .A0(T14312_Q));
KC_AOI22_X1 T3701 ( .Y(T3701_Y), .B1(T14163_Q), .B0(T9864_Y),     .A1(T14162_Q), .A0(T9865_Y));
KC_AOI22_X1 T3702 ( .Y(T3702_Y), .B1(T14161_Q), .B0(T9864_Y),     .A1(T14165_Q), .A0(T9865_Y));
KC_AOI22_X1 T3703 ( .Y(T3703_Y), .B1(T10503_Y), .B0(T14171_Q),     .A1(T3684_Y), .A0(T14166_Q));
KC_AOI22_X1 T3704 ( .Y(T3704_Y), .B1(T14171_Q), .B0(T9932_Y),     .A1(T14166_Q), .A0(T3719_Y));
KC_AOI22_X1 T3705 ( .Y(T3705_Y), .B1(T9823_Y), .B0(T14143_Q),     .A1(T9825_Y), .A0(T14180_Q));
KC_AOI22_X1 T3706 ( .Y(T3706_Y), .B1(T9864_Y), .B0(T14143_Q),     .A1(T9865_Y), .A0(T14180_Q));
KC_AOI22_X1 T3710 ( .Y(T3710_Y), .B1(T9862_Y), .B0(T14190_Q),     .A1(T9824_Y), .A0(T14191_Q));
KC_AOI22_X1 T3711 ( .Y(T3711_Y), .B1(T9823_Y), .B0(T14161_Q),     .A1(T9825_Y), .A0(T14165_Q));
KC_AOI22_X1 T3714 ( .Y(T3714_Y), .B1(T14145_Q), .B0(T9864_Y),     .A1(T14144_Q), .A0(T9865_Y));
KC_AOI22_X1 T3715 ( .Y(T3715_Y), .B1(T10503_Y), .B0(T14149_Q),     .A1(T3684_Y), .A0(T14142_Q));
KC_AOI22_X1 T3716 ( .Y(T3716_Y), .B1(T9823_Y), .B0(T14145_Q),     .A1(T9825_Y), .A0(T14144_Q));
KC_AOI22_X1 T3717 ( .Y(T3717_Y), .B1(T14146_Q), .B0(T9866_Y),     .A1(T14140_Q), .A0(T15222_Y));
KC_AOI22_X1 T3718 ( .Y(T3718_Y), .B1(T14149_Q), .B0(T9932_Y),     .A1(T14142_Q), .A0(T3719_Y));
KC_AOI22_X1 T3721 ( .Y(T3721_Y), .B1(T14361_Q), .B0(T3117_Y),     .A1(T14358_Q), .A0(T12329_Y));
KC_AOI22_X1 T3722 ( .Y(T3722_Y), .B1(T14334_Q), .B0(T9932_Y),     .A1(T14336_Q), .A0(T3719_Y));
KC_AOI22_X1 T3723 ( .Y(T3723_Y), .B1(T10503_Y), .B0(T14334_Q),     .A1(T3684_Y), .A0(T14336_Q));
KC_AOI22_X1 T3724 ( .Y(T3724_Y), .B1(T10504_Y), .B0(T14337_Q),     .A1(T15215_Y), .A0(T14335_Q));
KC_AOI22_X1 T3725 ( .Y(T3725_Y), .B1(T14337_Q), .B0(T16442_Y),     .A1(T14335_Q), .A0(T15254_Y));
KC_AOI22_X1 T3726 ( .Y(T3726_Y), .B1(T10503_Y), .B0(T14322_Q),     .A1(T3684_Y), .A0(T14308_Q));
KC_AOI22_X1 T3727 ( .Y(T3727_Y), .B1(T14322_Q), .B0(T9932_Y),     .A1(T14308_Q), .A0(T3719_Y));
KC_AOI22_X1 T3729 ( .Y(T3729_Y), .B1(T10503_Y), .B0(T14307_Q),     .A1(T3684_Y), .A0(T14310_Q));
KC_AOI22_X1 T3730 ( .Y(T3730_Y), .B1(T14307_Q), .B0(T9932_Y),     .A1(T14310_Q), .A0(T3719_Y));
KC_AOI22_X1 T3731 ( .Y(T3731_Y), .B1(T10504_Y), .B0(T14317_Q),     .A1(T15215_Y), .A0(T14313_Q));
KC_AOI22_X1 T3732 ( .Y(T3732_Y), .B1(T10503_Y), .B0(T14288_Q),     .A1(T3684_Y), .A0(T14292_Q));
KC_AOI22_X1 T3733 ( .Y(T3733_Y), .B1(T14302_Q), .B0(T9932_Y),     .A1(T14889_Q), .A0(T3719_Y));
KC_AOI22_X1 T3734 ( .Y(T3734_Y), .B1(T14288_Q), .B0(T9932_Y),     .A1(T14292_Q), .A0(T3719_Y));
KC_AOI22_X1 T5977 ( .Y(T5977_Y), .B1(T10501_Y), .B0(T14900_Q),     .A1(T10502_Y), .A0(T14505_Q));
KC_AOI22_X1 T5976 ( .Y(T5976_Y), .B1(T10501_Y), .B0(T14442_Q),     .A1(T10502_Y), .A0(T14439_Q));
KC_AOI22_X1 T3736 ( .Y(T3736_Y), .B1(T5579_Y), .B0(T14506_Q),     .A1(T16443_Y), .A0(T14902_Q));
KC_AOI22_X1 T3737 ( .Y(T3737_Y), .B1(T5579_Y), .B0(T14903_Q),     .A1(T16443_Y), .A0(T14904_Q));
KC_AOI22_X1 T3743 ( .Y(T3743_Y), .B1(T14900_Q), .B0(T9936_Y),     .A1(T14505_Q), .A0(T9937_Y));
KC_AOI22_X1 T3744 ( .Y(T3744_Y), .B1(T14905_Q), .B0(T3117_Y),     .A1(T14906_Q), .A0(T12329_Y));
KC_AOI22_X1 T3745 ( .Y(T3745_Y), .B1(T14903_Q), .B0(T3117_Y),     .A1(T14904_Q), .A0(T12329_Y));
KC_AOI22_X1 T3746 ( .Y(T3746_Y), .B1(T14506_Q), .B0(T3117_Y),     .A1(T14902_Q), .A0(T12329_Y));
KC_AOI22_X1 T3747 ( .Y(T3747_Y), .B1(T5579_Y), .B0(T14905_Q),     .A1(T16443_Y), .A0(T14906_Q));
KC_AOI22_X1 T3748 ( .Y(T3748_Y), .B1(T14442_Q), .B0(T9936_Y),     .A1(T14439_Q), .A0(T9937_Y));
KC_AOI22_X1 T3749 ( .Y(T3749_Y), .B1(T14441_Q), .B0(T16442_Y),     .A1(T14440_Q), .A0(T15254_Y));
KC_AOI22_X1 T3751 ( .Y(T3751_Y), .B1(T14448_Q), .B0(T9936_Y),     .A1(T14445_Q), .A0(T9937_Y));
KC_AOI22_X1 T3752 ( .Y(T3752_Y), .B1(T14443_Q), .B0(T16442_Y),     .A1(T14438_Q), .A0(T15254_Y));
KC_AOI22_X1 T3753 ( .Y(T3753_Y), .B1(T10501_Y), .B0(T14448_Q),     .A1(T10502_Y), .A0(T14445_Q));
KC_AOI22_X1 T3754 ( .Y(T3754_Y), .B1(T10504_Y), .B0(T14441_Q),     .A1(T15215_Y), .A0(T14440_Q));
KC_AOI22_X1 T3755 ( .Y(T3755_Y), .B1(T10504_Y), .B0(T14443_Q),     .A1(T15215_Y), .A0(T14438_Q));
KC_AOI22_X1 T3756 ( .Y(T3756_Y), .B1(T10504_Y), .B0(T14422_Q),     .A1(T15215_Y), .A0(T14431_Q));
KC_AOI22_X1 T3757 ( .Y(T3757_Y), .B1(T14414_Q), .B0(T16442_Y),     .A1(T14416_Q), .A0(T15254_Y));
KC_AOI22_X1 T3758 ( .Y(T3758_Y), .B1(T10504_Y), .B0(T14414_Q),     .A1(T15215_Y), .A0(T14416_Q));
KC_AOI22_X1 T3759 ( .Y(T3759_Y), .B1(T14422_Q), .B0(T16442_Y),     .A1(T14431_Q), .A0(T15254_Y));
KC_AOI22_X1 T3764 ( .Y(T3764_Y), .B1(T14395_Q), .B0(T3117_Y),     .A1(T14417_Q), .A0(T12329_Y));
KC_AOI22_X1 T3765 ( .Y(T3765_Y), .B1(T14413_Q), .B0(T9936_Y),     .A1(T14430_Q), .A0(T9937_Y));
KC_AOI22_X1 T3766 ( .Y(T3766_Y), .B1(T14398_Q), .B0(T9936_Y),     .A1(T14418_Q), .A0(T9937_Y));
KC_AOI22_X1 T3767 ( .Y(T3767_Y), .B1(T5579_Y), .B0(T14395_Q),     .A1(T16443_Y), .A0(T14417_Q));
KC_AOI22_X1 T3768 ( .Y(T3768_Y), .B1(T5579_Y), .B0(T14397_Q),     .A1(T16443_Y), .A0(T14415_Q));
KC_AOI22_X1 T3769 ( .Y(T3769_Y), .B1(T5579_Y), .B0(T14361_Q),     .A1(T16443_Y), .A0(T14358_Q));
KC_AOI22_X1 T3770 ( .Y(T3770_Y), .B1(T10501_Y), .B0(T14413_Q),     .A1(T10502_Y), .A0(T14430_Q));
KC_AOI22_X1 T3771 ( .Y(T3771_Y), .B1(T14397_Q), .B0(T3117_Y),     .A1(T14415_Q), .A0(T12329_Y));
KC_AOI22_X1 T3772 ( .Y(T3772_Y), .B1(T10501_Y), .B0(T14398_Q),     .A1(T10502_Y), .A0(T14418_Q));
KC_AOI22_X1 T15847 ( .Y(T15847_Y), .B1(T11985_Y), .B0(T15558_Y),     .A1(T11317_Y), .A0(T11410_Y));
KC_AOI22_X1 T3793 ( .Y(T3793_Y), .B1(T6031_S), .B0(T4997_Y),     .A1(T6031_Co), .A0(T15554_Y));
KC_AOI22_X1 T3811 ( .Y(T3811_Y), .B1(T11378_Y), .B0(T15865_Y),     .A1(T11353_Y), .A0(T11379_Y));
KC_AOI22_X1 T3817 ( .Y(T3817_Y), .B1(T11316_Y), .B0(T11393_Y),     .A1(T11311_Y), .A0(T11427_Y));
KC_AOI22_X1 T3829 ( .Y(T3829_Y), .B1(T13087_Y), .B0(T11424_Y),     .A1(T5842_Y), .A0(T11426_Y));
KC_AOI22_X1 T3847 ( .Y(T3847_Y), .B1(T4461_Y), .B0(T11981_Y),     .A1(T6740_Y), .A0(T11410_Y));
KC_AOI22_X1 T3848 ( .Y(T3848_Y), .B1(T5760_Y), .B0(T11372_Y),     .A1(T5827_Y), .A0(T11378_Y));
KC_AOI22_X1 T3858 ( .Y(T3858_Y), .B1(T3246_Q), .B0(T5141_Y),     .A1(T4493_Q), .A0(T11506_Y));
KC_AOI22_X1 T3859 ( .Y(T3859_Y), .B1(T3258_Q), .B0(T5141_Y),     .A1(T3885_Q), .A0(T11506_Y));
KC_AOI22_X1 T3862 ( .Y(T3862_Y), .B1(T3227_Q), .B0(T5141_Y),     .A1(T5130_Q), .A0(T11506_Y));
KC_AOI22_X1 T3863 ( .Y(T3863_Y), .B1(T5075_Q), .B0(T5141_Y),     .A1(T3895_Q), .A0(T11506_Y));
KC_AOI22_X1 T3864 ( .Y(T3864_Y), .B1(T5439_Q), .B0(T5141_Y),     .A1(T4491_Q), .A0(T11506_Y));
KC_AOI22_X1 T3867 ( .Y(T3867_Y), .B1(T5076_Q), .B0(T5141_Y),     .A1(T3900_Q), .A0(T11506_Y));
KC_AOI22_X1 T3943 ( .Y(T3943_Y), .B1(T11536_Y), .B0(T5141_Y),     .A1(T12164_Y), .A0(T5985_Y));
KC_AOI22_X1 T4030 ( .Y(T4030_Y), .B1(T16029_Y), .B0(T5992_Y),     .A1(T12957_Y), .A0(T15610_Y));
KC_AOI22_X1 T4065 ( .Y(T4065_Y), .B1(T6174_Y), .B0(T5112_Y),     .A1(T4057_Y), .A0(T5135_Y));
KC_AOI22_X1 T4066 ( .Y(T4066_Y), .B1(T2806_Y), .B0(T8503_Y),     .A1(T10615_Y), .A0(T4106_Y));
KC_AOI22_X1 T4088 ( .Y(T4088_Y), .B1(T10586_Y), .B0(T11715_Y),     .A1(T4075_Y), .A0(T6094_Y));
KC_AOI22_X1 T4089 ( .Y(T4089_Y), .B1(T4075_Y), .B0(T10617_Y),     .A1(T11715_Y), .A0(T5135_Y));
KC_AOI22_X1 T4090 ( .Y(T4090_Y), .B1(T11745_Y), .B0(T10583_Y),     .A1(T11658_Y), .A0(T6094_Y));
KC_AOI22_X1 T6535 ( .Y(T6535_Y), .B1(T4146_Y), .B0(T6590_S),     .A1(T6611_S), .A0(T10568_Y));
KC_AOI22_X1 T4110 ( .Y(T4110_Y), .B1(T6205_Y), .B0(T6841_S),     .A1(T6574_Y), .A0(T6567_S));
KC_AOI22_X1 T4111 ( .Y(T4111_Y), .B1(T11687_Y), .B0(T6568_S),     .A1(T10566_Y), .A0(T6591_S));
KC_AOI22_X1 T4112 ( .Y(T4112_Y), .B1(T16125_Y), .B0(T6568_S),     .A1(T6591_S), .A0(T10542_Y));
KC_AOI22_X1 T4113 ( .Y(T4113_Y), .B1(T16125_Y), .B0(T6567_S),     .A1(T16142_Y), .A0(T5528_Q));
KC_AOI22_X1 T4114 ( .Y(T4114_Y), .B1(T3475_Y), .B0(T6841_S),     .A1(T2924_Y), .A0(T6238_Y));
KC_AOI22_X1 T4115 ( .Y(T4115_Y), .B1(T4964_Q), .B0(T10543_Y),     .A1(T11781_Y), .A0(T6526_Q));
KC_AOI22_X1 T4116 ( .Y(T4116_Y), .B1(T4146_Y), .B0(T6568_S),     .A1(T6591_S), .A0(T10568_Y));
KC_AOI22_X1 T4117 ( .Y(T4117_Y), .B1(T4150_Y), .B0(T6567_S),     .A1(T11781_Y), .A0(T5525_Q));
KC_AOI22_X1 T4118 ( .Y(T4118_Y), .B1(T11789_Y), .B0(T6586_Y),     .A1(T11792_Y), .A0(T10581_Y));
KC_AOI22_X1 T4120 ( .Y(T4120_Y), .B1(T6211_Y), .B0(T6547_Y),     .A1(T10568_Y), .A0(T6586_Y));
KC_AOI22_X1 T4121 ( .Y(T4121_Y), .B1(T6207_Y), .B0(T6237_Y),     .A1(T8422_Y), .A0(T15631_Y));
KC_AOI22_X1 T4122 ( .Y(T4122_Y), .B1(T13325_Y), .B0(T5532_Q),     .A1(T11781_Y), .A0(T6555_Q));
KC_AOI22_X1 T4123 ( .Y(T4123_Y), .B1(T2923_Y), .B0(T15631_Y),     .A1(T3469_Y), .A0(T4147_Q));
KC_AOI22_X1 T4124 ( .Y(T4124_Y), .B1(T8408_Y), .B0(T6238_Y),     .A1(T12054_Y), .A0(T16102_Y));
KC_AOI22_X1 T4125 ( .Y(T4125_Y), .B1(T2892_Y), .B0(T15631_Y),     .A1(T6237_Y), .A0(T4178_Q));
KC_AOI22_X1 T4126 ( .Y(T4126_Y), .B1(T2924_Y), .B0(T15631_Y),     .A1(T6562_Y), .A0(T6237_Y));
KC_AOI22_X1 T4129 ( .Y(T4129_Y), .B1(T11687_Y), .B0(T6503_S),     .A1(T10566_Y), .A0(T6614_S));
KC_AOI22_X1 T4130 ( .Y(T4130_Y), .B1(T13325_Y), .B0(T3528_Q),     .A1(T11781_Y), .A0(T6549_Q));
KC_AOI22_X1 T4131 ( .Y(T4131_Y), .B1(T6205_Y), .B0(T6840_S),     .A1(T6574_Y), .A0(T6534_S));
KC_AOI22_X1 T4132 ( .Y(T4132_Y), .B1(T11687_Y), .B0(T4540_Y),     .A1(T10566_Y), .A0(T4609_Y));
KC_AOI22_X1 T4133 ( .Y(T4133_Y), .B1(T16125_Y), .B0(T6503_S),     .A1(T6614_S), .A0(T10542_Y));
KC_AOI22_X1 T4134 ( .Y(T4134_Y), .B1(T11780_Y), .B0(T6586_Y),     .A1(T4107_Y), .A0(T10581_Y));
KC_AOI22_X1 T4135 ( .Y(T4135_Y), .B1(T6205_Y), .B0(T6504_S),     .A1(T6574_Y), .A0(T6533_S));
KC_AOI22_X1 T4136 ( .Y(T4136_Y), .B1(T11687_Y), .B0(T6590_S),     .A1(T10566_Y), .A0(T6611_S));
KC_AOI22_X1 T4137 ( .Y(T4137_Y), .B1(T16125_Y), .B0(T6590_S),     .A1(T6611_S), .A0(T10542_Y));
KC_AOI22_X1 T4141 ( .Y(T4141_Y), .B1(T4139_Y), .B0(T6840_S),     .A1(T4149_Y), .A0(T6534_S));
KC_AOI22_X1 T4142 ( .Y(T4142_Y), .B1(T3477_Y), .B0(T6842_S),     .A1(T11795_Y), .A0(T4171_Q));
KC_AOI22_X1 T4143 ( .Y(T4143_Y), .B1(T6210_Y), .B0(T6590_S),     .A1(T3469_Y), .A0(T4179_Q));
KC_AOI22_X1 T4144 ( .Y(T4144_Y), .B1(T4149_Y), .B0(T6533_S),     .A1(T4139_Y), .A0(T6504_S));
KC_AOI22_X1 T4152 ( .Y(T4152_Y), .B1(T8429_Y), .B0(T11817_Y),     .A1(T10593_Y), .A0(T4609_Y));
KC_AOI22_X1 T4154 ( .Y(T4154_Y), .B1(T5516_Y), .B0(T6547_Y),     .A1(T6591_S), .A0(T10593_Y));
KC_AOI22_X1 T4155 ( .Y(T4155_Y), .B1(T11734_Y), .B0(T6547_Y),     .A1(T6611_S), .A0(T10593_Y));
KC_AOI22_X1 T4160 ( .Y(T4160_Y), .B1(T4156_Y), .B0(T11842_Y),     .A1(T4166_Y), .A0(T9163_Y));
KC_AOI22_X1 T4182 ( .Y(T4182_Y), .B1(T13387_Q), .B0(T9635_Y),     .A1(T13402_Q), .A0(T5088_Y));
KC_AOI22_X1 T4183 ( .Y(T4183_Y), .B1(T9664_Y), .B0(T13418_Q),     .A1(T3610_Y), .A0(T13417_Q));
KC_AOI22_X1 T4217 ( .Y(T4217_Y), .B1(T9822_Y), .B0(T13761_Q),     .A1(T3635_Y), .A0(T13780_Q));
KC_AOI22_X1 T4218 ( .Y(T4218_Y), .B1(T9822_Y), .B0(T13760_Q),     .A1(T3635_Y), .A0(T13778_Q));
KC_AOI22_X1 T4219 ( .Y(T4219_Y), .B1(T14913_Q), .B0(T9867_Y),     .A1(T13779_Q), .A0(T5134_Y));
KC_AOI22_X1 T4220 ( .Y(T4220_Y), .B1(T13761_Q), .B0(T9867_Y),     .A1(T13780_Q), .A0(T5134_Y));
KC_AOI22_X1 T4221 ( .Y(T4221_Y), .B1(T9822_Y), .B0(T13749_Q),     .A1(T3635_Y), .A0(T13762_Q));
KC_AOI22_X1 T4222 ( .Y(T4222_Y), .B1(T13760_Q), .B0(T9867_Y),     .A1(T13778_Q), .A0(T5134_Y));
KC_AOI22_X1 T4230 ( .Y(T4230_Y), .B1(T14825_Q), .B0(T9864_Y),     .A1(T14824_Q), .A0(T9865_Y));
KC_AOI22_X1 T4233 ( .Y(T4233_Y), .B1(T9822_Y), .B0(T14848_Q),     .A1(T3635_Y), .A0(T14849_Q));
KC_AOI22_X1 T4234 ( .Y(T4234_Y), .B1(T14848_Q), .B0(T9867_Y),     .A1(T14849_Q), .A0(T5134_Y));
KC_AOI22_X1 T4235 ( .Y(T4235_Y), .B1(T9823_Y), .B0(T14844_Q),     .A1(T9825_Y), .A0(T14847_Q));
KC_AOI22_X1 T4236 ( .Y(T4236_Y), .B1(T14844_Q), .B0(T9864_Y),     .A1(T14847_Q), .A0(T9865_Y));
KC_AOI22_X1 T4237 ( .Y(T4237_Y), .B1(T14846_Q), .B0(T9866_Y),     .A1(T14037_Q), .A0(T15222_Y));
KC_AOI22_X1 T4238 ( .Y(T4238_Y), .B1(T14845_Q), .B0(T9863_Y),     .A1(T14851_Q), .A0(T9868_Y));
KC_AOI22_X1 T4239 ( .Y(T4239_Y), .B1(T9823_Y), .B0(T13875_Q),     .A1(T9825_Y), .A0(T13877_Q));
KC_AOI22_X1 T4241 ( .Y(T4241_Y), .B1(T9862_Y), .B0(T13906_Q),     .A1(T9824_Y), .A0(T13907_Q));
KC_AOI22_X1 T4242 ( .Y(T4242_Y), .B1(T13906_Q), .B0(T9863_Y),     .A1(T13907_Q), .A0(T9868_Y));
KC_AOI22_X1 T4243 ( .Y(T4243_Y), .B1(T13889_Q), .B0(T9864_Y),     .A1(T14820_Q), .A0(T9865_Y));
KC_AOI22_X1 T4244 ( .Y(T4244_Y), .B1(T9822_Y), .B0(T13891_Q),     .A1(T3635_Y), .A0(T14822_Q));
KC_AOI22_X1 T4245 ( .Y(T4245_Y), .B1(T9823_Y), .B0(T13889_Q),     .A1(T9825_Y), .A0(T14820_Q));
KC_AOI22_X1 T4246 ( .Y(T4246_Y), .B1(T13888_Q), .B0(T9866_Y),     .A1(T14823_Q), .A0(T15222_Y));
KC_AOI22_X1 T4247 ( .Y(T4247_Y), .B1(T12084_Y), .B0(T13888_Q),     .A1(T15219_Y), .A0(T14823_Q));
KC_AOI22_X1 T4248 ( .Y(T4248_Y), .B1(T13891_Q), .B0(T9867_Y),     .A1(T14822_Q), .A0(T5134_Y));
KC_AOI22_X1 T4249 ( .Y(T4249_Y), .B1(T14917_Q), .B0(T9864_Y),     .A1(T14910_Q), .A0(T9865_Y));
KC_AOI22_X1 T4253 ( .Y(T4253_Y), .B1(T9862_Y), .B0(T14845_Q),     .A1(T9824_Y), .A0(T14851_Q));
KC_AOI22_X1 T4254 ( .Y(T4254_Y), .B1(T9862_Y), .B0(T13878_Q),     .A1(T9824_Y), .A0(T13905_Q));
KC_AOI22_X1 T4255 ( .Y(T4255_Y), .B1(T13902_Q), .B0(T9866_Y),     .A1(T13872_Q), .A0(T15222_Y));
KC_AOI22_X1 T4256 ( .Y(T4256_Y), .B1(T13874_Q), .B0(T9867_Y),     .A1(T13901_Q), .A0(T5134_Y));
KC_AOI22_X1 T4257 ( .Y(T4257_Y), .B1(T9822_Y), .B0(T13874_Q),     .A1(T3635_Y), .A0(T13901_Q));
KC_AOI22_X1 T4258 ( .Y(T4258_Y), .B1(T9823_Y), .B0(T13900_Q),     .A1(T9825_Y), .A0(T13899_Q));
KC_AOI22_X1 T4259 ( .Y(T4259_Y), .B1(T12084_Y), .B0(T13902_Q),     .A1(T15219_Y), .A0(T13872_Q));
KC_AOI22_X1 T4260 ( .Y(T4260_Y), .B1(T13875_Q), .B0(T9864_Y),     .A1(T13877_Q), .A0(T9865_Y));
KC_AOI22_X1 T4261 ( .Y(T4261_Y), .B1(T13878_Q), .B0(T9863_Y),     .A1(T13905_Q), .A0(T9868_Y));
KC_AOI22_X1 T4262 ( .Y(T4262_Y), .B1(T13900_Q), .B0(T9864_Y),     .A1(T13899_Q), .A0(T9865_Y));
KC_AOI22_X1 T4263 ( .Y(T4263_Y), .B1(T9822_Y), .B0(T14085_Q),     .A1(T3635_Y), .A0(T14027_Q));
KC_AOI22_X1 T4264 ( .Y(T4264_Y), .B1(T14085_Q), .B0(T9867_Y),     .A1(T14027_Q), .A0(T16063_Y));
KC_AOI22_X1 T4269 ( .Y(T4269_Y), .B1(T14038_Q), .B0(T9867_Y),     .A1(T14063_Q), .A0(T16063_Y));
KC_AOI22_X1 T4270 ( .Y(T4270_Y), .B1(T9822_Y), .B0(T14038_Q),     .A1(T3635_Y), .A0(T14063_Q));
KC_AOI22_X1 T4273 ( .Y(T4273_Y), .B1(T14043_Q), .B0(T9864_Y),     .A1(T14042_Q), .A0(T9865_Y));
KC_AOI22_X1 T5855 ( .Y(T5855_Y), .B1(T9823_Y), .B0(T14175_Q),     .A1(T9825_Y), .A0(T14871_Q));
KC_AOI22_X1 T4287 ( .Y(T4287_Y), .B1(T14286_Q), .B0(T9866_Y),     .A1(T14887_Q), .A0(T15222_Y));
KC_AOI22_X1 T4288 ( .Y(T4288_Y), .B1(T14294_Q), .B0(T9863_Y),     .A1(T14290_Q), .A0(T9868_Y));
KC_AOI22_X1 T4289 ( .Y(T4289_Y), .B1(T14311_Q), .B0(T9866_Y),     .A1(T14287_Q), .A0(T15222_Y));
KC_AOI22_X1 T4292 ( .Y(T4292_Y), .B1(T12084_Y), .B0(T14286_Q),     .A1(T15219_Y), .A0(T14887_Q));
KC_AOI22_X1 T4293 ( .Y(T4293_Y), .B1(T9822_Y), .B0(T14330_Q),     .A1(T3635_Y), .A0(T14329_Q));
KC_AOI22_X1 T4294 ( .Y(T4294_Y), .B1(T9822_Y), .B0(T14186_Q),     .A1(T3635_Y), .A0(T14886_Q));
KC_AOI22_X1 T4295 ( .Y(T4295_Y), .B1(T14186_Q), .B0(T9867_Y),     .A1(T14886_Q), .A0(T16063_Y));
KC_AOI22_X1 T4296 ( .Y(T4296_Y), .B1(T14285_Q), .B0(T9863_Y),     .A1(T14885_Q), .A0(T9868_Y));
KC_AOI22_X1 T4297 ( .Y(T4297_Y), .B1(T9862_Y), .B0(T14285_Q),     .A1(T9824_Y), .A0(T14885_Q));
KC_AOI22_X1 T4298 ( .Y(T4298_Y), .B1(T9862_Y), .B0(T14294_Q),     .A1(T9824_Y), .A0(T14290_Q));
KC_AOI22_X1 T4299 ( .Y(T4299_Y), .B1(T12084_Y), .B0(T14311_Q),     .A1(T15219_Y), .A0(T14287_Q));
KC_AOI22_X1 T4300 ( .Y(T4300_Y), .B1(T9822_Y), .B0(T14156_Q),     .A1(T3635_Y), .A0(T14188_Q));
KC_AOI22_X1 T4301 ( .Y(T4301_Y), .B1(T14164_Q), .B0(T9864_Y),     .A1(T14159_Q), .A0(T9865_Y));
KC_AOI22_X1 T4302 ( .Y(T4302_Y), .B1(T9823_Y), .B0(T14164_Q),     .A1(T9825_Y), .A0(T14159_Q));
KC_AOI22_X1 T4303 ( .Y(T4303_Y), .B1(T9823_Y), .B0(T14155_Q),     .A1(T9825_Y), .A0(T14157_Q));
KC_AOI22_X1 T4304 ( .Y(T4304_Y), .B1(T14156_Q), .B0(T9867_Y),     .A1(T14188_Q), .A0(T16063_Y));
KC_AOI22_X1 T4305 ( .Y(T4305_Y), .B1(T14155_Q), .B0(T9864_Y),     .A1(T14157_Q), .A0(T9865_Y));
KC_AOI22_X1 T4308 ( .Y(T4308_Y), .B1(T14175_Q), .B0(T9864_Y),     .A1(T14871_Q), .A0(T9865_Y));
KC_AOI22_X1 T4309 ( .Y(T4309_Y), .B1(T14868_Q), .B0(T9866_Y),     .A1(T14869_Q), .A0(T15222_Y));
KC_AOI22_X1 T4310 ( .Y(T4310_Y), .B1(T14139_Q), .B0(T9867_Y),     .A1(T14177_Q), .A0(T16063_Y));
KC_AOI22_X1 T4311 ( .Y(T4311_Y), .B1(T9822_Y), .B0(T14139_Q),     .A1(T3635_Y), .A0(T14177_Q));
KC_AOI22_X1 T4312 ( .Y(T4312_Y), .B1(T14178_Q), .B0(T9866_Y),     .A1(T14176_Q), .A0(T15222_Y));
KC_AOI22_X1 T4313 ( .Y(T4313_Y), .B1(T12084_Y), .B0(T14178_Q),     .A1(T15219_Y), .A0(T14176_Q));
KC_AOI22_X1 T4314 ( .Y(T4314_Y), .B1(T12084_Y), .B0(T14868_Q),     .A1(T15219_Y), .A0(T14869_Q));
KC_AOI22_X1 T4315 ( .Y(T4315_Y), .B1(T9822_Y), .B0(T14872_Q),     .A1(T3635_Y), .A0(T14870_Q));
KC_AOI22_X1 T4316 ( .Y(T4316_Y), .B1(T14872_Q), .B0(T9867_Y),     .A1(T14870_Q), .A0(T16063_Y));
KC_AOI22_X1 T4319 ( .Y(T4319_Y), .B1(T14350_Q), .B0(T9932_Y),     .A1(T14349_Q), .A0(T3719_Y));
KC_AOI22_X1 T4320 ( .Y(T4320_Y), .B1(T10503_Y), .B0(T14350_Q),     .A1(T3684_Y), .A0(T14349_Q));
KC_AOI22_X1 T4321 ( .Y(T4321_Y), .B1(T9822_Y), .B0(T14306_Q),     .A1(T3635_Y), .A0(T14320_Q));
KC_AOI22_X1 T4322 ( .Y(T4322_Y), .B1(T9822_Y), .B0(T14351_Q),     .A1(T3635_Y), .A0(T14328_Q));
KC_AOI22_X1 T4323 ( .Y(T4323_Y), .B1(T9867_Y), .B0(T14306_Q),     .A1(T14320_Q), .A0(T16063_Y));
KC_AOI22_X1 T4324 ( .Y(T4324_Y), .B1(T14330_Q), .B0(T9867_Y),     .A1(T14329_Q), .A0(T16063_Y));
KC_AOI22_X1 T4325 ( .Y(T4325_Y), .B1(T14351_Q), .B0(T9867_Y),     .A1(T14328_Q), .A0(T16063_Y));
KC_AOI22_X1 T5975 ( .Y(T5975_Y), .B1(T14504_Q), .B0(T9932_Y),     .A1(T14896_Q), .A0(T3719_Y));
KC_AOI22_X1 T5974 ( .Y(T5974_Y), .B1(T10503_Y), .B0(T14504_Q),     .A1(T3684_Y), .A0(T14896_Q));
KC_AOI22_X1 T4338 ( .Y(T4338_Y), .B1(T10503_Y), .B0(T14895_Q),     .A1(T3684_Y), .A0(T14503_Q));
KC_AOI22_X1 T4339 ( .Y(T4339_Y), .B1(T14895_Q), .B0(T9932_Y),     .A1(T14503_Q), .A0(T3719_Y));
KC_AOI22_X1 T4340 ( .Y(T4340_Y), .B1(T14898_Q), .B0(T9932_Y),     .A1(T14437_Q), .A0(T3719_Y));
KC_AOI22_X1 T4341 ( .Y(T4341_Y), .B1(T10503_Y), .B0(T14898_Q),     .A1(T3684_Y), .A0(T14437_Q));
KC_AOI22_X1 T4342 ( .Y(T4342_Y), .B1(T10503_Y), .B0(T14434_Q),     .A1(T3684_Y), .A0(T14435_Q));
KC_AOI22_X1 T4343 ( .Y(T4343_Y), .B1(T14434_Q), .B0(T9932_Y),     .A1(T14435_Q), .A0(T3719_Y));
KC_AOI22_X1 T4344 ( .Y(T4344_Y), .B1(T10503_Y), .B0(T14407_Q),     .A1(T3684_Y), .A0(T14429_Q));
KC_AOI22_X1 T4345 ( .Y(T4345_Y), .B1(T14407_Q), .B0(T9932_Y),     .A1(T14429_Q), .A0(T3719_Y));
KC_AOI22_X1 T4346 ( .Y(T4346_Y), .B1(T10503_Y), .B0(T14410_Q),     .A1(T3684_Y), .A0(T14391_Q));
KC_AOI22_X1 T4347 ( .Y(T4347_Y), .B1(T10503_Y), .B0(T14411_Q),     .A1(T3684_Y), .A0(T14390_Q));
KC_AOI22_X1 T4348 ( .Y(T4348_Y), .B1(T14410_Q), .B0(T9932_Y),     .A1(T14391_Q), .A0(T3719_Y));
KC_AOI22_X1 T4349 ( .Y(T4349_Y), .B1(T14411_Q), .B0(T9932_Y),     .A1(T14390_Q), .A0(T3719_Y));
KC_AOI22_X1 T4385 ( .Y(T4385_Y), .B1(T4405_Y), .B0(T3856_Y),     .A1(T14942_Q), .A0(T6089_Y));
KC_AOI22_X1 T4390 ( .Y(T4390_Y), .B1(T3826_Y), .B0(T11312_Y),     .A1(T13078_Y), .A0(T4487_Q));
KC_AOI22_X1 T4391 ( .Y(T4391_Y), .B1(T14523_Q), .B0(T11401_Y),     .A1(T11349_Y), .A0(T15845_Y));
KC_AOI22_X1 T4398 ( .Y(T4398_Y), .B1(T5760_Y), .B0(T11982_Y),     .A1(T4438_Y), .A0(T15845_Y));
KC_AOI22_X1 T4399 ( .Y(T4399_Y), .B1(T15845_Y), .B0(T15871_Y),     .A1(T11312_Y), .A0(T16241_Y));
KC_AOI22_X1 T4400 ( .Y(T4400_Y), .B1(T11328_Y), .B0(T11393_Y),     .A1(T12144_Y), .A0(T15871_Y));
KC_AOI22_X1 T4401 ( .Y(T4401_Y), .B1(T4395_Y), .B0(T15832_Y),     .A1(T4418_Y), .A0(T4386_Y));
KC_AOI22_X1 T4404 ( .Y(T4404_Y), .B1(T5777_Y), .B0(T15871_Y),     .A1(T5760_Y), .A0(T16241_Y));
KC_AOI22_X1 T15900 ( .Y(T15900_Y), .B1(T13295_Y), .B0(T5789_Y),     .A1(T12952_Y), .A0(T5815_Y));
KC_AOI22_X1 T6113 ( .Y(T6113_Y), .B1(T13091_Y), .B0(T4438_Y),     .A1(T11420_Y), .A0(T5789_Y));
KC_AOI22_X1 T4434 ( .Y(T4434_Y), .B1(T11401_Y), .B0(T15871_Y),     .A1(T12801_Y), .A0(T15908_Y));
KC_AOI22_X1 T4435 ( .Y(T4435_Y), .B1(T11363_Y), .B0(T5788_Y),     .A1(T11394_Y), .A0(T11421_Y));
KC_AOI22_X1 T4443 ( .Y(T4443_Y), .B1(T11400_Y), .B0(T5830_Y),     .A1(T15558_Y), .A0(T14546_Q));
KC_AOI22_X1 T4444 ( .Y(T4444_Y), .B1(T4464_Y), .B0(T16154_Y),     .A1(T5767_Y), .A0(T11367_Y));
KC_AOI22_X1 T4449 ( .Y(T4449_Y), .B1(T15876_Y), .B0(T3856_Y),     .A1(T15869_Y), .A0(T5815_Y));
KC_AOI22_X1 T4450 ( .Y(T4450_Y), .B1(T10901_Y), .B0(T3836_Y),     .A1(T5760_Y), .A0(T6089_Y));
KC_AOI22_X1 T4562 ( .Y(T4562_Y), .B1(T11537_Y), .B0(T4517_Y),     .A1(T12014_Y), .A0(T4474_Y));
KC_AOI22_X1 T4598 ( .Y(T4598_Y), .B1(T8321_Y), .B0(T4617_Y),     .A1(T6325_Y), .A0(T12238_Y));
KC_AOI22_X1 T16323 ( .Y(T16323_Y), .B1(T16325_Y), .B0(T7574_Y),     .A1(T7569_Y), .A0(T16329_Y));
KC_AOI22_X1 T16322 ( .Y(T16322_Y), .B1(T7824_Y), .B0(T15655_Y),     .A1(T16319_Y), .A0(T16325_Y));
KC_AOI22_X1 T6725 ( .Y(T6725_Y), .B1(T11864_Y), .B0(T167_Q),     .A1(T6801_Y), .A0(T163_Q));
KC_AOI22_X1 T6718 ( .Y(T6718_Y), .B1(T8389_Y), .B0(T319_Q),     .A1(T15739_Y), .A0(T165_Q));
KC_AOI22_X1 T6717 ( .Y(T6717_Y), .B1(T12426_Y), .B0(T5559_Q),     .A1(T12424_Y), .A0(T320_Q));
KC_AOI22_X1 T6715 ( .Y(T6715_Y), .B1(T12399_Y), .B0(T163_Q),     .A1(T12425_Y), .A0(T5252_Q));
KC_AOI22_X1 T6680 ( .Y(T6680_Y), .B1(T15739_Y), .B0(T363_Q),     .A1(T8389_Y), .A0(T524_Q));
KC_AOI22_X1 T6476 ( .Y(T6476_Y), .B1(T6818_Y), .B0(T153_Q),     .A1(T6828_Y), .A0(T5564_Q));
KC_AOI22_X1 T6472 ( .Y(T6472_Y), .B1(T12423_Y), .B0(T157_Q),     .A1(T12407_Y), .A0(T153_Q));
KC_AOI22_X1 T6268 ( .Y(T6268_Y), .B1(T6801_Y), .B0(T5243_Q),     .A1(T11864_Y), .A0(T4822_Q));
KC_AOI22_X1 T270 ( .Y(T270_Y), .B1(T12423_Y), .B0(T284_Q),     .A1(T12408_Y), .A0(T5226_Q));
KC_AOI22_X1 T16342 ( .Y(T16342_Y), .B1(T8735_Y), .B0(T554_Y),     .A1(T641_Y), .A0(T517_Q));
KC_AOI22_X1 T16341 ( .Y(T16341_Y), .B1(T8735_Y), .B0(T5537_Y),     .A1(T641_Y), .A0(T4827_Q));
KC_AOI22_X1 T16340 ( .Y(T16340_Y), .B1(T8735_Y), .B0(T2130_Y),     .A1(T641_Y), .A0(T512_Q));
KC_AOI22_X1 T6709 ( .Y(T6709_Y), .B1(T15310_Y), .B0(T5276_Q),     .A1(T6799_Y), .A0(T4799_Q));
KC_AOI22_X1 T6701 ( .Y(T6701_Y), .B1(T6829_Y), .B0(T5560_Q),     .A1(T6597_Y), .A0(T664_Q));
KC_AOI22_X1 T6668 ( .Y(T6668_Y), .B1(T922_Y), .B0(T523_Q),     .A1(T16116_Y), .A0(T519_Q));
KC_AOI22_X1 T6667 ( .Y(T6667_Y), .B1(T15734_Y), .B0(T363_Q),     .A1(T12427_Y), .A0(T5305_Q));
KC_AOI22_X1 T6661 ( .Y(T6661_Y), .B1(T922_Y), .B0(T5306_Q),     .A1(T16116_Y), .A0(T5305_Q));
KC_AOI22_X1 T6660 ( .Y(T6660_Y), .B1(T600_Y), .B0(T5283_Q),     .A1(T12435_Y), .A0(T5306_Q));
KC_AOI22_X1 T6349 ( .Y(T6349_Y), .B1(T600_Y), .B0(T4835_Q),     .A1(T12435_Y), .A0(T7085_Q));
KC_AOI22_X1 T6267 ( .Y(T6267_Y), .B1(T12425_Y), .B0(T278_Q),     .A1(T12406_Y), .A0(T5221_Q));
KC_AOI22_X1 T6263 ( .Y(T6263_Y), .B1(T12399_Y), .B0(T439_Q),     .A1(T12405_Y), .A0(T438_Q));
KC_AOI22_X1 T6262 ( .Y(T6262_Y), .B1(T6799_Y), .B0(T273_Q),     .A1(T15310_Y), .A0(T5221_Q));
KC_AOI22_X1 T6259 ( .Y(T6259_Y), .B1(T6264_Y), .B0(T438_Q),     .A1(T6288_Y), .A0(T627_Q));
KC_AOI22_X1 T16347 ( .Y(T16347_Y), .B1(T5358_Y), .B0(T956_Y),     .A1(T8756_Y), .A0(T8831_Y));
KC_AOI22_X1 T16344 ( .Y(T16344_Y), .B1(T9371_Y), .B0(T2242_Y),     .A1(T904_Y), .A0(T716_Q));
KC_AOI22_X1 T6697 ( .Y(T6697_Y), .B1(T600_Y), .B0(T6487_Q),     .A1(T12435_Y), .A0(T669_Q));
KC_AOI22_X1 T6696 ( .Y(T6696_Y), .B1(T12409_Y), .B0(T5262_Q),     .A1(T12407_Y), .A0(T4836_Q));
KC_AOI22_X1 T6695 ( .Y(T6695_Y), .B1(T12429_Y), .B0(T862_Q),     .A1(T12427_Y), .A0(T696_Q));
KC_AOI22_X1 T6658 ( .Y(T6658_Y), .B1(T12426_Y), .B0(T5309_Q),     .A1(T12424_Y), .A0(T1066_Q));
KC_AOI22_X1 T6657 ( .Y(T6657_Y), .B1(T12425_Y), .B0(T705_Q),     .A1(T12406_Y), .A0(T1046_Q));
KC_AOI22_X1 T6656 ( .Y(T6656_Y), .B1(T12426_Y), .B0(T935_Q),     .A1(T12424_Y), .A0(T1068_Q));
KC_AOI22_X1 T6328 ( .Y(T6328_Y), .B1(T922_Y), .B0(T5206_Q),     .A1(T16116_Y), .A0(T653_Q));
KC_AOI22_X1 T6323 ( .Y(T6323_Y), .B1(T12399_Y), .B0(T829_Q),     .A1(T12405_Y), .A0(T679_Q));
KC_AOI22_X1 T6322 ( .Y(T6322_Y), .B1(T600_Y), .B0(T5238_Q),     .A1(T12435_Y), .A0(T674_Q));
KC_AOI22_X1 T6255 ( .Y(T6255_Y), .B1(T12399_Y), .B0(T822_Q),     .A1(T12405_Y), .A0(T5199_Q));
KC_AOI22_X1 T6254 ( .Y(T6254_Y), .B1(T12399_Y), .B0(T790_Q),     .A1(T12405_Y), .A0(T627_Q));
KC_AOI22_X1 T16349 ( .Y(T16349_Y), .B1(T956_Y), .B0(T8772_Y),     .A1(T9365_Y), .A0(T8831_Y));
KC_AOI22_X1 T16279 ( .Y(T16279_Y), .B1(T1158_Q), .B0(T9032_Y),     .A1(T8997_Y), .A0(T1012_Q));
KC_AOI22_X1 T6690 ( .Y(T6690_Y), .B1(T11193_Y), .B0(T9298_Y),     .A1(T15781_Y), .A0(T715_Y));
KC_AOI22_X1 T6649 ( .Y(T6649_Y), .B1(T9330_Y), .B0(T637_Y),     .A1(T6650_Y), .A0(T1068_Q));
KC_AOI22_X1 T6038 ( .Y(T6038_Y), .B1(T922_Y), .B0(T674_Q),     .A1(T16116_Y), .A0(T828_Q));
KC_AOI22_X1 T6795 ( .Y(T6795_Y), .B1(T12706_Y), .B0(T715_Y),     .A1(T11171_Y), .A0(T9300_Y));
KC_AOI22_X1 T10869 ( .Y(T10869_Y), .B1(T14583_Q), .B0(T9576_Y),     .A1(T14585_Q), .A0(T15237_Y));
KC_AOI22_X1 T10868 ( .Y(T10868_Y), .B1(T9585_Y), .B0(T14583_Q),     .A1(T15197_Y), .A0(T14585_Q));
KC_AOI22_X1 T10831 ( .Y(T10831_Y), .B1(T10420_Y), .B0(T14672_Q),     .A1(T10423_Y), .A0(T14673_Q));
KC_AOI22_X1 T10828 ( .Y(T10828_Y), .B1(T7231_Y), .B0(T15220_Y),     .A1(T10374_Y), .A0(T12086_Y));
KC_AOI22_X1 T10827 ( .Y(T10827_Y), .B1(T13841_Q), .B0(T10421_Y),     .A1(T14669_Q), .A0(T15194_Y));
KC_AOI22_X1 T10826 ( .Y(T10826_Y), .B1(T10418_Y), .B0(T13841_Q),     .A1(T15248_Y), .A0(T14669_Q));
KC_AOI22_X1 T10825 ( .Y(T10825_Y), .B1(T6794_Q), .B0(T1344_Y),     .A1(T13831_Q), .A0(T1343_Y));
KC_AOI22_X1 T10824 ( .Y(T10824_Y), .B1(T10368_Y), .B0(T6794_Q),     .A1(T10366_Y), .A0(T13831_Q));
KC_AOI22_X1 T10815 ( .Y(T10815_Y), .B1(T13825_Q), .B0(T10422_Y),     .A1(T13823_Q), .A0(T10367_Y));
KC_AOI22_X1 T10814 ( .Y(T10814_Y), .B1(T13821_Q), .B0(T10422_Y),     .A1(T13839_Q), .A0(T10367_Y));
KC_AOI22_X1 T10813 ( .Y(T10813_Y), .B1(T7206_Y), .B0(T15220_Y),     .A1(T5678_Y), .A0(T12086_Y));
KC_AOI22_X1 T10794 ( .Y(T10794_Y), .B1(T14649_Q), .B0(T12327_Y),     .A1(T14652_Q), .A0(T10788_Y));
KC_AOI22_X1 T10791 ( .Y(T10791_Y), .B1(T10368_Y), .B0(T14651_Q),     .A1(T10366_Y), .A0(T14647_Q));
KC_AOI22_X1 T10790 ( .Y(T10790_Y), .B1(T14650_Q), .B0(T1344_Y),     .A1(T14644_Q), .A0(T1343_Y));
KC_AOI22_X1 T6793 ( .Y(T6793_Y), .B1(T7025_Y), .B0(T15220_Y),     .A1(T10371_Y), .A0(T12086_Y));
KC_AOI22_X1 T10816 ( .Y(T10816_Y), .B1(T10368_Y), .B0(T14748_Q),     .A1(T10366_Y), .A0(T14750_Q));
KC_AOI22_X1 T10812 ( .Y(T10812_Y), .B1(T7016_Y), .B0(T15220_Y),     .A1(T10370_Y), .A0(T12086_Y));
KC_AOI22_X1 T10811 ( .Y(T10811_Y), .B1(T14748_Q), .B0(T1344_Y),     .A1(T14750_Q), .A0(T1343_Y));
KC_AOI22_X1 T10789 ( .Y(T10789_Y), .B1(T14646_Q), .B0(T12327_Y),     .A1(T14639_Q), .A0(T10788_Y));
KC_AOI22_X1 T10786 ( .Y(T10786_Y), .B1(T12327_Y), .B0(T14641_Q),     .A1(T13999_Q), .A0(T10788_Y));
KC_AOI22_X1 T10741 ( .Y(T10741_Y), .B1(T12094_Y), .B0(T14597_Q),     .A1(T8000_Y), .A0(T14213_Q));
KC_AOI22_X1 T16441 ( .Y(T16441_Y), .B1(T8013_Y), .B0(T14612_Q),     .A1(T7711_Y), .A0(T2565_Y));
KC_AOI22_X1 T10809 ( .Y(T10809_Y), .B1(T10808_Y), .B0(T14661_Q),     .A1(T10369_Y), .A0(T2565_Y));
KC_AOI22_X1 T10878 ( .Y(T10878_Y), .B1(T7176_Y), .B0(T13583_Q),     .A1(T5662_Y), .A0(T9642_Y));
KC_AOI22_X1 T10877 ( .Y(T10877_Y), .B1(T9580_Y), .B0(T14721_Q),     .A1(T3640_Y), .A0(T14723_Q));
KC_AOI22_X1 T10867 ( .Y(T10867_Y), .B1(T14705_Q), .B0(T12075_Y),     .A1(T14704_Q), .A0(T7323_Y));
KC_AOI22_X1 T10866 ( .Y(T10866_Y), .B1(T9580_Y), .B0(T13604_Q),     .A1(T2027_Y), .A0(T13605_Q));
KC_AOI22_X1 T10803 ( .Y(T10803_Y), .B1(T14663_Q), .B0(T10358_Y),     .A1(T14741_Q), .A0(T9712_Y));
KC_AOI22_X1 T10802 ( .Y(T10802_Y), .B1(T10346_Y), .B0(T13715_Q),     .A1(T15245_Y), .A0(T13733_Q));
KC_AOI22_X1 T10801 ( .Y(T10801_Y), .B1(T9704_Y), .B0(T14663_Q),     .A1(T9705_Y), .A0(T14741_Q));
KC_AOI22_X1 T10797 ( .Y(T10797_Y), .B1(T10346_Y), .B0(T13735_Q),     .A1(T15245_Y), .A0(T13731_Q));
KC_AOI22_X1 T10796 ( .Y(T10796_Y), .B1(T13735_Q), .B0(T10361_Y),     .A1(T13731_Q), .A0(T15247_Y));
KC_AOI22_X1 T10782 ( .Y(T10782_Y), .B1(T9704_Y), .B0(T13785_Q),     .A1(T9705_Y), .A0(T13851_Q));
KC_AOI22_X1 T10781 ( .Y(T10781_Y), .B1(T7757_Y), .B0(T12086_Y),     .A1(T10363_Y), .A0(T2531_Y));
KC_AOI22_X1 T10780 ( .Y(T10780_Y), .B1(T14011_Q), .B0(T10361_Y),     .A1(T13955_Q), .A0(T15247_Y));
KC_AOI22_X1 T10779 ( .Y(T10779_Y), .B1(T13992_Q), .B0(T10362_Y),     .A1(T13991_Q), .A0(T10360_Y));
KC_AOI22_X1 T10778 ( .Y(T10778_Y), .B1(T13954_Q), .B0(T10362_Y),     .A1(T16178_Q), .A0(T10360_Y));
KC_AOI22_X1 T10777 ( .Y(T10777_Y), .B1(T14633_Q), .B0(T10358_Y),     .A1(T14632_Q), .A0(T9712_Y));
KC_AOI22_X1 T10776 ( .Y(T10776_Y), .B1(T9704_Y), .B0(T13996_Q),     .A1(T9705_Y), .A0(T13976_Q));
KC_AOI22_X1 T10770 ( .Y(T10770_Y), .B1(T14629_Q), .B0(T10359_Y),     .A1(T14627_Q), .A0(T4889_Y));
KC_AOI22_X1 T10766 ( .Y(T10766_Y), .B1(T9706_Y), .B0(T14629_Q),     .A1(T1545_Y), .A0(T14627_Q));
KC_AOI22_X1 T10759 ( .Y(T10759_Y), .B1(T10758_Y), .B0(T14607_Q),     .A1(T7991_Y), .A0(T2565_Y));
KC_AOI22_X1 T4893 ( .Y(T4893_Y), .B1(T12094_Y), .B0(T14458_Q),     .A1(T8000_Y), .A0(T14457_Q));
KC_AOI22_X1 T10876 ( .Y(T10876_Y), .B1(T10397_Y), .B0(T6461_Q),     .A1(T15204_Y), .A0(T13581_Q));
KC_AOI22_X1 T10875 ( .Y(T10875_Y), .B1(T12325_Y), .B0(T13686_Q),     .A1(T12324_Y), .A0(T13711_Q));
KC_AOI22_X1 T10874 ( .Y(T10874_Y), .B1(T12076_Y), .B0(T13686_Q),     .A1(T12074_Y), .A0(T13711_Q));
KC_AOI22_X1 T10769 ( .Y(T10769_Y), .B1(T13985_Q), .B0(T10359_Y),     .A1(T13990_Q), .A0(T4889_Y));
KC_AOI22_X1 T10768 ( .Y(T10768_Y), .B1(T14630_Q), .B0(T10359_Y),     .A1(T14631_Q), .A0(T4889_Y));
KC_AOI22_X1 T10767 ( .Y(T10767_Y), .B1(T9706_Y), .B0(T13972_Q),     .A1(T1545_Y), .A0(T13988_Q));
KC_AOI22_X1 T10742 ( .Y(T10742_Y), .B1(T2038_Y), .B0(T1450_Y),     .A1(T10525_Y), .A0(T16413_Q));
KC_AOI22_X1 T4906 ( .Y(T4906_Y), .B1(T2038_Y), .B0(T1724_Y),     .A1(T10525_Y), .A0(T1707_Q));
KC_AOI22_X1 T4907 ( .Y(T4907_Y), .B1(T9706_Y), .B0(T14075_Q),     .A1(T1545_Y), .A0(T10247_Q));
KC_AOI22_X1 T4908 ( .Y(T4908_Y), .B1(T14075_Q), .B0(T10359_Y),     .A1(T10247_Q), .A0(T4889_Y));
KC_AOI22_X1 T4909 ( .Y(T4909_Y), .B1(T14841_Q), .B0(T10361_Y),     .A1(T13923_Q), .A0(T15247_Y));
KC_AOI22_X1 T4910 ( .Y(T4910_Y), .B1(T13599_Q), .B0(T1547_Y),     .A1(T13601_Q), .A0(T15202_Y));
KC_AOI22_X1 T4913 ( .Y(T4913_Y), .B1(T1826_Q), .B0(T12269_Y),     .A1(T1803_Q), .A0(T6164_Y));
KC_AOI22_X1 T4914 ( .Y(T4914_Y), .B1(T1790_Q), .B0(T12269_Y),     .A1(T1785_Q), .A0(T6164_Y));
KC_AOI22_X1 T4915 ( .Y(T4915_Y), .B1(T1787_Q), .B0(T12269_Y),     .A1(T1790_Q), .A0(T12270_Y));
KC_AOI22_X1 T4938 ( .Y(T4938_Y), .B1(T11620_Y), .B0(T2112_Q),     .A1(T2182_Q), .A0(T11586_Y));
KC_AOI22_X1 T4939 ( .Y(T4939_Y), .B1(T2186_Q), .B0(T11586_Y),     .A1(T11012_Y), .A0(T11551_Y));
KC_AOI22_X1 T4940 ( .Y(T4940_Y), .B1(T13108_Q), .B0(T12030_Y),     .A1(T5481_Q), .A0(T5990_Y));
KC_AOI22_X1 T4941 ( .Y(T4941_Y), .B1(T2114_Q), .B0(T5848_Y),     .A1(T1753_Q), .A0(T11499_Y));
KC_AOI22_X1 T4944 ( .Y(T4944_Y), .B1(T5455_Q), .B0(T5944_Y),     .A1(T4970_Q), .A0(T5909_Y));
KC_AOI22_X1 T4945 ( .Y(T4945_Y), .B1(T5443_Y), .B0(T11499_Y),     .A1(T11480_Y), .A0(T8447_Y));
KC_AOI22_X1 T4952 ( .Y(T4952_Y), .B1(T4968_Y), .B0(T12268_Y),     .A1(T2345_Q), .A0(T11728_Y));
KC_AOI22_X1 T4953 ( .Y(T4953_Y), .B1(T2714_Y), .B0(T12268_Y),     .A1(T11728_Y), .A0(T2316_Q));
KC_AOI22_X1 T4956 ( .Y(T4956_Y), .B1(T9162_Y), .B0(T6015_Y),     .A1(T2671_Y), .A0(T15232_Y));
KC_AOI22_X1 T4957 ( .Y(T4957_Y), .B1(T15608_Y), .B0(T16009_Y),     .A1(T2243_Y), .A0(T6013_Y));
KC_AOI22_X1 T4958 ( .Y(T4958_Y), .B1(T2238_Y), .B0(T16096_Y),     .A1(T2851_Y), .A0(T12103_Y));
KC_AOI22_X1 T4959 ( .Y(T4959_Y), .B1(T2673_Y), .B0(T6015_Y),     .A1(T2134_Y), .A0(T11551_Y));
KC_AOI22_X1 T4961 ( .Y(T4961_Y), .B1(T2237_Q), .B0(T2876_Y),     .A1(T11728_Y), .A0(T16082_Q));
KC_AOI22_X1 T16256 ( .Y(T16256_Y), .B1(T5951_Y), .B0(T14366_Q),     .A1(T3161_Y), .A0(T14994_Y));
KC_AOI22_X1 T4988 ( .Y(T4988_Y), .B1(T7504_Y), .B0(T2531_Y),     .A1(T4290_Y), .A0(T16165_Y));
KC_AOI22_X1 T4989 ( .Y(T4989_Y), .B1(T2412_Y), .B0(T2535_Y),     .A1(T3545_Y), .A0(T2532_Y));
KC_AOI22_X1 T4990 ( .Y(T4990_Y), .B1(T6637_Y), .B0(T13782_Q),     .A1(T2973_Y), .A0(T4937_Y));
KC_AOI22_X1 T5000 ( .Y(T5000_Y), .B1(T3436_Y), .B0(T10546_Y),     .A1(T2899_Y), .A0(T10555_Y));
KC_AOI22_X1 T5001 ( .Y(T5001_Y), .B1(T3436_Y), .B0(T10546_Y),     .A1(T11688_Y), .A0(T12317_Y));
KC_AOI22_X1 T5005 ( .Y(T5005_Y), .B1(T3436_Y), .B0(T12048_Y),     .A1(T6073_Y), .A0(T12104_Y));
KC_AOI22_X1 T5006 ( .Y(T5006_Y), .B1(T12048_Y), .B0(T6182_Y),     .A1(T2851_Y), .A0(T12104_Y));
KC_AOI22_X1 T5007 ( .Y(T5007_Y), .B1(T8480_Y), .B0(T12009_Y),     .A1(T5069_Y), .A0(T15805_Q));
KC_AOI22_X1 T16259 ( .Y(T16259_Y), .B1(T5579_Y), .B0(T14364_Q),     .A1(T16443_Y), .A0(T14359_Q));
KC_AOI22_X1 T5031 ( .Y(T5031_Y), .B1(T9731_Y), .B0(T14047_Q),     .A1(T3640_Y), .A0(T14046_Q));
KC_AOI22_X1 T5032 ( .Y(T5032_Y), .B1(T9731_Y), .B0(T14044_Q),     .A1(T3640_Y), .A0(T14068_Q));
KC_AOI22_X1 T5035 ( .Y(T5035_Y), .B1(T13625_Q), .B0(T9637_Y),     .A1(T13626_Q), .A0(T6483_Y));
KC_AOI22_X1 T5036 ( .Y(T5036_Y), .B1(T10436_Y), .B0(T13625_Q),     .A1(T10437_Y), .A0(T13626_Q));
KC_AOI22_X1 T5043 ( .Y(T5043_Y), .B1(T3228_Q), .B0(T5141_Y),     .A1(T5129_Q), .A0(T11506_Y));
KC_AOI22_X1 T5085 ( .Y(T5085_Y), .B1(T12084_Y), .B0(T14828_Q),     .A1(T15219_Y), .A0(T14916_Q));
KC_AOI22_X1 T5086 ( .Y(T5086_Y), .B1(T9823_Y), .B0(T14921_Q),     .A1(T9825_Y), .A0(T14911_Q));
KC_AOI22_X1 T5087 ( .Y(T5087_Y), .B1(T12084_Y), .B0(T14826_Q),     .A1(T15219_Y), .A0(T14920_Q));
KC_AOI22_X1 T5089 ( .Y(T5089_Y), .B1(T13622_Q), .B0(T9665_Y),     .A1(T14779_Q), .A0(T15256_Y));
KC_AOI22_X1 T5090 ( .Y(T5090_Y), .B1(T3024_Y), .B0(T13622_Q),     .A1(T15211_Y), .A0(T14779_Q));
KC_AOI22_X1 T5091 ( .Y(T5091_Y), .B1(T3027_Y), .B0(T14794_Q),     .A1(T9636_Y), .A0(T14778_Q));
KC_AOI22_X1 T5092 ( .Y(T5092_Y), .B1(T14794_Q), .B0(T3611_Y),     .A1(T14778_Q), .A0(T6482_Y));
KC_AOI22_X1 T5093 ( .Y(T5093_Y), .B1(T3027_Y), .B0(T14760_Q),     .A1(T9636_Y), .A0(T13646_Q));
KC_AOI22_X1 T5094 ( .Y(T5094_Y), .B1(T3027_Y), .B0(T14759_Q),     .A1(T9636_Y), .A0(T13649_Q));
KC_AOI22_X1 T5095 ( .Y(T5095_Y), .B1(T3027_Y), .B0(T14763_Q),     .A1(T9636_Y), .A0(T13650_Q));
KC_AOI22_X1 T5096 ( .Y(T5096_Y), .B1(T14759_Q), .B0(T3611_Y),     .A1(T13649_Q), .A0(T6482_Y));
KC_AOI22_X1 T5097 ( .Y(T5097_Y), .B1(T3611_Y), .B0(T14760_Q),     .A1(T6482_Y), .A0(T13646_Q));
KC_AOI22_X1 T5098 ( .Y(T5098_Y), .B1(T14763_Q), .B0(T3611_Y),     .A1(T13650_Q), .A0(T6482_Y));
KC_AOI22_X1 T5102 ( .Y(T5102_Y), .B1(T11978_Y), .B0(T11427_Y),     .A1(T12159_Y), .A0(T15877_Y));
KC_AOI22_X1 T5103 ( .Y(T5103_Y), .B1(T5760_Y), .B0(T11353_Y),     .A1(T4403_Y), .A0(T11402_Y));
KC_AOI22_X1 T5104 ( .Y(T5104_Y), .B1(T6740_Y), .B0(T11376_Y),     .A1(T15868_Y), .A0(T11367_Y));
KC_AOI22_X1 T5106 ( .Y(T5106_Y), .B1(T12181_Y), .B0(T11969_Y),     .A1(T3853_Y), .A0(T14494_Q));
KC_AOI22_X1 T5110 ( .Y(T5110_Y), .B1(T11687_Y), .B0(T6842_S),     .A1(T10566_Y), .A0(T6610_S));
KC_AOI22_X1 T5136 ( .Y(T5136_Y), .B1(T12084_Y), .B0(T14846_Q),     .A1(T15219_Y), .A0(T14037_Q));
KC_AOI22_X1 T5137 ( .Y(T5137_Y), .B1(T13749_Q), .B0(T9867_Y),     .A1(T13762_Q), .A0(T5134_Y));
KC_AOI22_X1 T5138 ( .Y(T5138_Y), .B1(T9822_Y), .B0(T14913_Q),     .A1(T3635_Y), .A0(T13779_Q));
KC_AOI22_X1 T6886 ( .Y(T6886_Y), .B1(T9579_Y), .B0(T13356_Q),     .A1(T14980_Y), .A0(T13383_Q));
KC_AOI22_X1 T6859 ( .Y(T6859_Y), .B1(T6855_S), .B0(T6855_S),     .A1(T6855_Co), .A0(T6855_S));
KC_AOI22_X1 T5177 ( .Y(T5177_Y), .B1(T9664_Y), .B0(T13506_Q),     .A1(T3610_Y), .A0(T13507_Q));
KC_AOI22_X1 T5178 ( .Y(T5178_Y), .B1(T15045_Q), .B0(T12075_Y),     .A1(T13416_Q), .A0(T7323_Y));
KC_AOI22_X1 T5179 ( .Y(T5179_Y), .B1(T13409_Q), .B0(T9635_Y),     .A1(T13408_Q), .A0(T5088_Y));
KC_AOI22_X1 T5180 ( .Y(T5180_Y), .B1(T9664_Y), .B0(T13392_Q),     .A1(T3610_Y), .A0(T13393_Q));
KC_AOI22_X1 T5181 ( .Y(T5181_Y), .B1(T9664_Y), .B0(T13409_Q),     .A1(T3610_Y), .A0(T13408_Q));
KC_AOI22_X1 T5182 ( .Y(T5182_Y), .B1(T9664_Y), .B0(T13387_Q),     .A1(T3610_Y), .A0(T13402_Q));
KC_AOI22_X1 T6298 ( .Y(T6298_Y), .B1(T12399_Y), .B0(T5205_Q),     .A1(T12405_Y), .A0(T5196_Q));
KC_AOI22_X1 T10847 ( .Y(T10847_Y), .B1(T12325_Y), .B0(T14686_Q),     .A1(T12324_Y), .A0(T14685_Q));
KC_AOI22_X1 T7037 ( .Y(T7037_Y), .B1(T13493_Q), .B0(T12076_Y),     .A1(T16505_Y), .A0(T12074_Y));
KC_AOI22_X1 T7032 ( .Y(T7032_Y), .B1(T13485_Q), .B0(T9578_Y),     .A1(T13486_Q), .A0(T12073_Y));
KC_AOI22_X1 T7030 ( .Y(T7030_Y), .B1(T9575_Y), .B0(T13485_Q),     .A1(T9586_Y), .A0(T13486_Q));
KC_AOI22_X1 T6995 ( .Y(T6995_Y), .B1(T13452_Q), .B0(T9578_Y),     .A1(T13481_Q), .A0(T12073_Y));
KC_AOI22_X1 T6975 ( .Y(T6975_Y), .B1(T13465_Q), .B0(T12077_Y),     .A1(T13494_Q), .A0(T12078_Y));
KC_AOI22_X1 T6955 ( .Y(T6955_Y), .B1(T7364_Y), .B0(T442_Q),     .A1(T8384_Y), .A0(T5227_Q));
KC_AOI22_X1 T6929 ( .Y(T6929_Y), .B1(T12409_Y), .B0(T288_Q),     .A1(T12407_Y), .A0(T283_Q));
KC_AOI22_X1 T6921 ( .Y(T6921_Y), .B1(T12423_Y), .B0(T442_Q),     .A1(T12408_Y), .A0(T446_Q));
KC_AOI22_X1 T5207 ( .Y(T5207_Y), .B1(T13537_Q), .B0(T12076_Y),     .A1(T13518_Q), .A0(T12074_Y));
KC_AOI22_X1 T5209 ( .Y(T5209_Y), .B1(T14800_Q), .B0(T9637_Y),     .A1(T13556_Q), .A0(T6483_Y));
KC_AOI22_X1 T5210 ( .Y(T5210_Y), .B1(T13553_Q), .B0(T9635_Y),     .A1(T13552_Q), .A0(T5088_Y));
KC_AOI22_X1 T5211 ( .Y(T5211_Y), .B1(T13538_Q), .B0(T12077_Y),     .A1(T13517_Q), .A0(T12078_Y));
KC_AOI22_X1 T5212 ( .Y(T5212_Y), .B1(T13530_Q), .B0(T1547_Y),     .A1(T13532_Q), .A0(T15202_Y));
KC_AOI22_X1 T5213 ( .Y(T5213_Y), .B1(T9664_Y), .B0(T13524_Q),     .A1(T3610_Y), .A0(T14797_Q));
KC_AOI22_X1 T5214 ( .Y(T5214_Y), .B1(T13524_Q), .B0(T9635_Y),     .A1(T14797_Q), .A0(T5088_Y));
KC_AOI22_X1 T5215 ( .Y(T5215_Y), .B1(T9664_Y), .B0(T13553_Q),     .A1(T3610_Y), .A0(T13552_Q));
KC_AOI22_X1 T5216 ( .Y(T5216_Y), .B1(T9664_Y), .B0(T13423_Q),     .A1(T3610_Y), .A0(T14814_Q));
KC_AOI22_X1 T12389 ( .Y(T12389_Y), .B1(T15734_Y), .B0(T831_Q),     .A1(T15735_Y), .A0(T5195_Q));
KC_AOI22_X1 T7197 ( .Y(T7197_Y), .B1(T9585_Y), .B0(T14733_Q),     .A1(T15197_Y), .A0(T14730_Q));
KC_AOI22_X1 T7192 ( .Y(T7192_Y), .B1(T7194_Y), .B0(T13586_Q),     .A1(T7233_Y), .A0(T9642_Y));
KC_AOI22_X1 T7146 ( .Y(T7146_Y), .B1(T14733_Q), .B0(T9576_Y),     .A1(T14730_Q), .A0(T15237_Y));
KC_AOI22_X1 T7141 ( .Y(T7141_Y), .B1(T7143_Y), .B0(T13597_Q),     .A1(T7236_Y), .A0(T4937_Y));
KC_AOI22_X1 T7139 ( .Y(T7139_Y), .B1(T7142_Y), .B0(T13575_Q),     .A1(T7036_Y), .A0(T9642_Y));
KC_AOI22_X1 T7113 ( .Y(T7113_Y), .B1(T15739_Y), .B0(T434_Q),     .A1(T8389_Y), .A0(T5240_Q));
KC_AOI22_X1 T7109 ( .Y(T7109_Y), .B1(T15734_Y), .B0(T813_Q),     .A1(T15735_Y), .A0(T825_Q));
KC_AOI22_X1 T5231 ( .Y(T5231_Y), .B1(T13651_Q), .B0(T9637_Y),     .A1(T13637_Q), .A0(T6483_Y));
KC_AOI22_X1 T5232 ( .Y(T5232_Y), .B1(T14789_Q), .B0(T12076_Y),     .A1(T13683_Q), .A0(T12074_Y));
KC_AOI22_X1 T5233 ( .Y(T5233_Y), .B1(T6452_Y), .B0(T14810_Q),     .A1(T1632_Y), .A0(T14811_Q));
KC_AOI22_X1 T5234 ( .Y(T5234_Y), .B1(T13672_Q), .B0(T9665_Y),     .A1(T13675_Q), .A0(T15256_Y));
KC_AOI22_X1 T10649 ( .Y(T10649_Y), .B1(T10419_Y), .B0(T13706_Q),     .A1(T1338_Y), .A0(T13702_Q));
KC_AOI22_X1 T7298 ( .Y(T7298_Y), .B1(T6818_Y), .B0(T677_Q),     .A1(T6828_Y), .A0(T860_Q));
KC_AOI22_X1 T7295 ( .Y(T7295_Y), .B1(T6597_Y), .B0(T679_Q),     .A1(T6829_Y), .A0(T5238_Q));
KC_AOI22_X1 T7272 ( .Y(T7272_Y), .B1(T15737_Y), .B0(T320_Q),     .A1(T15311_Y), .A0(T5252_Q));
KC_AOI22_X1 T7240 ( .Y(T7240_Y), .B1(T12423_Y), .B0(T4855_Q),     .A1(T12408_Y), .A0(T860_Q));
KC_AOI22_X1 T5656 ( .Y(T5656_Y), .B1(T10358_Y), .B0(T14743_Q),     .A1(T9712_Y), .A0(T14744_Q));
KC_AOI22_X1 T5655 ( .Y(T5655_Y), .B1(T9707_Y), .B0(T13693_Q),     .A1(T10347_Y), .A0(T13736_Q));
KC_AOI22_X1 T5247 ( .Y(T5247_Y), .B1(T14758_Q), .B0(T9635_Y),     .A1(T14756_Q), .A0(T5088_Y));
KC_AOI22_X1 T5248 ( .Y(T5248_Y), .B1(T9664_Y), .B0(T14758_Q),     .A1(T3610_Y), .A0(T14756_Q));
KC_AOI22_X1 T5249 ( .Y(T5249_Y), .B1(T3027_Y), .B0(T14762_Q),     .A1(T9636_Y), .A0(T14764_Q));
KC_AOI22_X1 T5250 ( .Y(T5250_Y), .B1(T9664_Y), .B0(T13647_Q),     .A1(T3610_Y), .A0(T13763_Q));
KC_AOI22_X1 T10832 ( .Y(T10832_Y), .B1(T14670_Q), .B0(T10422_Y),     .A1(T13842_Q), .A0(T10367_Y));
KC_AOI22_X1 T7520 ( .Y(T7520_Y), .B1(T10420_Y), .B0(T13830_Q),     .A1(T10423_Y), .A0(T13843_Q));
KC_AOI22_X1 T7473 ( .Y(T7473_Y), .B1(T13797_Q), .B0(T12327_Y),     .A1(T13868_Q), .A0(T10788_Y));
KC_AOI22_X1 T7453 ( .Y(T7453_Y), .B1(T15311_Y), .B0(T359_Q),     .A1(T15737_Y), .A0(T5304_Q));
KC_AOI22_X1 T7441 ( .Y(T7441_Y), .B1(T12423_Y), .B0(T698_Q),     .A1(T12408_Y), .A0(T4858_Q));
KC_AOI22_X1 T7424 ( .Y(T7424_Y), .B1(T15737_Y), .B0(T343_Q),     .A1(T15311_Y), .A0(T190_Q));
KC_AOI22_X1 T5808 ( .Y(T5808_Y), .B1(T10346_Y), .B0(T13887_Q),     .A1(T15245_Y), .A0(T13886_Q));
KC_AOI22_X1 T5266 ( .Y(T5266_Y), .B1(T9731_Y), .B0(T14048_Q),     .A1(T3640_Y), .A0(T14853_Q));
KC_AOI22_X1 T5267 ( .Y(T5267_Y), .B1(T14921_Q), .B0(T9864_Y),     .A1(T14911_Q), .A0(T9865_Y));
KC_AOI22_X1 T5269 ( .Y(T5269_Y), .B1(T9763_Y), .B0(T14833_Q),     .A1(T3623_Y), .A0(T14830_Q));
KC_AOI22_X1 T5271 ( .Y(T5271_Y), .B1(T14922_Q), .B0(T9763_Y),     .A1(T14926_Q), .A0(T3623_Y));
KC_AOI22_X1 T5272 ( .Y(T5272_Y), .B1(T5792_Y), .B0(T14857_Q),     .A1(T4231_Y), .A0(T14994_Y));
KC_AOI22_X1 T7792 ( .Y(T7792_Y), .B1(T7793_Y), .B0(T13946_Q),     .A1(T7738_Y), .A0(T1484_Y));
KC_AOI22_X1 T7762 ( .Y(T7762_Y), .B1(T7150_Y), .B0(T15220_Y),     .A1(T7777_Y), .A0(T12086_Y));
KC_AOI22_X1 T7648 ( .Y(T7648_Y), .B1(T7640_Y), .B0(T725_Q),     .A1(T7652_Y), .A0(T5348_Q));
KC_AOI22_X1 T7573 ( .Y(T7573_Y), .B1(T8752_Y), .B0(T9381_Y),     .A1(T7564_Y), .A0(T918_Y));
KC_AOI22_X1 T5286 ( .Y(T5286_Y), .B1(T9706_Y), .B0(T14071_Q),     .A1(T1545_Y), .A0(T14059_Q));
KC_AOI22_X1 T5287 ( .Y(T5287_Y), .B1(T3688_Y), .B0(T16165_Y),     .A1(T3011_Y), .A0(T2532_Y));
KC_AOI22_X1 T16350 ( .Y(T16350_Y), .B1(T5358_Y), .B0(T8764_Y),     .A1(T8756_Y), .A0(T786_Y));
KC_AOI22_X1 T10762 ( .Y(T10762_Y), .B1(T10652_Y), .B0(T14613_Q),     .A1(T7975_Y), .A0(T1484_Y));
KC_AOI22_X1 T8005 ( .Y(T8005_Y), .B1(T7953_Y), .B0(T14608_Q),     .A1(T9992_Y), .A0(T2565_Y));
KC_AOI22_X1 T7939 ( .Y(T7939_Y), .B1(T14107_Q), .B0(T9893_Y),     .A1(T14254_Q), .A0(T15229_Y));
KC_AOI22_X1 T7927 ( .Y(T7927_Y), .B1(T14101_Q), .B0(T1584_Y),     .A1(T14114_Q), .A0(T1585_Y));
KC_AOI22_X1 T7907 ( .Y(T7907_Y), .B1(T8867_Y), .B0(T8397_Y),     .A1(T11264_Y), .A0(T8868_Y));
KC_AOI22_X1 T7887 ( .Y(T7887_Y), .B1(T985_Y), .B0(T8855_Y),     .A1(T1151_Q), .A0(T723_Y));
KC_AOI22_X1 T5323 ( .Y(T5323_Y), .B1(T9862_Y), .B0(T14877_Q),     .A1(T9824_Y), .A0(T14179_Q));
KC_AOI22_X1 T5326 ( .Y(T5326_Y), .B1(T5887_Y), .B0(T14198_Q),     .A1(T3669_Y), .A0(T14994_Y));
KC_AOI22_X1 T5328 ( .Y(T5328_Y), .B1(T9823_Y), .B0(T14163_Q),     .A1(T9825_Y), .A0(T14162_Q));
KC_AOI22_X1 T5329 ( .Y(T5329_Y), .B1(T5865_Y), .B0(T14881_Q),     .A1(T3137_Y), .A0(T14994_Y));
KC_AOI22_X1 T5332 ( .Y(T5332_Y), .B1(T14877_Q), .B0(T9863_Y),     .A1(T14179_Q), .A0(T9868_Y));
KC_AOI22_X1 T10705 ( .Y(T10705_Y), .B1(T14265_Q), .B0(T9892_Y),     .A1(T14249_Q), .A0(T9902_Y));
KC_AOI22_X1 T10667 ( .Y(T10667_Y), .B1(T14219_Q), .B0(T1584_Y),     .A1(T14208_Q), .A0(T1585_Y));
KC_AOI22_X1 T10664 ( .Y(T10664_Y), .B1(T10306_Y), .B0(T14217_Q),     .A1(T10009_Y), .A0(T14218_Q));
KC_AOI22_X1 T8133 ( .Y(T8133_Y), .B1(T8964_Y), .B0(T9441_Y),     .A1(T8642_Y), .A0(T10069_Y));
KC_AOI22_X1 T8051 ( .Y(T8051_Y), .B1(T12886_Y), .B0(T8948_Y),     .A1(T1214_Y), .A0(T1213_Y));
KC_AOI22_X1 T5368 ( .Y(T5368_Y), .B1(T14317_Q), .B0(T16442_Y),     .A1(T14313_Q), .A0(T15254_Y));
KC_AOI22_X1 T4832 ( .Y(T4832_Y), .B1(T14375_Q), .B0(T12088_Y),     .A1(T14381_Q), .A0(T8011_Y));
KC_AOI22_X1 T4830 ( .Y(T4830_Y), .B1(T12094_Y), .B0(T14371_Q),     .A1(T8000_Y), .A0(T14590_Q));
KC_AOI22_X1 T1576 ( .Y(T1576_Y), .B1(T7859_Y), .B0(T9011_Y),     .A1(T772_Q), .A0(T9034_Y));
KC_AOI22_X1 T1575 ( .Y(T1575_Y), .B1(T7811_Y), .B0(T9011_Y),     .A1(T5416_Q), .A0(T9034_Y));
KC_AOI22_X1 T1558 ( .Y(T1558_Y), .B1(T1001_Q), .B0(T8996_Y),     .A1(T1000_Q), .A0(T9002_Y));
KC_AOI22_X1 T10734 ( .Y(T10734_Y), .B1(T12094_Y), .B0(T14376_Q),     .A1(T8000_Y), .A0(T14383_Q));
KC_AOI22_X1 T5399 ( .Y(T5399_Y), .B1(T14456_Q), .B0(T12088_Y),     .A1(T14455_Q), .A0(T8011_Y));
KC_AOI22_X1 T5400 ( .Y(T5400_Y), .B1(T12094_Y), .B0(T14593_Q),     .A1(T8000_Y), .A0(T14454_Q));
KC_AOI22_X1 T5401 ( .Y(T5401_Y), .B1(T10504_Y), .B0(T14447_Q),     .A1(T15215_Y), .A0(T14444_Q));
KC_AOI22_X1 T5402 ( .Y(T5402_Y), .B1(T10504_Y), .B0(T14909_Q),     .A1(T15215_Y), .A0(T14908_Q));
KC_AOI22_X1 T5403 ( .Y(T5403_Y), .B1(T10504_Y), .B0(T14432_Q),     .A1(T15215_Y), .A0(T14419_Q));
KC_AOI22_X1 T5445 ( .Y(T5445_Y), .B1(T3245_Q), .B0(T5141_Y),     .A1(T3877_Q), .A0(T11506_Y));
KC_AOI22_X1 T5447 ( .Y(T5447_Y), .B1(T3244_Q), .B0(T5141_Y),     .A1(T3883_Q), .A0(T11506_Y));
KC_AOI22_X1 T5470 ( .Y(T5470_Y), .B1(T3967_Y), .B0(T8329_Y),     .A1(T11451_Y), .A0(T11505_Y));
KC_AOI22_X1 T5489 ( .Y(T5489_Y), .B1(T2819_Y), .B0(T2281_Q),     .A1(T10593_Y), .A0(T8352_Q));
KC_AOI22_X1 T5493 ( .Y(T5493_Y), .B1(T1785_Q), .B0(T11728_Y),     .A1(T3785_Y), .A0(T12268_Y));
KC_AOI22_X1 T6466 ( .Y(T6466_Y), .B1(T5566_Q), .B0(T4965_Y),     .A1(T16023_Q), .A0(T2876_Y));
KC_AOI22_X1 T5505 ( .Y(T5505_Y), .B1(T1829_Q), .B0(T4965_Y),     .A1(T2809_Q), .A0(T2876_Y));
KC_AOI22_X1 T5506 ( .Y(T5506_Y), .B1(T5522_Y), .B0(T16102_Y),     .A1(T2859_Y), .A0(T6182_Y));
KC_AOI22_X1 T5507 ( .Y(T5507_Y), .B1(T10974_Y), .B0(T6842_S),     .A1(T6610_S), .A0(T10568_Y));
KC_AOI22_X1 T5514 ( .Y(T5514_Y), .B1(T12061_Y), .B0(T6240_Y),     .A1(T11812_Y), .A0(T16270_Y));
KC_AOI22_X1 T5519 ( .Y(T5519_Y), .B1(T16050_Y), .B0(T10571_Y),     .A1(T10542_Y), .A0(T16102_Y));
KC_AOI22_X1 T5534 ( .Y(T5534_Y), .B1(T8431_Y), .B0(T11817_Y),     .A1(T10593_Y), .A0(T6614_S));
KC_AOI22_X1 T16348 ( .Y(T16348_Y), .B1(T8764_Y), .B0(T8772_Y),     .A1(T9365_Y), .A0(T786_Y));
KC_AOI22_X1 T16336 ( .Y(T16336_Y), .B1(T12607_Y), .B0(T9375_Y),     .A1(T16333_Y), .A0(T16332_Y));
KC_AOI22_X1 T16280 ( .Y(T16280_Y), .B1(T1006_Y), .B0(T8996_Y),     .A1(T5384_Q), .A0(T9002_Y));
KC_AOI22_X1 T6685 ( .Y(T6685_Y), .B1(T9503_Y), .B0(T715_Y),     .A1(T10344_Y), .A0(T15223_Y));
KC_AOI22_X1 T10830 ( .Y(T10830_Y), .B1(T14672_Q), .B0(T10422_Y),     .A1(T14673_Q), .A0(T10367_Y));
KC_AOI22_X1 T10817 ( .Y(T10817_Y), .B1(T7035_Y), .B0(T15220_Y),     .A1(T5679_Y), .A0(T12086_Y));
KC_AOI22_X1 T10804 ( .Y(T10804_Y), .B1(T9704_Y), .B0(T14743_Q),     .A1(T9705_Y), .A0(T14744_Q));
KC_AOI22_X1 T10795 ( .Y(T10795_Y), .B1(T10419_Y), .B0(T14003_Q),     .A1(T1338_Y), .A0(T14006_Q));
KC_AOI22_X1 T5550 ( .Y(T5550_Y), .B1(T6673_Y), .B0(T14069_Q),     .A1(T3614_Y), .A0(T14994_Y));
KC_AOI22_X1 T5551 ( .Y(T5551_Y), .B1(T9823_Y), .B0(T14825_Q),     .A1(T9825_Y), .A0(T14824_Q));
KC_AOI22_X1 T5552 ( .Y(T5552_Y), .B1(T14781_Q), .B0(T3611_Y),     .A1(T14780_Q), .A0(T6482_Y));
KC_AOI22_X1 T5554 ( .Y(T5554_Y), .B1(T5568_Q), .B0(T6352_Y),     .A1(T12833_Y), .A0(T2073_Y));
KC_AOI22_X1 T5555 ( .Y(T5555_Y), .B1(T8296_Y), .B0(T11613_Y),     .A1(T11999_Y), .A0(T8503_Y));
KC_NAND2_X2 T5637 ( .B(T5190_Q), .A(T5589_Q), .Y(T5637_Y));
KC_NAND2_X2 T5624 ( .B(T878_Y), .A(T15213_Y), .Y(T5624_Y));
KC_NAND2_X2 T5607 ( .B(T5606_Y), .A(T40_Y), .Y(T5607_Y));
KC_NAND2_X2 T5619 ( .B(T103_Q), .A(T15319_Y), .Y(T5619_Y));
KC_NAND2_X2 T5618 ( .B(T12369_Y), .A(T12371_Y), .Y(T5618_Y));
KC_NAND2_X2 T5605 ( .B(T106_Q), .A(T5202_Q), .Y(T5605_Y));
KC_NAND2_X2 T5596 ( .B(T15315_Y), .A(T106_Q), .Y(T5596_Y));
KC_NAND2_X2 T6862 ( .B(T16310_Y), .A(T1201_Y), .Y(T6862_Y));
KC_NAND2_X2 T5604 ( .B(T16479_Y), .A(T8559_Y), .Y(T5604_Y));
KC_NAND2_X2 T6934 ( .B(T150_Q), .A(T5222_Q), .Y(T6934_Y));
KC_NAND2_X2 T6914 ( .B(T11262_Y), .A(T228_Y), .Y(T6914_Y));
KC_NAND2_X2 T9272 ( .B(T257_Y), .A(T6319_Y), .Y(T9272_Y));
KC_NAND2_X2 T7122 ( .B(T16176_Y), .A(T13229_Q), .Y(T7122_Y));
KC_NAND2_X2 T7698 ( .B(T7583_Y), .A(T8747_Y), .Y(T7698_Y));
KC_NAND2_X2 T7682 ( .B(T8746_Y), .A(T7845_Y), .Y(T7682_Y));
KC_NAND2_X2 T7680 ( .B(T7581_Y), .A(T208_Q), .Y(T7680_Y));
KC_NAND2_X2 T7678 ( .B(T743_Y), .A(T7580_Y), .Y(T7678_Y));
KC_NAND2_X2 T7584 ( .B(T8746_Y), .A(T16176_Y), .Y(T7584_Y));
KC_NAND2_X2 T9397 ( .B(T12383_Y), .A(T15656_Y), .Y(T9397_Y));
KC_NAND2_X2 T9030 ( .B(T243_Y), .A(T9013_Y), .Y(T9030_Y));
KC_NAND2_X2 T8992 ( .B(T8993_S), .A(T8960_Y), .Y(T8992_Y));
KC_NAND2_X2 T8991 ( .B(T8994_Y), .A(T1364_Y), .Y(T8991_Y));
KC_NAND2_X2 T9181 ( .B(T15118_Y), .A(T15100_Y), .Y(T9181_Y));
KC_NAND2_X2 T9158 ( .B(T4800_Y), .A(T9180_Y), .Y(T9158_Y));
KC_NAND2_X2 T9092 ( .B(T9087_Y), .A(T15150_Y), .Y(T9092_Y));
KC_NAND2_X2 T9091 ( .B(T15100_Y), .A(T4818_Y), .Y(T9091_Y));
KC_NAND2_X2 T9267 ( .B(T265_Y), .A(T288_Q), .Y(T9267_Y));
KC_NAND2_X2 T9266 ( .B(T1477_Y), .A(T9267_Y), .Y(T9266_Y));
KC_NAND2_X2 T9261 ( .B(T332_Y), .A(T306_Q), .Y(T9261_Y));
KC_NAND2_X2 T7121 ( .B(T6368_Y), .A(T7087_Y), .Y(T7121_Y));
KC_NAND2_X2 T7120 ( .B(T318_Y), .A(T313_Q), .Y(T7120_Y));
KC_NAND2_X2 T7105 ( .B(T321_Y), .A(T275_Q), .Y(T7105_Y));
KC_NAND2_X2 T7104 ( .B(T6612_Y), .A(T7105_Y), .Y(T7104_Y));
KC_NAND2_X2 T7087 ( .B(T348_Y), .A(T158_Q), .Y(T7087_Y));
KC_NAND2_X2 T7084 ( .B(T6377_Y), .A(T7120_Y), .Y(T7084_Y));
KC_NAND2_X2 T9260 ( .B(T6607_Y), .A(T9261_Y), .Y(T9260_Y));
KC_NAND2_X2 T7679 ( .B(T7628_Y), .A(T739_Y), .Y(T7679_Y));
KC_NAND2_X2 T7670 ( .B(T7819_Y), .A(T7662_Y), .Y(T7670_Y));
KC_NAND2_X2 T7669 ( .B(T7626_Y), .A(T7823_Y), .Y(T7669_Y));
KC_NAND2_X2 T7627 ( .B(T8679_Y), .A(T350_Y), .Y(T7627_Y));
KC_NAND2_X2 T7626 ( .B(T8654_Y), .A(T350_Y), .Y(T7626_Y));
KC_NAND2_X2 T7579 ( .B(T7826_Y), .A(T7570_Y), .Y(T7579_Y));
KC_NAND2_X2 T7578 ( .B(T7661_Y), .A(T7821_Y), .Y(T7578_Y));
KC_NAND2_X2 T7577 ( .B(T7578_Y), .A(T739_Y), .Y(T7577_Y));
KC_NAND2_X2 T9398 ( .B(T7677_Y), .A(T6944_Y), .Y(T9398_Y));
KC_NAND2_X2 T9387 ( .B(T9386_Y), .A(T9388_Y), .Y(T9387_Y));
KC_NAND2_X2 T9386 ( .B(T612_Y), .A(T8775_Y), .Y(T9386_Y));
KC_NAND2_X2 T7918 ( .B(T8140_Y), .A(T7817_Y), .Y(T7918_Y));
KC_NAND2_X2 T7917 ( .B(T1213_Y), .A(T350_Y), .Y(T7917_Y));
KC_NAND2_X2 T7916 ( .B(T8080_Y), .A(T7917_Y), .Y(T7916_Y));
KC_NAND2_X2 T7911 ( .B(T8665_Y), .A(T371_Y), .Y(T7911_Y));
KC_NAND2_X2 T7910 ( .B(T7818_Y), .A(T8139_Y), .Y(T7910_Y));
KC_NAND2_X2 T7863 ( .B(T7860_Y), .A(T8138_Y), .Y(T7863_Y));
KC_NAND2_X2 T7860 ( .B(T8610_Y), .A(T350_Y), .Y(T7860_Y));
KC_NAND2_X2 T7833 ( .B(T5354_Q), .A(T235_Q), .Y(T7833_Y));
KC_NAND2_X2 T7832 ( .B(T924_Y), .A(T7828_Y), .Y(T7832_Y));
KC_NAND2_X2 T7831 ( .B(T235_Q), .A(T921_Y), .Y(T7831_Y));
KC_NAND2_X2 T7830 ( .B(T8143_Y), .A(T8777_Y), .Y(T7830_Y));
KC_NAND2_X2 T7828 ( .B(T8775_Y), .A(T920_Y), .Y(T7828_Y));
KC_NAND2_X2 T7825 ( .B(T16514_Y), .A(T920_Y), .Y(T7825_Y));
KC_NAND2_X2 T7824 ( .B(T9386_Y), .A(T7827_Y), .Y(T7824_Y));
KC_NAND2_X2 T7823 ( .B(T9116_Y), .A(T8777_Y), .Y(T7823_Y));
KC_NAND2_X2 T7822 ( .B(T7826_Y), .A(T7828_Y), .Y(T7822_Y));
KC_NAND2_X2 T7821 ( .B(T8964_Y), .A(T8777_Y), .Y(T7821_Y));
KC_NAND2_X2 T7819 ( .B(T9067_Y), .A(T8777_Y), .Y(T7819_Y));
KC_NAND2_X2 T7818 ( .B(T8625_Y), .A(T350_Y), .Y(T7818_Y));
KC_NAND2_X2 T7817 ( .B(T9325_Y), .A(T350_Y), .Y(T7817_Y));
KC_NAND2_X2 T9014 ( .B(T9029_Y), .A(T9013_Y), .Y(T9014_Y));
KC_NAND2_X2 T8149 ( .B(T9449_Y), .A(T1429_Y), .Y(T8149_Y));
KC_NAND2_X2 T8148 ( .B(T9068_Y), .A(T8865_Y), .Y(T8148_Y));
KC_NAND2_X2 T8147 ( .B(T9449_Y), .A(T1439_Y), .Y(T8147_Y));
KC_NAND2_X2 T8146 ( .B(T9449_Y), .A(T9071_Y), .Y(T8146_Y));
KC_NAND2_X2 T8145 ( .B(T16286_Y), .A(T9021_Y), .Y(T8145_Y));
KC_NAND2_X2 T8144 ( .B(T16286_Y), .A(T9027_Y), .Y(T8144_Y));
KC_NAND2_X2 T8140 ( .B(T9058_Y), .A(T8865_Y), .Y(T8140_Y));
KC_NAND2_X2 T8139 ( .B(T233_Y), .A(T8865_Y), .Y(T8139_Y));
KC_NAND2_X2 T8138 ( .B(T8871_Y), .A(T8865_Y), .Y(T8138_Y));
KC_NAND2_X2 T8137 ( .B(T6800_Y), .A(T8865_Y), .Y(T8137_Y));
KC_NAND2_X2 T8109 ( .B(T393_Y), .A(T15488_Y), .Y(T8109_Y));
KC_NAND2_X2 T8104 ( .B(T613_Y), .A(T8962_Y), .Y(T8104_Y));
KC_NAND2_X2 T8103 ( .B(T8962_Y), .A(T1330_Y), .Y(T8103_Y));
KC_NAND2_X2 T8102 ( .B(T8079_Y), .A(T7857_Y), .Y(T8102_Y));
KC_NAND2_X2 T8100 ( .B(T16513_Y), .A(T1330_Y), .Y(T8100_Y));
KC_NAND2_X2 T8099 ( .B(T8104_Y), .A(T8078_Y), .Y(T8099_Y));
KC_NAND2_X2 T8083 ( .B(T7858_Y), .A(T1284_Y), .Y(T8083_Y));
KC_NAND2_X2 T8082 ( .B(T8104_Y), .A(T7917_Y), .Y(T8082_Y));
KC_NAND2_X2 T8081 ( .B(T1206_Y), .A(T8103_Y), .Y(T8081_Y));
KC_NAND2_X2 T8080 ( .B(T8079_Y), .A(T8103_Y), .Y(T8080_Y));
KC_NAND2_X2 T8078 ( .B(T8963_Y), .A(T1330_Y), .Y(T8078_Y));
KC_NAND2_X2 T8077 ( .B(T1273_Y), .A(T8079_Y), .Y(T8077_Y));
KC_NAND2_X2 T8053 ( .B(T7863_Y), .A(T1284_Y), .Y(T8053_Y));
KC_NAND2_X2 T9174 ( .B(T9137_Y), .A(T9117_Y), .Y(T9174_Y));
KC_NAND2_X2 T9173 ( .B(T16286_Y), .A(T9170_Y), .Y(T9173_Y));
KC_NAND2_X2 T9172 ( .B(T16286_Y), .A(T9171_Y), .Y(T9172_Y));
KC_NAND2_X2 T9152 ( .B(T9169_Y), .A(T9121_Y), .Y(T9152_Y));
KC_NAND2_X2 T9151 ( .B(T9168_Y), .A(T9121_Y), .Y(T9151_Y));
KC_NAND2_X2 T9129 ( .B(T9120_Y), .A(T9072_Y), .Y(T9129_Y));
KC_NAND2_X2 T9128 ( .B(T9118_Y), .A(T9069_Y), .Y(T9128_Y));
KC_NAND2_X2 T9127 ( .B(T9120_Y), .A(T9069_Y), .Y(T9127_Y));
KC_NAND2_X2 T9126 ( .B(T4801_Y), .A(T9123_Y), .Y(T9126_Y));
KC_NAND2_X2 T9125 ( .B(T16286_Y), .A(T9136_Y), .Y(T9125_Y));
KC_NAND2_X2 T9093 ( .B(T9137_Y), .A(T9072_Y), .Y(T9093_Y));
KC_NAND2_X2 T9079 ( .B(T9137_Y), .A(T9069_Y), .Y(T9079_Y));
KC_NAND2_X2 T9078 ( .B(T9120_Y), .A(T9117_Y), .Y(T9078_Y));
KC_NAND2_X2 T9077 ( .B(T9118_Y), .A(T9072_Y), .Y(T9077_Y));
KC_NAND2_X2 T7097 ( .B(T6375_Y), .A(T7082_Y), .Y(T7097_Y));
KC_NAND2_X2 T7082 ( .B(T347_Y), .A(T460_Q), .Y(T7082_Y));
KC_NAND2_X2 T7307 ( .B(T6348_Y), .A(T5265_Q), .Y(T7307_Y));
KC_NAND2_X2 T7306 ( .B(T6618_Y), .A(T7307_Y), .Y(T7306_Y));
KC_NAND2_X2 T7250 ( .B(T6346_Y), .A(T4835_Q), .Y(T7250_Y));
KC_NAND2_X2 T7249 ( .B(T6366_Y), .A(T7250_Y), .Y(T7249_Y));
KC_NAND2_X2 T7662 ( .B(T9321_Y), .A(T382_Y), .Y(T7662_Y));
KC_NAND2_X2 T7661 ( .B(T8632_Y), .A(T382_Y), .Y(T7661_Y));
KC_NAND2_X2 T7901 ( .B(T8072_Y), .A(T16388_Y), .Y(T7901_Y));
KC_NAND2_X2 T7900 ( .B(T16388_Y), .A(T16420_Y), .Y(T7900_Y));
KC_NAND2_X2 T7827 ( .B(T8776_Y), .A(T920_Y), .Y(T7827_Y));
KC_NAND2_X2 T7816 ( .B(T612_Y), .A(T16514_Y), .Y(T7816_Y));
KC_NAND2_X2 T9015 ( .B(T9053_S), .A(T1421_Y), .Y(T9015_Y));
KC_NAND2_X2 T8131 ( .B(T9019_Y), .A(T9442_Y), .Y(T8131_Y));
KC_NAND2_X2 T8130 ( .B(T1328_Y), .A(T8981_Y), .Y(T8130_Y));
KC_NAND2_X2 T8129 ( .B(T233_Y), .A(T9442_Y), .Y(T8129_Y));
KC_NAND2_X2 T8128 ( .B(T8120_Y), .A(T8980_Y), .Y(T8128_Y));
KC_NAND2_X2 T8127 ( .B(T559_Y), .A(T8864_Y), .Y(T8127_Y));
KC_NAND2_X2 T8126 ( .B(T9148_Y), .A(T9442_Y), .Y(T8126_Y));
KC_NAND2_X2 T8125 ( .B(T8983_Y), .A(T7829_Y), .Y(T8125_Y));
KC_NAND2_X2 T8119 ( .B(T8116_Y), .A(T750_Q), .Y(T8119_Y));
KC_NAND2_X2 T8101 ( .B(T613_Y), .A(T16513_Y), .Y(T8101_Y));
KC_NAND2_X2 T8073 ( .B(T1323_Y), .A(T566_Q), .Y(T8073_Y));
KC_NAND2_X2 T8065 ( .B(T1323_Y), .A(T5378_Q), .Y(T8065_Y));
KC_NAND2_X2 T8046 ( .B(T8041_Y), .A(T1205_Y), .Y(T8046_Y));
KC_NAND2_X2 T8038 ( .B(T9007_Y), .A(T16310_Y), .Y(T8038_Y));
KC_NAND2_X2 T9113 ( .B(T9109_Y), .A(T606_Q), .Y(T9113_Y));
KC_NAND2_X2 T9112 ( .B(T9107_Y), .A(T5406_Q), .Y(T9112_Y));
KC_NAND2_X2 T9065 ( .B(T567_Q), .A(T561_Q), .Y(T9065_Y));
KC_NAND2_X2 T6919 ( .B(T453_Q), .A(T310_Y), .Y(T6919_Y));
KC_NAND2_X2 T1143 ( .B(T8636_Y), .A(T8633_Y), .Y(T1143_Y));
KC_NAND2_X2 T9319 ( .B(T7599_Y), .A(T8762_Y), .Y(T9319_Y));
KC_NAND2_X2 T7684 ( .B(T7847_Y), .A(T931_Y), .Y(T7684_Y));
KC_NAND2_X2 T7646 ( .B(T907_Y), .A(T12417_Y), .Y(T7646_Y));
KC_NAND2_X2 T7645 ( .B(T907_Y), .A(T12414_Y), .Y(T7645_Y));
KC_NAND2_X2 T7644 ( .B(T907_Y), .A(T12415_Y), .Y(T7644_Y));
KC_NAND2_X2 T7563 ( .B(T907_Y), .A(T12416_Y), .Y(T7563_Y));
KC_NAND2_X2 T9420 ( .B(T8736_Y), .A(T9416_Y), .Y(T9420_Y));
KC_NAND2_X2 T7847 ( .B(T1095_Q), .A(T8794_Y), .Y(T7847_Y));
KC_NAND2_X2 T7846 ( .B(T928_Y), .A(T7582_Y), .Y(T7846_Y));
KC_NAND2_X2 T9009 ( .B(T747_Q), .A(T9433_Y), .Y(T9009_Y));
KC_NAND2_X2 T9007 ( .B(T4843_Q), .A(T977_Q), .Y(T9007_Y));
KC_NAND2_X2 T8121 ( .B(T9018_Y), .A(T9442_Y), .Y(T8121_Y));
KC_NAND2_X2 T8120 ( .B(T8978_Y), .A(T8977_Y), .Y(T8120_Y));
KC_NAND2_X2 T8117 ( .B(T5379_Q), .A(T977_Q), .Y(T8117_Y));
KC_NAND2_X2 T8116 ( .B(T5383_Q), .A(T977_Q), .Y(T8116_Y));
KC_NAND2_X2 T8067 ( .B(T8946_Y), .A(T977_Q), .Y(T8067_Y));
KC_NAND2_X2 T8066 ( .B(T8117_Y), .A(T1255_Y), .Y(T8066_Y));
KC_NAND2_X2 T8064 ( .B(T1327_Y), .A(T8941_Y), .Y(T8064_Y));
KC_NAND2_X2 T8063 ( .B(T1255_Y), .A(T1198_Y), .Y(T8063_Y));
KC_NAND2_X2 T9444 ( .B(T9459_Q), .A(T9002_Y), .Y(T9444_Y));
KC_NAND2_X2 T9161 ( .B(T11268_Y), .A(T8901_Y), .Y(T9161_Y));
KC_NAND2_X2 T9052 ( .B(T8397_Y), .A(T9442_Y), .Y(T9052_Y));
KC_NAND2_X2 T9051 ( .B(T9068_Y), .A(T9442_Y), .Y(T9051_Y));
KC_NAND2_X2 T9050 ( .B(T9058_Y), .A(T9442_Y), .Y(T9050_Y));
KC_NAND2_X2 T9043 ( .B(T1005_Q), .A(T9002_Y), .Y(T9043_Y));
KC_NAND2_X2 T9042 ( .B(T1152_Q), .A(T9002_Y), .Y(T9042_Y));
KC_NAND2_X2 T9041 ( .B(T1154_Q), .A(T9002_Y), .Y(T9041_Y));
KC_NAND2_X2 T9318 ( .B(T7599_Y), .A(T8762_Y), .Y(T9318_Y));
KC_NAND2_X2 T9316 ( .B(T7599_Y), .A(T8758_Y), .Y(T9316_Y));
KC_NAND2_X2 T9308 ( .B(T8707_Y), .A(T6694_Y), .Y(T9308_Y));
KC_NAND2_X2 T9306 ( .B(T8670_Y), .A(T6694_Y), .Y(T9306_Y));
KC_NAND2_X2 T7418 ( .B(T9370_Y), .A(T7839_Y), .Y(T7418_Y));
KC_NAND2_X2 T7414 ( .B(T497_Y), .A(T7555_Y), .Y(T7414_Y));
KC_NAND2_X2 T7413 ( .B(T549_Y), .A(T7555_Y), .Y(T7413_Y));
KC_NAND2_X2 T7412 ( .B(T6691_Y), .A(T7555_Y), .Y(T7412_Y));
KC_NAND2_X2 T7410 ( .B(T9370_Y), .A(T7555_Y), .Y(T7410_Y));
KC_NAND2_X2 T7637 ( .B(T1724_Y), .A(T15431_Y), .Y(T7637_Y));
KC_NAND2_X2 T7635 ( .B(T638_Y), .A(T5308_Q), .Y(T7635_Y));
KC_NAND2_X2 T7618 ( .B(T727_Y), .A(T8682_Y), .Y(T7618_Y));
KC_NAND2_X2 T7617 ( .B(T8715_Y), .A(T6694_Y), .Y(T7617_Y));
KC_NAND2_X2 T7616 ( .B(T9374_Y), .A(T8670_Y), .Y(T7616_Y));
KC_NAND2_X2 T7614 ( .B(T6694_Y), .A(T9370_Y), .Y(T7614_Y));
KC_NAND2_X2 T7599 ( .B(T886_Y), .A(T9361_Y), .Y(T7599_Y));
KC_NAND2_X2 T7593 ( .B(T9373_Y), .A(T8670_Y), .Y(T7593_Y));
KC_NAND2_X2 T7592 ( .B(T15223_Y), .A(T1131_Q), .Y(T7592_Y));
KC_NAND2_X2 T7591 ( .B(T9374_Y), .A(T8682_Y), .Y(T7591_Y));
KC_NAND2_X2 T7590 ( .B(T9373_Y), .A(T8682_Y), .Y(T7590_Y));
KC_NAND2_X2 T7557 ( .B(T15454_Y), .A(T10942_Y), .Y(T7557_Y));
KC_NAND2_X2 T9406 ( .B(T15457_Y), .A(T992_Q), .Y(T9406_Y));
KC_NAND2_X2 T9369 ( .B(T4872_Y), .A(T8828_Y), .Y(T9369_Y));
KC_NAND2_X2 T7881 ( .B(T948_Y), .A(T8846_Y), .Y(T7881_Y));
KC_NAND2_X2 T7870 ( .B(T958_Y), .A(T131_Q), .Y(T7870_Y));
KC_NAND2_X2 T7869 ( .B(T988_Y), .A(T8827_Y), .Y(T7869_Y));
KC_NAND2_X2 T7868 ( .B(T10880_Y), .A(T16275_Y), .Y(T7868_Y));
KC_NAND2_X2 T7867 ( .B(T16274_Y), .A(T16275_Y), .Y(T7867_Y));
KC_NAND2_X2 T7848 ( .B(T783_Y), .A(T8794_Y), .Y(T7848_Y));
KC_NAND2_X2 T7844 ( .B(T8791_Y), .A(T8796_Y), .Y(T7844_Y));
KC_NAND2_X2 T7842 ( .B(T8792_Y), .A(T16159_Y), .Y(T7842_Y));
KC_NAND2_X2 T7841 ( .B(T947_Y), .A(T8795_Y), .Y(T7841_Y));
KC_NAND2_X2 T7802 ( .B(T8831_Y), .A(T8828_Y), .Y(T7802_Y));
KC_NAND2_X2 T7801 ( .B(T8827_Y), .A(T15999_Y), .Y(T7801_Y));
KC_NAND2_X2 T9000 ( .B(T961_Y), .A(T972_Y), .Y(T9000_Y));
KC_NAND2_X2 T8999 ( .B(T4862_Q), .A(T9002_Y), .Y(T8999_Y));
KC_NAND2_X2 T8112 ( .B(T972_Y), .A(T16440_Y), .Y(T8112_Y));
KC_NAND2_X2 T8093 ( .B(T972_Y), .A(T1724_Y), .Y(T8093_Y));
KC_NAND2_X2 T9045 ( .B(T996_Q), .A(T9002_Y), .Y(T9045_Y));
KC_NAND2_X2 T9044 ( .B(T9458_Q), .A(T9002_Y), .Y(T9044_Y));
KC_NAND2_X2 T9508 ( .B(T9301_Y), .A(T6694_Y), .Y(T9508_Y));
KC_NAND2_X2 T9309 ( .B(T6826_Y), .A(T6694_Y), .Y(T9309_Y));
KC_NAND2_X2 T9307 ( .B(T9303_Y), .A(T6694_Y), .Y(T9307_Y));
KC_NAND2_X2 T7551 ( .B(T1044_Q), .A(T596_Y), .Y(T7551_Y));
KC_NAND2_X2 T7411 ( .B(T585_Y), .A(T7357_Y), .Y(T7411_Y));
KC_NAND2_X2 T7799 ( .B(T7845_Y), .A(T7623_Y), .Y(T7799_Y));
KC_NAND2_X2 T7741 ( .B(T7636_Y), .A(T1113_Q), .Y(T7741_Y));
KC_NAND2_X2 T7719 ( .B(T7636_Y), .A(T1128_Q), .Y(T7719_Y));
KC_NAND2_X2 T7638 ( .B(T7636_Y), .A(T1094_Q), .Y(T7638_Y));
KC_NAND2_X2 T7615 ( .B(T636_Y), .A(T9505_Y), .Y(T7615_Y));
KC_NAND2_X2 T7558 ( .B(T7636_Y), .A(T5334_Q), .Y(T7558_Y));
KC_NAND2_X2 T10331 ( .B(T7845_Y), .A(T15031_Y), .Y(T10331_Y));
KC_NAND2_X2 T10329 ( .B(T7845_Y), .A(T15839_Y), .Y(T10329_Y));
KC_NAND2_X2 T10328 ( .B(T7845_Y), .A(T15840_Y), .Y(T10328_Y));
KC_NAND2_X2 T10317 ( .B(T7999_Y), .A(T12095_Y), .Y(T10317_Y));
KC_NAND2_X2 T10316 ( .B(T12095_Y), .A(T15800_Y), .Y(T10316_Y));
KC_NAND2_X2 T8029 ( .B(T15664_Y), .A(T9891_Y), .Y(T8029_Y));
KC_NAND2_X2 T7999 ( .B(T7834_Y), .A(T8783_Y), .Y(T7999_Y));
KC_NAND2_X2 T7998 ( .B(T7834_Y), .A(T8781_Y), .Y(T7998_Y));
KC_NAND2_X2 T7997 ( .B(T7834_Y), .A(T15461_Y), .Y(T7997_Y));
KC_NAND2_X2 T7977 ( .B(T7834_Y), .A(T1050_Y), .Y(T7977_Y));
KC_NAND2_X2 T7976 ( .B(T10048_Y), .A(T1131_Q), .Y(T7976_Y));
KC_NAND2_X2 T7843 ( .B(T15664_Y), .A(T1095_Q), .Y(T7843_Y));
KC_NAND2_X2 T7840 ( .B(T16384_Y), .A(T9891_Y), .Y(T7840_Y));
KC_NAND2_X2 T10047 ( .B(T7977_Y), .A(T12095_Y), .Y(T10047_Y));
KC_NAND2_X2 T10046 ( .B(T8032_Y), .A(T5376_Q), .Y(T10046_Y));
KC_NAND2_X2 T10045 ( .B(T1249_Q), .A(T8032_Y), .Y(T10045_Y));
KC_NAND2_X2 T10044 ( .B(T12095_Y), .A(T8975_Y), .Y(T10044_Y));
KC_NAND2_X2 T10043 ( .B(T7998_Y), .A(T12095_Y), .Y(T10043_Y));
KC_NAND2_X2 T10026 ( .B(T7997_Y), .A(T12095_Y), .Y(T10026_Y));
KC_NAND2_X2 T10008 ( .B(T16149_Y), .A(T10000_Y), .Y(T10008_Y));
KC_NAND2_X2 T9987 ( .B(T10161_Y), .A(T10942_Y), .Y(T9987_Y));
KC_NAND2_X2 T8111 ( .B(T1341_Y), .A(T1196_Y), .Y(T8111_Y));
KC_NAND2_X2 T8110 ( .B(T1346_Y), .A(T10027_Y), .Y(T8110_Y));
KC_NAND2_X2 T8057 ( .B(T15487_Y), .A(T10008_Y), .Y(T8057_Y));
KC_NAND2_X2 T10175 ( .B(T1013_Q), .A(T977_Q), .Y(T10175_Y));
KC_NAND2_X2 T8025 ( .B(T16377_Y), .A(T7845_Y), .Y(T8025_Y));
KC_NAND2_X2 T10174 ( .B(T972_Y), .A(T10172_Y), .Y(T10174_Y));
KC_NAND2_X2 T10173 ( .B(T10175_Y), .A(T15999_Y), .Y(T10173_Y));
KC_NAND2_X2 T10159 ( .B(T1257_Y), .A(T10130_Y), .Y(T10159_Y));
KC_NAND2_X2 T10144 ( .B(T13125_Y), .A(T10934_Y), .Y(T10144_Y));
KC_NAND2_X2 T10143 ( .B(T972_Y), .A(T5814_Y), .Y(T10143_Y));
KC_NAND2_X2 T10142 ( .B(T2717_Y), .A(T5814_Y), .Y(T10142_Y));
KC_NAND2_X2 T10131 ( .B(T4831_Y), .A(T972_Y), .Y(T10131_Y));
KC_NAND2_X2 T10404 ( .B(T1633_Y), .A(T6595_Y), .Y(T10404_Y));
KC_NAND2_X2 T7182 ( .B(T361_Y), .A(T2589_Y), .Y(T7182_Y));
KC_NAND2_X2 T7351 ( .B(T403_Y), .A(T5331_Y), .Y(T7351_Y));
KC_NAND2_X2 T7350 ( .B(T6802_Y), .A(T6839_Y), .Y(T7350_Y));
KC_NAND2_X2 T7340 ( .B(T6802_Y), .A(T6839_Y), .Y(T7340_Y));
KC_NAND2_X2 T7339 ( .B(T403_Y), .A(T5331_Y), .Y(T7339_Y));
KC_NAND2_X2 T5674 ( .B(T6747_Y), .A(T2589_Y), .Y(T5674_Y));
KC_NAND2_X2 T5673 ( .B(T1633_Y), .A(T6595_Y), .Y(T5673_Y));
KC_NAND2_X2 T1357 ( .B(T1363_Y), .A(T1738_Y), .Y(T1357_Y));
KC_NAND2_X2 T10380 ( .B(T4884_Y), .A(T16448_Y), .Y(T10380_Y));
KC_NAND2_X2 T10389 ( .B(T10388_Y), .A(T12083_Y), .Y(T10389_Y));
KC_NAND2_X2 T6993 ( .B(T9539_Y), .A(T12081_Y), .Y(T6993_Y));
KC_NAND2_X2 T6992 ( .B(T12083_Y), .A(T10388_Y), .Y(T6992_Y));
KC_NAND2_X2 T6991 ( .B(T15393_Y), .A(T4884_Y), .Y(T6991_Y));
KC_NAND2_X2 T6990 ( .B(T15670_Y), .A(T4884_Y), .Y(T6990_Y));
KC_NAND2_X2 T6983 ( .B(T12081_Y), .A(T9539_Y), .Y(T6983_Y));
KC_NAND2_X2 T6982 ( .B(T4884_Y), .A(T16448_Y), .Y(T6982_Y));
KC_NAND2_X2 T7541 ( .B(T9719_Y), .A(T2534_Y), .Y(T7541_Y));
KC_NAND2_X2 T7489 ( .B(T2534_Y), .A(T9719_Y), .Y(T7489_Y));
KC_NAND2_X2 T10322 ( .B(T7990_Y), .A(T1586_Y), .Y(T10322_Y));
KC_NAND2_X2 T10018 ( .B(T10013_Y), .A(T9889_Y), .Y(T10018_Y));
KC_NAND2_X2 T10017 ( .B(T9889_Y), .A(T10013_Y), .Y(T10017_Y));
KC_NAND2_X2 T10016 ( .B(T15393_Y), .A(T1476_Y), .Y(T10016_Y));
KC_NAND2_X2 T9995 ( .B(T1476_Y), .A(T7703_Y), .Y(T9995_Y));
KC_NAND2_X2 T6890 ( .B(T6894_Y), .A(T6889_Y), .Y(T6890_Y));
KC_NAND2_X2 T7334 ( .B(T2451_Y), .A(T2589_Y), .Y(T7334_Y));
KC_NAND2_X2 T7320 ( .B(T403_Y), .A(T5331_Y), .Y(T7320_Y));
KC_NAND2_X2 T5664 ( .B(T6802_Y), .A(T6839_Y), .Y(T5664_Y));
KC_NAND2_X2 T5663 ( .B(T403_Y), .A(T5331_Y), .Y(T5663_Y));
KC_NAND2_X2 T5651 ( .B(T1633_Y), .A(T6595_Y), .Y(T5651_Y));
KC_NAND2_X2 T5650 ( .B(T2451_Y), .A(T2589_Y), .Y(T5650_Y));
KC_NAND2_X2 T5648 ( .B(T6802_Y), .A(T6839_Y), .Y(T5648_Y));
KC_NAND2_X2 T7782 ( .B(T7707_Y), .A(T7703_Y), .Y(T7782_Y));
KC_NAND2_X2 T7781 ( .B(T9809_Y), .A(T12328_Y), .Y(T7781_Y));
KC_NAND2_X2 T7705 ( .B(T15393_Y), .A(T7707_Y), .Y(T7705_Y));
KC_NAND2_X2 T7704 ( .B(T12328_Y), .A(T9809_Y), .Y(T7704_Y));
KC_NAND2_X2 T10320 ( .B(T6802_Y), .A(T6839_Y), .Y(T10320_Y));
KC_NAND2_X2 T8004 ( .B(T16397_Y), .A(T5331_Y), .Y(T8004_Y));
KC_NAND2_X2 T8003 ( .B(T1633_Y), .A(T6595_Y), .Y(T8003_Y));
KC_NAND2_X2 T8002 ( .B(T3683_Y), .A(T2589_Y), .Y(T8002_Y));
KC_NAND2_X2 T7322 ( .B(T1633_Y), .A(T6595_Y), .Y(T7322_Y));
KC_NAND2_X2 T5649 ( .B(T13710_Q), .A(T1637_Y), .Y(T5649_Y));
KC_NAND2_X2 T7702 ( .B(T1660_Q), .A(T1661_Q), .Y(T7702_Y));
KC_NAND2_X2 T10309 ( .B(T10305_Y), .A(T15069_Y), .Y(T10309_Y));
KC_NAND2_X2 T1687 ( .B(T16407_Y), .A(T2000_Y), .Y(T1687_Y));
KC_NAND2_X2 T1750 ( .B(T5794_Y), .A(T10224_Y), .Y(T1750_Y));
KC_NAND2_X2 T1762 ( .B(T5945_Y), .A(T5452_Q), .Y(T1762_Y));
KC_NAND2_X2 T1763 ( .B(T5904_Y), .A(T11493_Y), .Y(T1763_Y));
KC_NAND2_X2 T1766 ( .B(T16475_Y), .A(T1850_Y), .Y(T1766_Y));
KC_NAND2_X2 T1768 ( .B(T5903_Y), .A(T2150_Q), .Y(T1768_Y));
KC_NAND2_X2 T1782 ( .B(T4925_Q), .A(T12270_Y), .Y(T1782_Y));
KC_NAND2_X2 T1791 ( .B(T1820_Q), .A(T4965_Y), .Y(T1791_Y));
KC_NAND2_X2 T1793 ( .B(T1807_Q), .A(T11728_Y), .Y(T1793_Y));
KC_NAND2_X2 T1797 ( .B(T1807_Q), .A(T12270_Y), .Y(T1797_Y));
KC_NAND2_X2 T1810 ( .B(T1823_Q), .A(T12270_Y), .Y(T1810_Y));
KC_NAND2_X2 T1813 ( .B(T1822_Q), .A(T4965_Y), .Y(T1813_Y));
KC_NAND2_X2 T1814 ( .B(T1821_Q), .A(T4965_Y), .Y(T1814_Y));
KC_NAND2_X2 T1818 ( .B(T1826_Q), .A(T12270_Y), .Y(T1818_Y));
KC_NAND2_X2 T1985 ( .B(T15478_Y), .A(T2008_Q), .Y(T1985_Y));
KC_NAND2_X2 T1990 ( .B(T2008_Q), .A(T2015_Q), .Y(T1990_Y));
KC_NAND2_X2 T1991 ( .B(T11949_Y), .A(T15478_Y), .Y(T1991_Y));
KC_NAND2_X2 T1992 ( .B(T11949_Y), .A(T1142_Y), .Y(T1992_Y));
KC_NAND2_X2 T1993 ( .B(T11949_Y), .A(T2008_Q), .Y(T1993_Y));
KC_NAND2_X2 T1994 ( .B(T2008_Q), .A(T2023_Q), .Y(T1994_Y));
KC_NAND2_X2 T1999 ( .B(T1991_Y), .A(T5881_Y), .Y(T1999_Y));
KC_NAND2_X2 T2030 ( .B(T15503_Y), .A(T16268_Y), .Y(T2030_Y));
KC_NAND2_X2 T2031 ( .B(T2033_Y), .A(T10079_Y), .Y(T2031_Y));
KC_NAND2_X2 T2034 ( .B(T2550_Y), .A(T12736_Y), .Y(T2034_Y));
KC_NAND2_X2 T2035 ( .B(T10079_Y), .A(T5367_Y), .Y(T2035_Y));
KC_NAND2_X2 T2037 ( .B(T1117_Y), .A(T16365_Y), .Y(T2037_Y));
KC_NAND2_X2 T2038 ( .B(T2604_Y), .A(T2034_Y), .Y(T2038_Y));
KC_NAND2_X2 T2039 ( .B(T1518_Y), .A(T16411_Y), .Y(T2039_Y));
KC_NAND2_X2 T2040 ( .B(T10062_Y), .A(T2550_Y), .Y(T2040_Y));
KC_NAND2_X2 T2068 ( .B(T13131_Y), .A(T16274_Y), .Y(T2068_Y));
KC_NAND2_X2 T2072 ( .B(T8219_Y), .A(T8313_Y), .Y(T2072_Y));
KC_NAND2_X2 T15829 ( .B(T8183_Y), .A(T8182_Y), .Y(T15829_Y));
KC_NAND2_X2 T2104 ( .B(T15942_Y), .A(T16018_Q), .Y(T2104_Y));
KC_NAND2_X2 T2105 ( .B(T11489_Y), .A(T2109_Y), .Y(T2105_Y));
KC_NAND2_X2 T2132 ( .B(T15942_Y), .A(T16007_Q), .Y(T2132_Y));
KC_NAND2_X2 T2140 ( .B(T15942_Y), .A(T2835_Q), .Y(T2140_Y));
KC_NAND2_X2 T2145 ( .B(T15942_Y), .A(T2275_Q), .Y(T2145_Y));
KC_NAND2_X2 T2149 ( .B(T8497_Y), .A(T2722_Y), .Y(T2149_Y));
KC_NAND2_X2 T2165 ( .B(T15942_Y), .A(T2281_Q), .Y(T2165_Y));
KC_NAND2_X2 T2168 ( .B(T15942_Y), .A(T6007_Y), .Y(T2168_Y));
KC_NAND2_X2 T2170 ( .B(T2165_Y), .A(T11529_Y), .Y(T2170_Y));
KC_NAND2_X2 T2171 ( .B(T16156_Y), .A(T2839_Y), .Y(T2171_Y));
KC_NAND2_X2 T2172 ( .B(T5924_Y), .A(T15959_Y), .Y(T2172_Y));
KC_NAND2_X2 T2173 ( .B(T2167_Y), .A(T2167_Y), .Y(T2173_Y));
KC_NAND2_X2 T2215 ( .B(T6003_Y), .A(T12108_Y), .Y(T2215_Y));
KC_NAND2_X2 T2216 ( .B(T6003_Y), .A(T12103_Y), .Y(T2216_Y));
KC_NAND2_X2 T2217 ( .B(T12263_Y), .A(T15234_Y), .Y(T2217_Y));
KC_NAND2_X2 T2231 ( .B(T6003_Y), .A(T16270_Y), .Y(T2231_Y));
KC_NAND2_X2 T2259 ( .B(T11652_Y), .A(T16042_Y), .Y(T2259_Y));
KC_NAND2_X2 T2260 ( .B(T2819_Y), .A(T2249_Q), .Y(T2260_Y));
KC_NAND2_X2 T2261 ( .B(T2264_Y), .A(T16041_Y), .Y(T2261_Y));
KC_NAND2_X2 T2266 ( .B(T2876_Y), .A(T12108_Y), .Y(T2266_Y));
KC_NAND2_X2 T2267 ( .B(T2819_Y), .A(T2275_Q), .Y(T2267_Y));
KC_NAND2_X2 T2268 ( .B(T2876_Y), .A(T16270_Y), .Y(T2268_Y));
KC_NAND2_X2 T2271 ( .B(T2876_Y), .A(T12101_Y), .Y(T2271_Y));
KC_NAND2_X2 T2282 ( .B(T2876_Y), .A(T12105_Y), .Y(T2282_Y));
KC_NAND2_X2 T2283 ( .B(T2876_Y), .A(T12102_Y), .Y(T2283_Y));
KC_NAND2_X2 T2284 ( .B(T2876_Y), .A(T12107_Y), .Y(T2284_Y));
KC_NAND2_X2 T2293 ( .B(T10597_Y), .A(T2247_Y), .Y(T2293_Y));
KC_NAND2_X2 T2298 ( .B(T10626_Y), .A(T2240_Y), .Y(T2298_Y));
KC_NAND2_X2 T2299 ( .B(T2876_Y), .A(T12106_Y), .Y(T2299_Y));
KC_NAND2_X2 T2300 ( .B(T2876_Y), .A(T12103_Y), .Y(T2300_Y));
KC_NAND2_X2 T2325 ( .B(T10557_Y), .A(T12105_Y), .Y(T2325_Y));
KC_NAND2_X2 T2326 ( .B(T6227_Y), .A(T11776_Y), .Y(T2326_Y));
KC_NAND2_X2 T2327 ( .B(T2326_Y), .A(T6227_Y), .Y(T2327_Y));
KC_NAND2_X2 T2328 ( .B(T1832_Q), .A(T1833_Q), .Y(T2328_Y));
KC_NAND2_X2 T2332 ( .B(T2329_Y), .A(T12101_Y), .Y(T2332_Y));
KC_NAND2_X2 T2333 ( .B(T6198_Y), .A(T11772_Y), .Y(T2333_Y));
KC_NAND2_X2 T2334 ( .B(T11750_Y), .A(T11837_Y), .Y(T2334_Y));
KC_NAND2_X2 T2335 ( .B(T2328_Y), .A(T11775_Y), .Y(T2335_Y));
KC_NAND2_X2 T2338 ( .B(T2362_Y), .A(T2373_Y), .Y(T2338_Y));
KC_NAND2_X2 T2339 ( .B(T2338_Y), .A(T15628_Y), .Y(T2339_Y));
KC_NAND2_X2 T2372 ( .B(T1856_Q), .A(T2388_Q), .Y(T2372_Y));
KC_NAND2_X2 T2446 ( .B(T3589_Y), .A(T14984_Y), .Y(T2446_Y));
KC_NAND2_X2 T2447 ( .B(T2449_Y), .A(T14984_Y), .Y(T2447_Y));
KC_NAND2_X2 T2454 ( .B(T14859_Q), .A(T16079_Q), .Y(T2454_Y));
KC_NAND2_X2 T2457 ( .B(T2464_Y), .A(T2458_Y), .Y(T2457_Y));
KC_NAND2_X2 T2458 ( .B(T3605_Y), .A(T14984_Y), .Y(T2458_Y));
KC_NAND2_X2 T2459 ( .B(T12080_Y), .A(T9774_Y), .Y(T2459_Y));
KC_NAND2_X2 T2460 ( .B(T2478_Y), .A(T9745_Y), .Y(T2460_Y));
KC_NAND2_X2 T2464 ( .B(T15442_Y), .A(T13895_Q), .Y(T2464_Y));
KC_NAND2_X2 T2465 ( .B(T9779_Y), .A(T9854_Y), .Y(T2465_Y));
KC_NAND2_X2 T2466 ( .B(T13895_Q), .A(T16079_Q), .Y(T2466_Y));
KC_NAND2_X2 T2467 ( .B(T9772_Y), .A(T2674_Y), .Y(T2467_Y));
KC_NAND2_X2 T2476 ( .B(T13835_Q), .A(T16079_Q), .Y(T2476_Y));
KC_NAND2_X2 T2477 ( .B(T10493_Y), .A(T9854_Y), .Y(T2477_Y));
KC_NAND2_X2 T2478 ( .B(T13716_Q), .A(T16079_Q), .Y(T2478_Y));
KC_NAND2_X2 T2480 ( .B(T15419_Y), .A(T610_Y), .Y(T2480_Y));
KC_NAND2_X2 T2481 ( .B(T9772_Y), .A(T11174_Y), .Y(T2481_Y));
KC_NAND2_X2 T2482 ( .B(T634_Y), .A(T15419_Y), .Y(T2482_Y));
KC_NAND2_X2 T2500 ( .B(T882_Y), .A(T2861_Y), .Y(T2500_Y));
KC_NAND2_X2 T2501 ( .B(T16447_Y), .A(T16195_Y), .Y(T2501_Y));
KC_NAND2_X2 T2502 ( .B(T883_Y), .A(T882_Y), .Y(T2502_Y));
KC_NAND2_X2 T2507 ( .B(T5314_Y), .A(T5318_Y), .Y(T2507_Y));
KC_NAND2_X2 T2508 ( .B(T9780_Y), .A(T9874_Y), .Y(T2508_Y));
KC_NAND2_X2 T2520 ( .B(T2592_Q), .A(T2591_Q), .Y(T2520_Y));
KC_NAND2_X2 T2545 ( .B(T2575_Q), .A(T10518_Y), .Y(T2545_Y));
KC_NAND2_X2 T2547 ( .B(T13032_Y), .A(T2013_Y), .Y(T2547_Y));
KC_NAND2_X2 T2548 ( .B(T2564_Y), .A(T3692_Y), .Y(T2548_Y));
KC_NAND2_X2 T2549 ( .B(T13894_Q), .A(T10251_Y), .Y(T2549_Y));
KC_NAND2_X2 T2558 ( .B(T14995_Y), .A(T4307_Y), .Y(T2558_Y));
KC_NAND2_X2 T2559 ( .B(T14995_Y), .A(T3103_Y), .Y(T2559_Y));
KC_NAND2_X2 T2560 ( .B(T10942_Y), .A(T10941_Y), .Y(T2560_Y));
KC_NAND2_X2 T2597 ( .B(T10102_Y), .A(T15518_Y), .Y(T2597_Y));
KC_NAND2_X2 T2598 ( .B(T2717_Y), .A(T11662_Y), .Y(T2598_Y));
KC_NAND2_X2 T2608 ( .B(T13032_Y), .A(T10526_Y), .Y(T2608_Y));
KC_NAND2_X2 T2609 ( .B(T2832_Q), .A(T10090_Y), .Y(T2609_Y));
KC_NAND2_X2 T2610 ( .B(T10105_Y), .A(T12735_Y), .Y(T2610_Y));
KC_NAND2_X2 T2611 ( .B(T2057_Y), .A(T10080_Y), .Y(T2611_Y));
KC_NAND2_X2 T2614 ( .B(T3720_Y), .A(T14995_Y), .Y(T2614_Y));
KC_NAND2_X2 T2632 ( .B(T4981_Y), .A(T15535_Y), .Y(T2632_Y));
KC_NAND2_X2 T2633 ( .B(T10880_Y), .A(T10188_Y), .Y(T2633_Y));
KC_NAND2_X2 T2652 ( .B(T5751_Y), .A(T10277_Y), .Y(T2652_Y));
KC_NAND2_X2 T2653 ( .B(T10277_Y), .A(T5421_Q), .Y(T2653_Y));
KC_NAND2_X2 T2654 ( .B(T10280_Y), .A(T5749_Y), .Y(T2654_Y));
KC_NAND2_X2 T2655 ( .B(T10278_Y), .A(T5421_Q), .Y(T2655_Y));
KC_NAND2_X2 T2660 ( .B(T5724_Y), .A(T2063_Y), .Y(T2660_Y));
KC_NAND2_X2 T2661 ( .B(T5717_Y), .A(T5710_Y), .Y(T2661_Y));
KC_NAND2_X2 T2662 ( .B(T5717_Y), .A(T5425_Q), .Y(T2662_Y));
KC_NAND2_X2 T2663 ( .B(T5710_Y), .A(T5424_Q), .Y(T2663_Y));
KC_NAND2_X2 T2664 ( .B(T5424_Q), .A(T5425_Q), .Y(T2664_Y));
KC_NAND2_X2 T15827 ( .B(T15754_Y), .A(T5019_Y), .Y(T15827_Y));
KC_NAND2_X2 T2675 ( .B(T15696_Y), .A(T5714_Y), .Y(T2675_Y));
KC_NAND2_X2 T2676 ( .B(T11009_Y), .A(T2675_Y), .Y(T2676_Y));
KC_NAND2_X2 T2677 ( .B(T15696_Y), .A(T5425_Q), .Y(T2677_Y));
KC_NAND2_X2 T2678 ( .B(T5766_Y), .A(T15753_Y), .Y(T2678_Y));
KC_NAND2_X2 T2680 ( .B(T2696_Y), .A(T11338_Y), .Y(T2680_Y));
KC_NAND2_X2 T2681 ( .B(T11357_Y), .A(T5758_Y), .Y(T2681_Y));
KC_NAND2_X2 T2682 ( .B(T15442_Y), .A(T2656_Y), .Y(T2682_Y));
KC_NAND2_X2 T2683 ( .B(T2682_Y), .A(T10890_Y), .Y(T2683_Y));
KC_NAND2_X2 T2684 ( .B(T10891_Y), .A(T2695_Y), .Y(T2684_Y));
KC_NAND2_X2 T2686 ( .B(T11964_Y), .A(T14954_Q), .Y(T2686_Y));
KC_NAND2_X2 T2703 ( .B(T2706_Y), .A(T2124_Y), .Y(T2703_Y));
KC_NAND2_X2 T2722 ( .B(T15942_Y), .A(T2249_Q), .Y(T2722_Y));
KC_NAND2_X2 T2754 ( .B(T3411_Y), .A(T6235_Y), .Y(T2754_Y));
KC_NAND2_X2 T2777 ( .B(T5070_Y), .A(T5570_Y), .Y(T2777_Y));
KC_NAND2_X2 T2778 ( .B(T5570_Y), .A(T6526_Q), .Y(T2778_Y));
KC_NAND2_X2 T2779 ( .B(T2794_Q), .A(T2793_Q), .Y(T2779_Y));
KC_NAND2_X2 T2797 ( .B(T16023_Q), .A(T5990_Y), .Y(T2797_Y));
KC_NAND2_X2 T2800 ( .B(T6007_Y), .A(T11641_Y), .Y(T2800_Y));
KC_NAND2_X2 T2802 ( .B(T11633_Y), .A(T15234_Y), .Y(T2802_Y));
KC_NAND2_X2 T2803 ( .B(T6007_Y), .A(T11604_Y), .Y(T2803_Y));
KC_NAND2_X2 T2804 ( .B(T15942_Y), .A(T2843_Q), .Y(T2804_Y));
KC_NAND2_X2 T2805 ( .B(T16038_Y), .A(T10740_Y), .Y(T2805_Y));
KC_NAND2_X2 T2816 ( .B(T2819_Y), .A(T2835_Q), .Y(T2816_Y));
KC_NAND2_X2 T2817 ( .B(T11727_Y), .A(T15138_Q), .Y(T2817_Y));
KC_NAND2_X2 T2820 ( .B(T15942_Y), .A(T16023_Q), .Y(T2820_Y));
KC_NAND2_X2 T2821 ( .B(T5010_Y), .A(T2820_Y), .Y(T2821_Y));
KC_NAND2_X2 T2824 ( .B(T11666_Y), .A(T16305_Y), .Y(T2824_Y));
KC_NAND2_X2 T2849 ( .B(T3530_Y), .A(T1285_Y), .Y(T2849_Y));
KC_NAND2_X2 T2859 ( .B(T6180_Y), .A(T3526_Y), .Y(T2859_Y));
KC_NAND2_X2 T2860 ( .B(T12066_Y), .A(T6561_Y), .Y(T2860_Y));
KC_NAND2_X2 T2866 ( .B(T10591_Y), .A(T12065_Y), .Y(T2866_Y));
KC_NAND2_X2 T2867 ( .B(T4705_Y), .A(T10591_Y), .Y(T2867_Y));
KC_NAND2_X2 T2880 ( .B(T12038_Y), .A(T15621_Y), .Y(T2880_Y));
KC_NAND2_X2 T2881 ( .B(T15762_Y), .A(T6224_Y), .Y(T2881_Y));
KC_NAND2_X2 T2886 ( .B(T16131_Y), .A(T10573_Y), .Y(T2886_Y));
KC_NAND2_X2 T2887 ( .B(T2320_Y), .A(T10557_Y), .Y(T2887_Y));
KC_NAND2_X2 T2888 ( .B(T8417_Y), .A(T6193_Y), .Y(T2888_Y));
KC_NAND2_X2 T2891 ( .B(T2324_Y), .A(T2894_Y), .Y(T2891_Y));
KC_NAND2_X2 T2892 ( .B(T4999_Y), .A(T6572_Y), .Y(T2892_Y));
KC_NAND2_X2 T2896 ( .B(T15633_Y), .A(T11810_Y), .Y(T2896_Y));
KC_NAND2_X2 T2897 ( .B(T2901_Y), .A(T15632_Y), .Y(T2897_Y));
KC_NAND2_X2 T2898 ( .B(T6240_Y), .A(T15953_Y), .Y(T2898_Y));
KC_NAND2_X2 T2899 ( .B(T5518_Y), .A(T2901_Y), .Y(T2899_Y));
KC_NAND2_X2 T2900 ( .B(T2318_Y), .A(T2907_Y), .Y(T2900_Y));
KC_NAND2_X2 T2901 ( .B(T6223_Y), .A(T15627_Y), .Y(T2901_Y));
KC_NAND2_X2 T2902 ( .B(T6576_Y), .A(T2324_Y), .Y(T2902_Y));
KC_NAND2_X2 T2903 ( .B(T15627_Y), .A(T2354_Y), .Y(T2903_Y));
KC_NAND2_X2 T2907 ( .B(T6223_Y), .A(T6197_Y), .Y(T2907_Y));
KC_NAND2_X2 T2908 ( .B(T2320_Y), .A(T11774_Y), .Y(T2908_Y));
KC_NAND2_X2 T2909 ( .B(T2320_Y), .A(T15627_Y), .Y(T2909_Y));
KC_NAND2_X2 T2910 ( .B(T4054_Y), .A(T2948_Y), .Y(T2910_Y));
KC_NAND2_X2 T2911 ( .B(T11837_Y), .A(T6506_Y), .Y(T2911_Y));
KC_NAND2_X2 T2912 ( .B(T2908_Y), .A(T6195_Y), .Y(T2912_Y));
KC_NAND2_X2 T2915 ( .B(T4055_Y), .A(T2941_Y), .Y(T2915_Y));
KC_NAND2_X2 T2916 ( .B(T6561_Y), .A(T10554_Y), .Y(T2916_Y));
KC_NAND2_X2 T2932 ( .B(T2944_Q), .A(T2943_Q), .Y(T2932_Y));
KC_NAND2_X2 T2934 ( .B(T11005_Y), .A(T10570_Y), .Y(T2934_Y));
KC_NAND2_X2 T2935 ( .B(T6538_Y), .A(T4096_Y), .Y(T2935_Y));
KC_NAND2_X2 T2936 ( .B(T15643_Y), .A(T6537_Y), .Y(T2936_Y));
KC_NAND2_X2 T2937 ( .B(T3436_Y), .A(T6538_Y), .Y(T2937_Y));
KC_NAND2_X2 T2938 ( .B(T5540_Y), .A(T2959_Y), .Y(T2938_Y));
KC_NAND2_X2 T2939 ( .B(T6561_Y), .A(T11836_Y), .Y(T2939_Y));
KC_NAND2_X2 T3012 ( .B(T14984_Y), .A(T3586_Y), .Y(T3012_Y));
KC_NAND2_X2 T3013 ( .B(T1633_Y), .A(T6595_Y), .Y(T3013_Y));
KC_NAND2_X2 T3014 ( .B(T2451_Y), .A(T2589_Y), .Y(T3014_Y));
KC_NAND2_X2 T3020 ( .B(T2676_Y), .A(T15683_Y), .Y(T3020_Y));
KC_NAND2_X2 T3031 ( .B(T1633_Y), .A(T6595_Y), .Y(T3031_Y));
KC_NAND2_X2 T3045 ( .B(T2496_Y), .A(T10471_Y), .Y(T3045_Y));
KC_NAND2_X2 T3051 ( .B(T2451_Y), .A(T2589_Y), .Y(T3051_Y));
KC_NAND2_X2 T3068 ( .B(T3078_Y), .A(T3728_Y), .Y(T3068_Y));
KC_NAND2_X2 T3069 ( .B(T3683_Y), .A(T2589_Y), .Y(T3069_Y));
KC_NAND2_X2 T3093 ( .B(T3146_Y), .A(T14995_Y), .Y(T3093_Y));
KC_NAND2_X2 T3184 ( .B(T11309_Y), .A(T5747_Y), .Y(T3184_Y));
KC_NAND2_X2 T3200 ( .B(T5074_Q), .A(T3998_Y), .Y(T3200_Y));
KC_NAND2_X2 T3201 ( .B(T11356_Y), .A(T13067_Q), .Y(T3201_Y));
KC_NAND2_X2 T3202 ( .B(T3221_Y), .A(T11337_Y), .Y(T3202_Y));
KC_NAND2_X2 T3203 ( .B(T3816_Y), .A(T5806_Y), .Y(T3203_Y));
KC_NAND2_X2 T3204 ( .B(T11985_Y), .A(T11983_Y), .Y(T3204_Y));
KC_NAND2_X2 T3207 ( .B(T11370_Y), .A(T15865_Y), .Y(T3207_Y));
KC_NAND2_X2 T3223 ( .B(T14541_Q), .A(T14543_Q), .Y(T3223_Y));
KC_NAND2_X2 T3224 ( .B(T5039_Y), .A(T14540_Q), .Y(T3224_Y));
KC_NAND2_X2 T3286 ( .B(T5923_Y), .A(T3298_Y), .Y(T3286_Y));
KC_NAND2_X2 T3297 ( .B(T3299_Y), .A(T3307_Y), .Y(T3297_Y));
KC_NAND2_X2 T3328 ( .B(T3316_Y), .A(T11545_Y), .Y(T3328_Y));
KC_NAND2_X2 T3354 ( .B(T16035_Y), .A(T5072_Y), .Y(T3354_Y));
KC_NAND2_X2 T3355 ( .B(T5070_Y), .A(T5072_Y), .Y(T3355_Y));
KC_NAND2_X2 T3368 ( .B(T10970_Y), .A(T10585_Y), .Y(T3368_Y));
KC_NAND2_X2 T3369 ( .B(T6065_Y), .A(T12317_Y), .Y(T3369_Y));
KC_NAND2_X2 T3370 ( .B(T11625_Y), .A(T12045_Y), .Y(T3370_Y));
KC_NAND2_X2 T3374 ( .B(T15760_Q), .A(T4179_Q), .Y(T3374_Y));
KC_NAND2_X2 T3375 ( .B(T4179_Q), .A(T4176_Q), .Y(T3375_Y));
KC_NAND2_X2 T3376 ( .B(T16037_Y), .A(T12043_Y), .Y(T3376_Y));
KC_NAND2_X2 T3379 ( .B(T8385_Y), .A(T11746_Y), .Y(T3379_Y));
KC_NAND2_X2 T3382 ( .B(T11661_Y), .A(T6585_Y), .Y(T3382_Y));
KC_NAND2_X2 T3383 ( .B(T11647_Y), .A(T6585_Y), .Y(T3383_Y));
KC_NAND2_X2 T3384 ( .B(T6065_Y), .A(T11818_Y), .Y(T3384_Y));
KC_NAND2_X2 T3393 ( .B(T6048_Y), .A(T11627_Y), .Y(T3393_Y));
KC_NAND2_X2 T3394 ( .B(T6526_Q), .A(T6549_Q), .Y(T3394_Y));
KC_NAND2_X2 T3395 ( .B(T6080_Y), .A(T6067_Y), .Y(T3395_Y));
KC_NAND2_X2 T3396 ( .B(T6080_Y), .A(T3516_Y), .Y(T3396_Y));
KC_NAND2_X2 T3397 ( .B(T3399_Y), .A(T12043_Y), .Y(T3397_Y));
KC_NAND2_X2 T3400 ( .B(T11627_Y), .A(T5525_Q), .Y(T3400_Y));
KC_NAND2_X2 T3401 ( .B(T3411_Y), .A(T11643_Y), .Y(T3401_Y));
KC_NAND2_X2 T3415 ( .B(T6160_Y), .A(T6236_Y), .Y(T3415_Y));
KC_NAND2_X2 T3416 ( .B(T6236_Y), .A(T12044_Y), .Y(T3416_Y));
KC_NAND2_X2 T3417 ( .B(T6547_Y), .A(T11818_Y), .Y(T3417_Y));
KC_NAND2_X2 T3424 ( .B(T6067_Y), .A(T6120_Y), .Y(T3424_Y));
KC_NAND2_X2 T3426 ( .B(T15616_Y), .A(T5510_Y), .Y(T3426_Y));
KC_NAND2_X2 T3427 ( .B(T6547_Y), .A(T6139_Y), .Y(T3427_Y));
KC_NAND2_X2 T3428 ( .B(T4060_Y), .A(T6532_Y), .Y(T3428_Y));
KC_NAND2_X2 T3429 ( .B(T6112_Y), .A(T11746_Y), .Y(T3429_Y));
KC_NAND2_X2 T3435 ( .B(T3385_Y), .A(T4024_Y), .Y(T3435_Y));
KC_NAND2_X2 T3436 ( .B(T6098_Y), .A(T11746_Y), .Y(T3436_Y));
KC_NAND2_X2 T3437 ( .B(T10610_Y), .A(T12265_Y), .Y(T3437_Y));
KC_NAND2_X2 T3438 ( .B(T10611_Y), .A(T12265_Y), .Y(T3438_Y));
KC_NAND2_X2 T3439 ( .B(T16167_Y), .A(T10585_Y), .Y(T3439_Y));
KC_NAND2_X2 T3443 ( .B(T11746_Y), .A(T6096_Y), .Y(T3443_Y));
KC_NAND2_X2 T3444 ( .B(T12263_Y), .A(T16102_Y), .Y(T3444_Y));
KC_NAND2_X2 T3445 ( .B(T16167_Y), .A(T12317_Y), .Y(T3445_Y));
KC_NAND2_X2 T3446 ( .B(T6080_Y), .A(T3368_Y), .Y(T3446_Y));
KC_NAND2_X2 T3447 ( .B(T6138_Y), .A(T6049_Y), .Y(T3447_Y));
KC_NAND2_X2 T3448 ( .B(T6106_Y), .A(T15234_Y), .Y(T3448_Y));
KC_NAND2_X2 T3465 ( .B(T2800_Y), .A(T11816_Y), .Y(T3465_Y));
KC_NAND2_X2 T3466 ( .B(T11673_Y), .A(T3517_Y), .Y(T3466_Y));
KC_NAND2_X2 T3467 ( .B(T16102_Y), .A(T6585_Y), .Y(T3467_Y));
KC_NAND2_X2 T3468 ( .B(T6209_Y), .A(T6156_Y), .Y(T3468_Y));
KC_NAND2_X2 T3469 ( .B(T16138_Y), .A(T11802_Y), .Y(T3469_Y));
KC_NAND2_X2 T3473 ( .B(T11644_Y), .A(T6158_Y), .Y(T3473_Y));
KC_NAND2_X2 T3474 ( .B(T5109_Y), .A(T10550_Y), .Y(T3474_Y));
KC_NAND2_X2 T3475 ( .B(T5047_Y), .A(T5519_Y), .Y(T3475_Y));
KC_NAND2_X2 T3477 ( .B(T3465_Y), .A(T10548_Y), .Y(T3477_Y));
KC_NAND2_X2 T3478 ( .B(T6550_Y), .A(T4164_Q), .Y(T3478_Y));
KC_NAND2_X2 T3479 ( .B(T10553_Y), .A(T12108_Y), .Y(T3479_Y));
KC_NAND2_X2 T3480 ( .B(T8407_Y), .A(T6560_Y), .Y(T3480_Y));
KC_NAND2_X2 T3481 ( .B(T6193_Y), .A(T6560_Y), .Y(T3481_Y));
KC_NAND2_X2 T3489 ( .B(T6561_Y), .A(T11742_Y), .Y(T3489_Y));
KC_NAND2_X2 T3490 ( .B(T11822_Y), .A(T8426_Y), .Y(T3490_Y));
KC_NAND2_X2 T3506 ( .B(T6489_Y), .A(T3522_Q), .Y(T3506_Y));
KC_NAND2_X2 T3508 ( .B(T11843_Y), .A(T3521_Q), .Y(T3508_Y));
KC_NAND2_X2 T3509 ( .B(T6490_Y), .A(T6561_Y), .Y(T3509_Y));
KC_NAND2_X2 T3510 ( .B(T11835_Y), .A(T3525_Q), .Y(T3510_Y));
KC_NAND2_X2 T3511 ( .B(T6512_Y), .A(T11835_Y), .Y(T3511_Y));
KC_NAND2_X2 T3512 ( .B(T6512_Y), .A(T3519_Q), .Y(T3512_Y));
KC_NAND2_X2 T3514 ( .B(T11833_Y), .A(T11832_Y), .Y(T3514_Y));
KC_NAND2_X2 T3515 ( .B(T8426_Y), .A(T11823_Y), .Y(T3515_Y));
KC_NAND2_X2 T3607 ( .B(T6802_Y), .A(T6839_Y), .Y(T3607_Y));
KC_NAND2_X2 T3608 ( .B(T622_Y), .A(T5331_Y), .Y(T3608_Y));
KC_NAND2_X2 T3621 ( .B(T622_Y), .A(T5331_Y), .Y(T3621_Y));
KC_NAND2_X2 T3626 ( .B(T6802_Y), .A(T6839_Y), .Y(T3626_Y));
KC_NAND2_X2 T3651 ( .B(T6802_Y), .A(T6839_Y), .Y(T3651_Y));
KC_NAND2_X2 T3654 ( .B(T1633_Y), .A(T6595_Y), .Y(T3654_Y));
KC_NAND2_X2 T3666 ( .B(T622_Y), .A(T5331_Y), .Y(T3666_Y));
KC_NAND2_X2 T3667 ( .B(T3683_Y), .A(T2589_Y), .Y(T3667_Y));
KC_NAND2_X2 T3668 ( .B(T1633_Y), .A(T6595_Y), .Y(T3668_Y));
KC_NAND2_X2 T3712 ( .B(T622_Y), .A(T5331_Y), .Y(T3712_Y));
KC_NAND2_X2 T3787 ( .B(T5781_Y), .A(T3841_Y), .Y(T3787_Y));
KC_NAND2_X2 T3788 ( .B(T145_Q), .A(T15908_Y), .Y(T3788_Y));
KC_NAND2_X2 T3789 ( .B(T4486_Y), .A(T15868_Y), .Y(T3789_Y));
KC_NAND2_X2 T3790 ( .B(T15870_Y), .A(T11379_Y), .Y(T3790_Y));
KC_NAND2_X2 T3791 ( .B(T15825_Y), .A(T15835_Y), .Y(T3791_Y));
KC_NAND2_X2 T3794 ( .B(T4486_Y), .A(T144_Q), .Y(T3794_Y));
KC_NAND2_X2 T3795 ( .B(T15888_Y), .A(T145_Q), .Y(T3795_Y));
KC_NAND2_X2 T3796 ( .B(T5801_Y), .A(T4465_Q), .Y(T3796_Y));
KC_NAND2_X2 T3797 ( .B(T4486_Y), .A(T15888_Y), .Y(T3797_Y));
KC_NAND2_X2 T3800 ( .B(T15845_Y), .A(T16153_Y), .Y(T3800_Y));
KC_NAND2_X2 T3801 ( .B(T11983_Y), .A(T11379_Y), .Y(T3801_Y));
KC_NAND2_X2 T3802 ( .B(T11353_Y), .A(T16153_Y), .Y(T3802_Y));
KC_NAND2_X2 T3803 ( .B(T5767_Y), .A(T11365_Y), .Y(T3803_Y));
KC_NAND2_X2 T3804 ( .B(T15868_Y), .A(T5763_Y), .Y(T3804_Y));
KC_NAND2_X2 T3805 ( .B(T11336_Y), .A(T15877_Y), .Y(T3805_Y));
KC_NAND2_X2 T3806 ( .B(T4389_Y), .A(T5767_Y), .Y(T3806_Y));
KC_NAND2_X2 T3815 ( .B(T15870_Y), .A(T5763_Y), .Y(T3815_Y));
KC_NAND2_X2 T3816 ( .B(T15845_Y), .A(T11410_Y), .Y(T3816_Y));
KC_NAND2_X2 T3824 ( .B(T11367_Y), .A(T11410_Y), .Y(T3824_Y));
KC_NAND2_X2 T3825 ( .B(T5815_Y), .A(T15908_Y), .Y(T3825_Y));
KC_NAND2_X2 T3826 ( .B(T15907_Y), .A(T15908_Y), .Y(T3826_Y));
KC_NAND2_X2 T3827 ( .B(T5788_Y), .A(T16154_Y), .Y(T3827_Y));
KC_NAND2_X2 T3831 ( .B(T11410_Y), .A(T144_Q), .Y(T3831_Y));
KC_NAND2_X2 T3832 ( .B(T4438_Y), .A(T144_Q), .Y(T3832_Y));
KC_NAND2_X2 T3833 ( .B(T11367_Y), .A(T144_Q), .Y(T3833_Y));
KC_NAND2_X2 T3834 ( .B(T15897_Y), .A(T15908_Y), .Y(T3834_Y));
KC_NAND2_X2 T3835 ( .B(T11322_Y), .A(T5826_Y), .Y(T3835_Y));
KC_NAND2_X2 T3836 ( .B(T5815_Y), .A(T5830_Y), .Y(T3836_Y));
KC_NAND2_X2 T3839 ( .B(T5801_Y), .A(T144_Q), .Y(T3839_Y));
KC_NAND2_X2 T3840 ( .B(T15877_Y), .A(T4500_Y), .Y(T3840_Y));
KC_NAND2_X2 T3841 ( .B(T5767_Y), .A(T11378_Y), .Y(T3841_Y));
KC_NAND2_X2 T3842 ( .B(T11378_Y), .A(T15908_Y), .Y(T3842_Y));
KC_NAND2_X2 T3843 ( .B(T4486_Y), .A(T11408_Y), .Y(T3843_Y));
KC_NAND2_X2 T3849 ( .B(T5788_Y), .A(T4487_Q), .Y(T3849_Y));
KC_NAND2_X2 T3850 ( .B(T4486_Y), .A(T16154_Y), .Y(T3850_Y));
KC_NAND2_X2 T3851 ( .B(T12174_Y), .A(T15896_Y), .Y(T3851_Y));
KC_NAND2_X2 T3857 ( .B(T5852_Y), .A(T11367_Y), .Y(T3857_Y));
KC_NAND2_X2 T3860 ( .B(T2073_Y), .A(T5985_Y), .Y(T3860_Y));
KC_NAND2_X2 T3866 ( .B(T15919_Y), .A(T15919_Y), .Y(T3866_Y));
KC_NAND2_X2 T3871 ( .B(T5868_Y), .A(T5140_Y), .Y(T3871_Y));
KC_NAND2_X2 T3901 ( .B(T10228_Y), .A(T4523_Y), .Y(T3901_Y));
KC_NAND2_X2 T3902 ( .B(T15580_Y), .A(T4508_Y), .Y(T3902_Y));
KC_NAND2_X2 T3905 ( .B(T5458_Y), .A(T5892_Y), .Y(T3905_Y));
KC_NAND2_X2 T3906 ( .B(T11023_Y), .A(T15961_Y), .Y(T3906_Y));
KC_NAND2_X2 T3912 ( .B(T3933_Y), .A(T3935_Q), .Y(T3912_Y));
KC_NAND2_X2 T3913 ( .B(T3908_Y), .A(T10958_Y), .Y(T3913_Y));
KC_NAND2_X2 T3914 ( .B(T5892_Y), .A(T3933_Y), .Y(T3914_Y));
KC_NAND2_X2 T3916 ( .B(T5458_Y), .A(T13115_Y), .Y(T3916_Y));
KC_NAND2_X2 T3917 ( .B(T5986_Y), .A(T12205_Y), .Y(T3917_Y));
KC_NAND2_X2 T3918 ( .B(T5099_Y), .A(T6204_Y), .Y(T3918_Y));
KC_NAND2_X2 T3919 ( .B(T15945_Y), .A(T11534_Y), .Y(T3919_Y));
KC_NAND2_X2 T3941 ( .B(T3949_Y), .A(T11616_Y), .Y(T3941_Y));
KC_NAND2_X2 T3944 ( .B(T15587_Y), .A(T3968_Q), .Y(T3944_Y));
KC_NAND2_X2 T3945 ( .B(T11577_Y), .A(T3965_Q), .Y(T3945_Y));
KC_NAND2_X2 T3946 ( .B(T5973_Y), .A(T11577_Y), .Y(T3946_Y));
KC_NAND2_X2 T3947 ( .B(T3968_Q), .A(T3974_Q), .Y(T3947_Y));
KC_NAND2_X2 T3949 ( .B(T3974_Q), .A(T5981_Y), .Y(T3949_Y));
KC_NAND2_X2 T3975 ( .B(T11615_Y), .A(T5476_Y), .Y(T3975_Y));
KC_NAND2_X2 T3976 ( .B(T6022_Y), .A(T4586_Y), .Y(T3976_Y));
KC_NAND2_X2 T3977 ( .B(T4583_Y), .A(T4584_Y), .Y(T3977_Y));
KC_NAND2_X2 T3978 ( .B(T6025_Y), .A(T5122_Y), .Y(T3978_Y));
KC_NAND2_X2 T4015 ( .B(T6077_Y), .A(T4748_Y), .Y(T4015_Y));
KC_NAND2_X2 T4016 ( .B(T5466_Y), .A(T4748_Y), .Y(T4016_Y));
KC_NAND2_X2 T4017 ( .B(T12043_Y), .A(T6045_Y), .Y(T4017_Y));
KC_NAND2_X2 T4024 ( .B(T6062_Y), .A(T5070_Y), .Y(T4024_Y));
KC_NAND2_X2 T4025 ( .B(T4052_Q), .A(T8167_Y), .Y(T4025_Y));
KC_NAND2_X2 T4031 ( .B(T6175_Y), .A(T5530_Q), .Y(T4031_Y));
KC_NAND2_X2 T4032 ( .B(T11638_Y), .A(T4179_Q), .Y(T4032_Y));
KC_NAND2_X2 T4033 ( .B(T11671_Y), .A(T5525_Q), .Y(T4033_Y));
KC_NAND2_X2 T4034 ( .B(T6034_Y), .A(T4147_Q), .Y(T4034_Y));
KC_NAND2_X2 T4035 ( .B(T6175_Y), .A(T6034_Y), .Y(T4035_Y));
KC_NAND2_X2 T4036 ( .B(T4147_Q), .A(T5530_Q), .Y(T4036_Y));
KC_NAND2_X2 T4057 ( .B(T4068_Y), .A(T6174_Y), .Y(T4057_Y));
KC_NAND2_X2 T4058 ( .B(T8502_Y), .A(T5135_Y), .Y(T4058_Y));
KC_NAND2_X2 T4059 ( .B(T4060_Y), .A(T11711_Y), .Y(T4059_Y));
KC_NAND2_X2 T4060 ( .B(T4589_Y), .A(T11709_Y), .Y(T4060_Y));
KC_NAND2_X2 T4061 ( .B(T6078_Y), .A(T11709_Y), .Y(T4061_Y));
KC_NAND2_X2 T4062 ( .B(T4023_Y), .A(T15760_Q), .Y(T4062_Y));
KC_NAND2_X2 T4067 ( .B(T4061_Y), .A(T12279_Y), .Y(T4067_Y));
KC_NAND2_X2 T4068 ( .B(T15619_Y), .A(T10581_Y), .Y(T4068_Y));
KC_NAND2_X2 T4069 ( .B(T3433_Y), .A(T6547_Y), .Y(T4069_Y));
KC_NAND2_X2 T4073 ( .B(T6137_Y), .A(T6135_Y), .Y(T4073_Y));
KC_NAND2_X2 T4074 ( .B(T6135_Y), .A(T5510_Y), .Y(T4074_Y));
KC_NAND2_X2 T4075 ( .B(T4074_Y), .A(T11710_Y), .Y(T4075_Y));
KC_NAND2_X2 T4076 ( .B(T6098_Y), .A(T15620_Y), .Y(T4076_Y));
KC_NAND2_X2 T4077 ( .B(T15912_Y), .A(T16124_Y), .Y(T4077_Y));
KC_NAND2_X2 T4078 ( .B(T2752_Q), .A(T4081_Y), .Y(T4078_Y));
KC_NAND2_X2 T4079 ( .B(T4080_Y), .A(T11710_Y), .Y(T4079_Y));
KC_NAND2_X2 T4082 ( .B(T12268_Y), .A(T15233_Y), .Y(T4082_Y));
KC_NAND2_X2 T4083 ( .B(T10617_Y), .A(T6096_Y), .Y(T4083_Y));
KC_NAND2_X2 T4084 ( .B(T6157_Y), .A(T11715_Y), .Y(T4084_Y));
KC_NAND2_X2 T4085 ( .B(T4027_Y), .A(T10584_Y), .Y(T4085_Y));
KC_NAND2_X2 T4091 ( .B(T4084_Y), .A(T10586_Y), .Y(T4091_Y));
KC_NAND2_X2 T4092 ( .B(T6157_Y), .A(T10586_Y), .Y(T4092_Y));
KC_NAND2_X2 T4093 ( .B(T2803_Y), .A(T4062_Y), .Y(T4093_Y));
KC_NAND2_X2 T4119 ( .B(T6207_Y), .A(T6587_Y), .Y(T4119_Y));
KC_NAND2_X2 T4127 ( .B(T10566_Y), .A(T10581_Y), .Y(T4127_Y));
KC_NAND2_X2 T4128 ( .B(T12287_Y), .A(T4137_Y), .Y(T4128_Y));
KC_NAND2_X2 T4139 ( .B(T4127_Y), .A(T4120_Y), .Y(T4139_Y));
KC_NAND2_X2 T4140 ( .B(T11687_Y), .A(T10581_Y), .Y(T4140_Y));
KC_NAND2_X2 T4202 ( .B(T15441_Y), .A(T16449_Y), .Y(T4202_Y));
KC_NAND2_X2 T4203 ( .B(T12082_Y), .A(T10431_Y), .Y(T4203_Y));
KC_NAND2_X2 T4204 ( .B(T10431_Y), .A(T12082_Y), .Y(T4204_Y));
KC_NAND2_X2 T4205 ( .B(T16449_Y), .A(T3073_Y), .Y(T4205_Y));
KC_NAND2_X2 T4265 ( .B(T3679_Y), .A(T3073_Y), .Y(T4265_Y));
KC_NAND2_X2 T4266 ( .B(T2530_Y), .A(T9858_Y), .Y(T4266_Y));
KC_NAND2_X2 T4267 ( .B(T9858_Y), .A(T2530_Y), .Y(T4267_Y));
KC_NAND2_X2 T4268 ( .B(T15441_Y), .A(T3679_Y), .Y(T4268_Y));
KC_NAND2_X2 T4318 ( .B(T10115_Y), .A(T12761_Y), .Y(T4318_Y));
KC_NAND2_X2 T4382 ( .B(T4403_Y), .A(T15871_Y), .Y(T4382_Y));
KC_NAND2_X2 T4383 ( .B(T5838_Y), .A(T16154_Y), .Y(T4383_Y));
KC_NAND2_X2 T4387 ( .B(T4403_Y), .A(T11378_Y), .Y(T4387_Y));
KC_NAND2_X2 T4388 ( .B(T5838_Y), .A(T11378_Y), .Y(T4388_Y));
KC_NAND2_X2 T4389 ( .B(T3794_Y), .A(T5800_Y), .Y(T4389_Y));
KC_NAND2_X2 T4392 ( .B(T11389_Y), .A(T5763_Y), .Y(T4392_Y));
KC_NAND2_X2 T4393 ( .B(T4394_Y), .A(T11365_Y), .Y(T4393_Y));
KC_NAND2_X2 T4394 ( .B(T5838_Y), .A(T16153_Y), .Y(T4394_Y));
KC_NAND2_X2 T4403 ( .B(T15907_Y), .A(T14942_Q), .Y(T4403_Y));
KC_NAND2_X2 T4431 ( .B(T4452_Y), .A(T3825_Y), .Y(T4431_Y));
KC_NAND2_X2 T4432 ( .B(T4478_Y), .A(T15907_Y), .Y(T4432_Y));
KC_NAND2_X2 T4436 ( .B(T5821_Y), .A(T5823_Y), .Y(T4436_Y));
KC_NAND2_X2 T4437 ( .B(T11370_Y), .A(T14546_Q), .Y(T4437_Y));
KC_NAND2_X2 T4438 ( .B(T4394_Y), .A(T3826_Y), .Y(T4438_Y));
KC_NAND2_X2 T4439 ( .B(T16153_Y), .A(T4463_Y), .Y(T4439_Y));
KC_NAND2_X2 T4440 ( .B(T4439_Y), .A(T4487_Q), .Y(T4440_Y));
KC_NAND2_X2 T4441 ( .B(T5826_Y), .A(T5821_Y), .Y(T4441_Y));
KC_NAND2_X2 T4445 ( .B(T4457_Y), .A(T15908_Y), .Y(T4445_Y));
KC_NAND2_X2 T4446 ( .B(T3856_Y), .A(T5815_Y), .Y(T4446_Y));
KC_NAND2_X2 T4448 ( .B(T11365_Y), .A(T4500_Y), .Y(T4448_Y));
KC_NAND2_X2 T4452 ( .B(T3856_Y), .A(T15908_Y), .Y(T4452_Y));
KC_NAND2_X2 T4471 ( .B(T4560_Y), .A(T4474_Y), .Y(T4471_Y));
KC_NAND2_X2 T4478 ( .B(T14549_Q), .A(T14548_Q), .Y(T4478_Y));
KC_NAND2_X2 T4481 ( .B(T5930_Y), .A(T4477_Y), .Y(T4481_Y));
KC_NAND2_X2 T4506 ( .B(T5929_Y), .A(T4489_Y), .Y(T4506_Y));
KC_NAND2_X2 T4507 ( .B(T3901_Y), .A(T12355_Y), .Y(T4507_Y));
KC_NAND2_X2 T4508 ( .B(T10629_Y), .A(T4482_Y), .Y(T4508_Y));
KC_NAND2_X2 T4510 ( .B(T5140_Y), .A(T4528_Q), .Y(T4510_Y));
KC_NAND2_X2 T4515 ( .B(T4482_Y), .A(T4518_Y), .Y(T4515_Y));
KC_NAND2_X2 T4516 ( .B(T4489_Y), .A(T4535_Y), .Y(T4516_Y));
KC_NAND2_X2 T4519 ( .B(T4527_Q), .A(T4526_Q), .Y(T4519_Y));
KC_NAND2_X2 T4520 ( .B(T5139_Y), .A(T4532_Y), .Y(T4520_Y));
KC_NAND2_X2 T4544 ( .B(T4575_Q), .A(T4572_Q), .Y(T4544_Y));
KC_NAND2_X2 T4545 ( .B(T5952_Y), .A(T11541_Y), .Y(T4545_Y));
KC_NAND2_X2 T4549 ( .B(T11542_Y), .A(T11538_Y), .Y(T4549_Y));
KC_NAND2_X2 T4550 ( .B(T4560_Y), .A(T4559_Y), .Y(T4550_Y));
KC_NAND2_X2 T4553 ( .B(T15592_Y), .A(T11555_Y), .Y(T4553_Y));
KC_NAND2_X2 T4556 ( .B(T4576_Q), .A(T4578_Q), .Y(T4556_Y));
KC_NAND2_X2 T4557 ( .B(T4588_Y), .A(T2073_Y), .Y(T4557_Y));
KC_NAND2_X2 T4558 ( .B(T4557_Y), .A(T5946_Y), .Y(T4558_Y));
KC_NAND2_X2 T4580 ( .B(T6021_Y), .A(T6344_Y), .Y(T4580_Y));
KC_NAND2_X2 T4581 ( .B(T6021_Y), .A(T4607_Q), .Y(T4581_Y));
KC_NAND2_X2 T4582 ( .B(T4597_Y), .A(T4621_Y), .Y(T4582_Y));
KC_NAND2_X2 T4595 ( .B(T11607_Y), .A(T11608_Y), .Y(T4595_Y));
KC_NAND2_X2 T4596 ( .B(T4607_Q), .A(T4608_Q), .Y(T4596_Y));
KC_NAND2_X2 T16047 ( .B(T4634_Y), .A(T4726_Y), .Y(T16047_Y));
KC_NAND2_X2 T4631 ( .B(T5145_Y), .A(T6467_Y), .Y(T4631_Y));
KC_NAND2_X2 T4632 ( .B(T4694_Y), .A(T6448_Y), .Y(T4632_Y));
KC_NAND2_X2 T4633 ( .B(T5152_Y), .A(T6448_Y), .Y(T4633_Y));
KC_NAND2_X2 T4634 ( .B(T5145_Y), .A(T6448_Y), .Y(T4634_Y));
KC_NAND2_X2 T4635 ( .B(T4694_Y), .A(T6467_Y), .Y(T4635_Y));
KC_NAND2_X2 T4636 ( .B(T5152_Y), .A(T6467_Y), .Y(T4636_Y));
KC_NAND2_X2 T4637 ( .B(T4635_Y), .A(T4725_Y), .Y(T4637_Y));
KC_NAND2_X2 T4639 ( .B(T6166_Y), .A(T4664_Y), .Y(T4639_Y));
KC_NAND2_X2 T4640 ( .B(T4632_Y), .A(T12855_Y), .Y(T4640_Y));
KC_NAND2_X2 T4642 ( .B(T12031_Y), .A(T8460_Y), .Y(T4642_Y));
KC_NAND2_X2 T4643 ( .B(T4664_Y), .A(T4725_Y), .Y(T4643_Y));
KC_NAND2_X2 T4644 ( .B(T8460_Y), .A(T12034_Y), .Y(T4644_Y));
KC_NAND2_X2 T4645 ( .B(T4726_Y), .A(T4632_Y), .Y(T4645_Y));
KC_NAND2_X2 T4646 ( .B(T4631_Y), .A(T4725_Y), .Y(T4646_Y));
KC_NAND2_X2 T4647 ( .B(T8459_Y), .A(T12034_Y), .Y(T4647_Y));
KC_NAND2_X2 T4648 ( .B(T12031_Y), .A(T8459_Y), .Y(T4648_Y));
KC_NAND2_X2 T4652 ( .B(T4636_Y), .A(T4725_Y), .Y(T4652_Y));
KC_NAND2_X2 T4653 ( .B(T8458_Y), .A(T12034_Y), .Y(T4653_Y));
KC_NAND2_X2 T4654 ( .B(T4633_Y), .A(T12855_Y), .Y(T4654_Y));
KC_NAND2_X2 T4655 ( .B(T12034_Y), .A(T8461_Y), .Y(T4655_Y));
KC_NAND2_X2 T4656 ( .B(T8462_Y), .A(T12034_Y), .Y(T4656_Y));
KC_NAND2_X2 T4657 ( .B(T4633_Y), .A(T4726_Y), .Y(T4657_Y));
KC_NAND2_X2 T4658 ( .B(T4634_Y), .A(T12855_Y), .Y(T4658_Y));
KC_NAND2_X2 T4659 ( .B(T8456_Y), .A(T12034_Y), .Y(T4659_Y));
KC_NAND2_X2 T4660 ( .B(T12031_Y), .A(T8456_Y), .Y(T4660_Y));
KC_NAND2_X2 T4694 ( .B(T4717_Q), .A(T4713_Q), .Y(T4694_Y));
KC_NAND2_X2 T4698 ( .B(T4071_Y), .A(T4691_Y), .Y(T4698_Y));
KC_NAND2_X2 T4700 ( .B(T11707_Y), .A(T10601_Y), .Y(T4700_Y));
KC_NAND2_X2 T4703 ( .B(T5144_Y), .A(T4706_Y), .Y(T4703_Y));
KC_NAND2_X2 T4706 ( .B(T10576_Y), .A(T6090_Y), .Y(T4706_Y));
KC_NAND2_X2 T4729 ( .B(T4706_Y), .A(T4733_Y), .Y(T4729_Y));
KC_NAND2_X2 T4731 ( .B(T6203_Y), .A(T15629_Y), .Y(T4731_Y));
KC_NAND2_X2 T4732 ( .B(T4742_Y), .A(T4752_Y), .Y(T4732_Y));
KC_NAND2_X2 T4733 ( .B(T4732_Y), .A(T15255_Y), .Y(T4733_Y));
KC_NAND2_X2 T4738 ( .B(T4740_Y), .A(T4743_Y), .Y(T4738_Y));
KC_NAND2_X2 T4762 ( .B(T16146_Y), .A(T15949_Y), .Y(T4762_Y));
KC_NAND2_X2 T4763 ( .B(T16146_Y), .A(T15687_Y), .Y(T4763_Y));
KC_NAND2_X2 T4764 ( .B(T16146_Y), .A(T4792_Y), .Y(T4764_Y));
KC_NAND2_X2 T4765 ( .B(T16146_Y), .A(T298_Y), .Y(T4765_Y));
KC_NAND2_X2 T4766 ( .B(T16146_Y), .A(T4791_Y), .Y(T4766_Y));
KC_NAND2_X2 T4767 ( .B(T16146_Y), .A(T4795_Y), .Y(T4767_Y));
KC_NAND2_X2 T4768 ( .B(T16146_Y), .A(T4794_Y), .Y(T4768_Y));
KC_NAND2_X2 T4769 ( .B(T16146_Y), .A(T4793_Y), .Y(T4769_Y));
KC_NAND2_X2 T4770 ( .B(T16146_Y), .A(T4789_Y), .Y(T4770_Y));
KC_NAND2_X2 T4771 ( .B(T16146_Y), .A(T4785_Y), .Y(T4771_Y));
KC_NAND2_X2 T4772 ( .B(T16146_Y), .A(T4790_Y), .Y(T4772_Y));
KC_NAND2_X2 T4773 ( .B(T16146_Y), .A(T4786_Y), .Y(T4773_Y));
KC_NAND2_X2 T4774 ( .B(T16146_Y), .A(T4780_Y), .Y(T4774_Y));
KC_NAND2_X2 T4775 ( .B(T16146_Y), .A(T4779_Y), .Y(T4775_Y));
KC_NAND2_X2 T4776 ( .B(T16146_Y), .A(T4778_Y), .Y(T4776_Y));
KC_NAND2_X2 T4777 ( .B(T16146_Y), .A(T4781_Y), .Y(T4777_Y));
KC_NAND2_X2 T9454 ( .B(T9453_Y), .A(T9013_Y), .Y(T9454_Y));
KC_NAND2_X2 T9453 ( .B(T11296_Y), .A(T9089_Y), .Y(T9453_Y));
KC_NAND2_X2 T9450 ( .B(T9093_Y), .A(T9079_Y), .Y(T9450_Y));
KC_NAND2_X2 T9389 ( .B(T917_Y), .A(T7826_Y), .Y(T9389_Y));
KC_NAND2_X2 T9388 ( .B(T16332_Y), .A(T382_Y), .Y(T9388_Y));
KC_NAND2_X2 T16189 ( .B(T15538_Y), .A(T4842_Y), .Y(T16189_Y));
KC_NAND2_X2 T9478 ( .B(T15538_Y), .A(T15540_Y), .Y(T9478_Y));
KC_NAND2_X2 T9446 ( .B(T605_Q), .A(T15795_Q), .Y(T9446_Y));
KC_NAND2_X2 T9438 ( .B(T10941_Y), .A(T9432_Y), .Y(T9438_Y));
KC_NAND2_X2 T9437 ( .B(T16274_Y), .A(T9031_Y), .Y(T9437_Y));
KC_NAND2_X2 T9436 ( .B(T9432_Y), .A(T4872_Y), .Y(T9436_Y));
KC_NAND2_X2 T9374 ( .B(T786_Y), .A(T8757_Y), .Y(T9374_Y));
KC_NAND2_X2 T9373 ( .B(T902_Y), .A(T8757_Y), .Y(T9373_Y));
KC_NAND2_X2 T9370 ( .B(T8757_Y), .A(T8829_Y), .Y(T9370_Y));
KC_NAND2_X2 T9331 ( .B(T637_Y), .A(T8682_Y), .Y(T9331_Y));
KC_NAND2_X2 T10345 ( .B(T4858_Q), .A(T15665_Y), .Y(T10345_Y));
KC_NAND2_X2 T10344 ( .B(T1037_Q), .A(T15751_Y), .Y(T10344_Y));
KC_NAND2_X2 T10303 ( .B(T10161_Y), .A(T16275_Y), .Y(T10303_Y));
KC_NAND2_X2 T9405 ( .B(T7949_Y), .A(T16384_Y), .Y(T9405_Y));
KC_NAND2_X2 T9332 ( .B(T1066_Q), .A(T656_Y), .Y(T9332_Y));
KC_NAND2_X2 T4865 ( .B(T1275_Y), .A(T5382_Y), .Y(T4865_Y));
KC_NAND2_X2 T10308 ( .B(T10032_Y), .A(T15087_Y), .Y(T10308_Y));
KC_NAND2_X2 T4905 ( .B(T10525_Y), .A(T16433_Q), .Y(T4905_Y));
KC_NAND2_X2 T4912 ( .B(T10627_Y), .A(T2279_Y), .Y(T4912_Y));
KC_NAND2_X2 T16267 ( .B(T10880_Y), .A(T13131_Y), .Y(T16267_Y));
KC_NAND2_X2 T4933 ( .B(T4934_Y), .A(T2040_Y), .Y(T4933_Y));
KC_NAND2_X2 T4934 ( .B(T10100_Y), .A(T5367_Y), .Y(T4934_Y));
KC_NAND2_X2 T4935 ( .B(T16371_Y), .A(T2604_Y), .Y(T4935_Y));
KC_NAND2_X2 T4942 ( .B(T11499_Y), .A(T11639_Y), .Y(T4942_Y));
KC_NAND2_X2 T4943 ( .B(T15942_Y), .A(T16010_Q), .Y(T4943_Y));
KC_NAND2_X2 T4946 ( .B(T6464_Y), .A(T16082_Q), .Y(T4946_Y));
KC_NAND2_X2 T4954 ( .B(T6003_Y), .A(T12106_Y), .Y(T4954_Y));
KC_NAND2_X2 T16265 ( .B(T10184_Y), .A(T16264_Y), .Y(T16265_Y));
KC_NAND2_X2 T16262 ( .B(T3177_Y), .A(T14995_Y), .Y(T16262_Y));
KC_NAND2_X2 T4981 ( .B(T10540_Y), .A(T12148_Y), .Y(T4981_Y));
KC_NAND2_X2 T4982 ( .B(T5024_Y), .A(T10518_Y), .Y(T4982_Y));
KC_NAND2_X2 T4984 ( .B(T1132_Y), .A(T16275_Y), .Y(T4984_Y));
KC_NAND2_X2 T4985 ( .B(T9854_Y), .A(T9747_Y), .Y(T4985_Y));
KC_NAND2_X2 T4986 ( .B(T13960_Q), .A(T16079_Q), .Y(T4986_Y));
KC_NAND2_X2 T4991 ( .B(T15943_Y), .A(T2848_Y), .Y(T4991_Y));
KC_NAND2_X2 T4992 ( .B(T15696_Y), .A(T5749_Y), .Y(T4992_Y));
KC_NAND2_X2 T4993 ( .B(T10269_Y), .A(T6729_Y), .Y(T4993_Y));
KC_NAND2_X2 T4994 ( .B(T4995_Y), .A(T10279_Y), .Y(T4994_Y));
KC_NAND2_X2 T4995 ( .B(T5714_Y), .A(T10278_Y), .Y(T4995_Y));
KC_NAND2_X2 T4998 ( .B(T6576_Y), .A(T15762_Y), .Y(T4998_Y));
KC_NAND2_X2 T4999 ( .B(T6101_Y), .A(T15712_Y), .Y(T4999_Y));
KC_NAND2_X2 T5002 ( .B(T11831_Y), .A(T2874_Q), .Y(T5002_Y));
KC_NAND2_X2 T5003 ( .B(T6160_Y), .A(T16101_Y), .Y(T5003_Y));
KC_NAND2_X2 T5008 ( .B(T2276_Q), .A(T2854_Y), .Y(T5008_Y));
KC_NAND2_X2 T5037 ( .B(T14984_Y), .A(T3544_Y), .Y(T5037_Y));
KC_NAND2_X2 T5038 ( .B(T14984_Y), .A(T2966_Y), .Y(T5038_Y));
KC_NAND2_X2 T5039 ( .B(T15699_Y), .A(T15863_Y), .Y(T5039_Y));
KC_NAND2_X2 T5042 ( .B(T5043_Y), .A(T3920_Y), .Y(T5042_Y));
KC_NAND2_X2 T5045 ( .B(T15616_Y), .A(T16102_Y), .Y(T5045_Y));
KC_NAND2_X2 T5046 ( .B(T10545_Y), .A(T3447_Y), .Y(T5046_Y));
KC_NAND2_X2 T5047 ( .B(T10568_Y), .A(T10545_Y), .Y(T5047_Y));
KC_NAND2_X2 T5048 ( .B(T15616_Y), .A(T11818_Y), .Y(T5048_Y));
KC_NAND2_X2 T5049 ( .B(T15711_Y), .A(T15616_Y), .Y(T5049_Y));
KC_NAND2_X2 T5050 ( .B(T10968_Y), .A(T16149_Y), .Y(T5050_Y));
KC_NAND2_X2 T5051 ( .B(T3362_Y), .A(T6138_Y), .Y(T5051_Y));
KC_NAND2_X2 T5052 ( .B(T5523_Y), .A(T10623_Y), .Y(T5052_Y));
KC_NAND2_X2 T5056 ( .B(T15233_Y), .A(T11641_Y), .Y(T5056_Y));
KC_NAND2_X2 T5058 ( .B(T3413_Y), .A(T6048_Y), .Y(T5058_Y));
KC_NAND2_X2 T5059 ( .B(T16034_Y), .A(T10584_Y), .Y(T5059_Y));
KC_NAND2_X2 T5082 ( .B(T6802_Y), .A(T6839_Y), .Y(T5082_Y));
KC_NAND2_X2 T5099 ( .B(T12227_Y), .A(T5989_Y), .Y(T5099_Y));
KC_NAND2_X2 T5101 ( .B(T5788_Y), .A(T11428_Y), .Y(T5101_Y));
KC_NAND2_X2 T5105 ( .B(T11365_Y), .A(T5763_Y), .Y(T5105_Y));
KC_NAND2_X2 T5111 ( .B(T3397_Y), .A(T16140_Y), .Y(T5111_Y));
KC_NAND2_X2 T5112 ( .B(T6000_Y), .A(T4066_Y), .Y(T5112_Y));
KC_NAND2_X2 T16251 ( .B(T15441_Y), .A(T7707_Y), .Y(T16251_Y));
KC_NAND2_X2 T16250 ( .B(T7707_Y), .A(T3073_Y), .Y(T16250_Y));
KC_NAND2_X2 T16248 ( .B(T12761_Y), .A(T10115_Y), .Y(T16248_Y));
KC_NAND2_X2 T5139 ( .B(T4532_Y), .A(T12024_Y), .Y(T5139_Y));
KC_NAND2_X2 T5144 ( .B(T15756_Y), .A(T16144_Y), .Y(T5144_Y));
KC_NAND2_X2 T5145 ( .B(T6171_Y), .A(T4717_Q), .Y(T5145_Y));
KC_NAND2_X2 T5634 ( .B(T83_Q), .A(T5185_Q), .Y(T5634_Y));
KC_NAND2_X2 T5617 ( .B(T16479_Y), .A(T8543_Y), .Y(T5617_Y));
KC_NAND2_X2 T9317 ( .B(T7599_Y), .A(T8758_Y), .Y(T9317_Y));
KC_NAND2_X2 T7542 ( .B(T15393_Y), .A(T1476_Y), .Y(T7542_Y));
KC_NAND2_X2 T7490 ( .B(T1476_Y), .A(T7703_Y), .Y(T7490_Y));
KC_NAND2_X2 T7685 ( .B(T928_Y), .A(T8771_Y), .Y(T7685_Y));
KC_NAND2_X2 T7636 ( .B(T15223_Y), .A(T927_Y), .Y(T7636_Y));
KC_NAND2_X2 T5288 ( .B(T3110_Y), .A(T14995_Y), .Y(T5288_Y));
KC_NAND2_X2 T7826 ( .B(T612_Y), .A(T8776_Y), .Y(T7826_Y));
KC_NAND2_X2 T7820 ( .B(T15084_Y), .A(T8777_Y), .Y(T7820_Y));
KC_NAND2_X2 T5330 ( .B(T14995_Y), .A(T3108_Y), .Y(T5330_Y));
KC_NAND2_X2 T9008 ( .B(T762_Q), .A(T9002_Y), .Y(T9008_Y));
KC_NAND2_X2 T8079 ( .B(T613_Y), .A(T8963_Y), .Y(T8079_Y));
KC_NAND2_X2 T8062 ( .B(T16311_Y), .A(T1349_Y), .Y(T8062_Y));
KC_NAND2_X2 T5369 ( .B(T1518_Y), .A(T10526_Y), .Y(T5369_Y));
KC_NAND2_X2 T9182 ( .B(T9180_Y), .A(T15150_Y), .Y(T9182_Y));
KC_NAND2_X2 T15852 ( .B(T8175_Y), .A(T8174_Y), .Y(T15852_Y));
KC_NAND2_X2 T5427 ( .B(T5766_Y), .A(T10241_Y), .Y(T5427_Y));
KC_NAND2_X2 T5436 ( .B(T15942_Y), .A(T5987_Q), .Y(T5436_Y));
KC_NAND2_X2 T5448 ( .B(T3896_Y), .A(T4505_Y), .Y(T5448_Y));
KC_NAND2_X2 T5457 ( .B(T4508_Y), .A(T4515_Y), .Y(T5457_Y));
KC_NAND2_X2 T5458 ( .B(T5914_Y), .A(T11505_Y), .Y(T5458_Y));
KC_NAND2_X2 T5459 ( .B(T11523_Y), .A(T10632_Y), .Y(T5459_Y));
KC_NAND2_X2 T5468 ( .B(T5972_Y), .A(T5860_Y), .Y(T5468_Y));
KC_NAND2_X2 T5517 ( .B(T6225_Y), .A(T12103_Y), .Y(T5517_Y));
KC_NAND2_X2 T5520 ( .B(T6240_Y), .A(T2329_Y), .Y(T5520_Y));
KC_NAND2_X2 T5521 ( .B(T6513_Y), .A(T11742_Y), .Y(T5521_Y));
KC_NAND2_X2 T5522 ( .B(T11815_Y), .A(T11822_Y), .Y(T5522_Y));
KC_NAND2_X2 T5533 ( .B(T15640_Y), .A(T11813_Y), .Y(T5533_Y));
KC_NAND2_X2 T9399 ( .B(T9414_Y), .A(T7676_Y), .Y(T9399_Y));
KC_NAND2_X2 T5553 ( .B(T11367_Y), .A(T14550_Q), .Y(T5553_Y));
KC_NAND2_X2 T5556 ( .B(T16034_Y), .A(T11996_Y), .Y(T5556_Y));
KC_BUF_X5 T29 ( .Y(T29_Y), .A(T13068_Y));
KC_BUF_X5 T35 ( .Y(T35_Y), .A(T13075_Y));
KC_BUF_X5 T5593 ( .Y(T5593_Y), .A(T13075_Y));
KC_BUF_X5 T56 ( .Y(T56_Y), .A(T70_Y));
KC_BUF_X5 T82 ( .Y(T82_Y), .A(T70_Y));
KC_BUF_X5 T90 ( .Y(T90_Y), .A(T15321_Y));
KC_BUF_X5 T97 ( .Y(T97_Y), .A(T15321_Y));
KC_BUF_X5 T138 ( .Y(T138_Y), .A(T13288_Y));
KC_BUF_X5 T175 ( .Y(T175_Y), .A(T13288_Y));
KC_BUF_X5 T178 ( .Y(T178_Y), .A(T13935_Q));
KC_BUF_X5 T197 ( .Y(T197_Y), .A(T5423_Y));
KC_BUF_X5 T198 ( .Y(T198_Y), .A(T202_Y));
KC_BUF_X5 T280 ( .Y(T280_Y), .A(T293_Q));
KC_BUF_X5 T309 ( .Y(T309_Y), .A(T685_Y));
KC_BUF_X5 T352 ( .Y(T352_Y), .A(T14588_Q));
KC_BUF_X5 T400 ( .Y(T400_Y), .A(T1335_Y));
KC_BUF_X5 T428 ( .Y(T428_Y), .A(T16482_Q));
KC_BUF_X5 T429 ( .Y(T429_Y), .A(T15828_Q));
KC_BUF_X5 T433 ( .Y(T433_Y), .A(T6949_Y));
KC_BUF_X5 T465 ( .Y(T465_Y), .A(T15369_Y));
KC_BUF_X5 T466 ( .Y(T466_Y), .A(T15369_Y));
KC_BUF_X5 T495 ( .Y(T495_Y), .A(T685_Y));
KC_BUF_X5 T503 ( .Y(T503_Y), .A(T13933_Q));
KC_BUF_X5 T510 ( .Y(T510_Y), .A(T13932_Q));
KC_BUF_X5 T575 ( .Y(T575_Y), .A(T15484_Y));
KC_BUF_X5 T582 ( .Y(T582_Y), .A(T15484_Y));
KC_BUF_X5 T594 ( .Y(T594_Y), .A(T14452_Q));
KC_BUF_X5 T640 ( .Y(T640_Y), .A(T13932_Q));
KC_BUF_X5 T644 ( .Y(T644_Y), .A(T13933_Q));
KC_BUF_X5 T685 ( .Y(T685_Y), .A(T13934_Q));
KC_BUF_X5 T686 ( .Y(T686_Y), .A(T14097_Q));
KC_BUF_X5 T693 ( .Y(T693_Y), .A(T13935_Q));
KC_BUF_X5 T706 ( .Y(T706_Y), .A(T708_Y));
KC_BUF_X5 T707 ( .Y(T707_Y), .A(T5298_Y));
KC_BUF_X5 T708 ( .Y(T708_Y), .A(T707_Y));
KC_BUF_X5 T792 ( .Y(T792_Y), .A(T15335_Y));
KC_BUF_X5 T798 ( .Y(T798_Y), .A(T15335_Y));
KC_BUF_X5 T810 ( .Y(T810_Y), .A(T685_Y));
KC_BUF_X5 T836 ( .Y(T836_Y), .A(T8688_Y));
KC_BUF_X5 T846 ( .Y(T846_Y), .A(T14097_Q));
KC_BUF_X5 T855 ( .Y(T855_Y), .A(T685_Y));
KC_BUF_X5 T890 ( .Y(T890_Y), .A(T15411_Y));
KC_BUF_X5 T891 ( .Y(T891_Y), .A(T15411_Y));
KC_BUF_X5 T911 ( .Y(T911_Y), .A(T13262_Y));
KC_BUF_X5 T923 ( .Y(T923_Y), .A(T685_Y));
KC_BUF_X5 T958 ( .Y(T958_Y), .A(T12703_Y));
KC_BUF_X5 T971 ( .Y(T971_Y), .A(T16415_Y));
KC_BUF_X5 T990 ( .Y(T990_Y), .A(T14982_Y));
KC_BUF_X5 T991 ( .Y(T991_Y), .A(T990_Y));
KC_BUF_X5 T1023 ( .Y(T1023_Y), .A(T15951_Y));
KC_BUF_X5 T1030 ( .Y(T1030_Y), .A(T15673_Y));
KC_BUF_X5 T1047 ( .Y(T1047_Y), .A(T685_Y));
KC_BUF_X5 T1074 ( .Y(T1074_Y), .A(T14588_Q));
KC_BUF_X5 T1112 ( .Y(T1112_Y), .A(T1244_Y));
KC_BUF_X5 T1115 ( .Y(T1115_Y), .A(T14588_Q));
KC_BUF_X5 T1120 ( .Y(T1120_Y), .A(T14588_Q));
KC_BUF_X5 T1140 ( .Y(T1140_Y), .A(T991_Y));
KC_BUF_X5 T1145 ( .Y(T1145_Y), .A(T8189_Y));
KC_BUF_X5 T1147 ( .Y(T1147_Y), .A(T943_Y));
KC_BUF_X5 T1163 ( .Y(T1163_Y), .A(T1147_Y));
KC_BUF_X5 T1229 ( .Y(T1229_Y), .A(T15496_Y));
KC_BUF_X5 T1240 ( .Y(T1240_Y), .A(T15496_Y));
KC_BUF_X5 T1243 ( .Y(T1243_Y), .A(T5480_Q));
KC_BUF_X5 T1318 ( .Y(T1318_Y), .A(T15342_Y));
KC_BUF_X5 T1325 ( .Y(T1325_Y), .A(T1403_Y));
KC_BUF_X5 T1356 ( .Y(T1356_Y), .A(T14983_Y));
KC_BUF_X5 T1363 ( .Y(T1363_Y), .A(T4902_Y));
KC_BUF_X5 T1373 ( .Y(T1373_Y), .A(T5413_Y));
KC_BUF_X5 T1374 ( .Y(T1374_Y), .A(T1373_Y));
KC_BUF_X5 T1376 ( .Y(T1376_Y), .A(T1381_Y));
KC_BUF_X5 T1381 ( .Y(T1381_Y), .A(T1382_Y));
KC_BUF_X5 T1382 ( .Y(T1382_Y), .A(T4881_Y));
KC_BUF_X5 T1384 ( .Y(T1384_Y), .A(T13057_Q));
KC_BUF_X5 T1385 ( .Y(T1385_Y), .A(T4882_Y));
KC_BUF_X5 T1390 ( .Y(T1390_Y), .A(T15342_Y));
KC_BUF_X5 T1403 ( .Y(T1403_Y), .A(T2059_Y));
KC_BUF_X5 T1463 ( .Y(T1463_Y), .A(T15415_Y));
KC_BUF_X5 T1464 ( .Y(T1464_Y), .A(T15415_Y));
KC_BUF_X5 T1510 ( .Y(T1510_Y), .A(T4897_Y));
KC_BUF_X5 T1514 ( .Y(T1514_Y), .A(T1516_Y));
KC_BUF_X5 T1515 ( .Y(T1515_Y), .A(T1514_Y));
KC_BUF_X5 T1516 ( .Y(T1516_Y), .A(T1613_Y));
KC_BUF_X5 T1525 ( .Y(T1525_Y), .A(T2059_Y));
KC_BUF_X5 T1534 ( .Y(T1534_Y), .A(T8671_Y));
KC_BUF_X5 T1540 ( .Y(T1540_Y), .A(T8671_Y));
KC_BUF_X5 T1549 ( .Y(T1549_Y), .A(T1964_Y));
KC_BUF_X5 T1560 ( .Y(T1560_Y), .A(T2059_Y));
KC_BUF_X5 T1569 ( .Y(T1569_Y), .A(T11279_Y));
KC_BUF_X5 T1589 ( .Y(T1589_Y), .A(T2011_Y));
KC_BUF_X5 T1598 ( .Y(T1598_Y), .A(T15176_Y));
KC_BUF_X5 T1600 ( .Y(T1600_Y), .A(T1601_Y));
KC_BUF_X5 T1601 ( .Y(T1601_Y), .A(T5371_Y));
KC_BUF_X5 T1604 ( .Y(T1604_Y), .A(T1600_Y));
KC_BUF_X5 T1608 ( .Y(T1608_Y), .A(T1609_Y));
KC_BUF_X5 T1609 ( .Y(T1609_Y), .A(T15168_Q));
KC_BUF_X5 T1610 ( .Y(T1610_Y), .A(T1615_Y));
KC_BUF_X5 T1611 ( .Y(T1611_Y), .A(T1610_Y));
KC_BUF_X5 T1612 ( .Y(T1612_Y), .A(T1611_Y));
KC_BUF_X5 T1613 ( .Y(T1613_Y), .A(T1612_Y));
KC_BUF_X5 T1614 ( .Y(T1614_Y), .A(T1740_Y));
KC_BUF_X5 T1615 ( .Y(T1615_Y), .A(T1614_Y));
KC_BUF_X5 T1638 ( .Y(T1638_Y), .A(T1964_Y));
KC_BUF_X5 T1650 ( .Y(T1650_Y), .A(T1964_Y));
KC_BUF_X5 T1651 ( .Y(T1651_Y), .A(T1964_Y));
KC_BUF_X5 T1722 ( .Y(T1722_Y), .A(T14998_Y));
KC_BUF_X5 T1740 ( .Y(T1740_Y), .A(T1608_Y));
KC_BUF_X5 T1747 ( .Y(T1747_Y), .A(T13102_Q));
KC_BUF_X5 T1754 ( .Y(T1754_Y), .A(T4924_Q));
KC_BUF_X5 T1824 ( .Y(T1824_Y), .A(T5513_Q));
KC_BUF_X5 T1862 ( .Y(T1862_Y), .A(T15347_Y));
KC_BUF_X5 T1866 ( .Y(T1866_Y), .A(T15347_Y));
KC_BUF_X5 T1963 ( .Y(T1963_Y), .A(T2059_Y));
KC_BUF_X5 T1964 ( .Y(T1964_Y), .A(T14368_Q));
KC_BUF_X5 T1965 ( .Y(T1965_Y), .A(T6848_Y));
KC_BUF_X5 T2007 ( .Y(T2007_Y), .A(T15843_Y));
KC_BUF_X5 T2013 ( .Y(T2013_Y), .A(T10083_Y));
KC_BUF_X5 T2027 ( .Y(T2027_Y), .A(T16193_Y));
KC_BUF_X5 T2047 ( .Y(T2047_Y), .A(T1964_Y));
KC_BUF_X5 T2050 ( .Y(T2050_Y), .A(T16253_Y));
KC_BUF_X5 T2058 ( .Y(T2058_Y), .A(T15511_Y));
KC_BUF_X5 T2059 ( .Y(T2059_Y), .A(T13266_Y));
KC_BUF_X5 T2075 ( .Y(T2075_Y), .A(T1984_Q));
KC_BUF_X5 T2078 ( .Y(T2078_Y), .A(T1356_Y));
KC_BUF_X5 T2083 ( .Y(T2083_Y), .A(T13266_Y));
KC_BUF_X5 T2097 ( .Y(T2097_Y), .A(T15191_Q));
KC_BUF_X5 T2124 ( .Y(T2124_Y), .A(T2766_Y));
KC_BUF_X5 T2131 ( .Y(T2131_Y), .A(T2097_Y));
KC_BUF_X5 T2156 ( .Y(T2156_Y), .A(T2131_Y));
KC_BUF_X5 T2342 ( .Y(T2342_Y), .A(T15990_Q));
KC_BUF_X5 T2343 ( .Y(T2343_Y), .A(T15038_Y));
KC_BUF_X5 T2349 ( .Y(T2349_Y), .A(T11783_Y));
KC_BUF_X5 T2350 ( .Y(T2350_Y), .A(T2250_Y));
KC_BUF_X5 T2377 ( .Y(T2377_Y), .A(T2377_A));
KC_BUF_X5 T2378 ( .Y(T2378_Y), .A(T2378_A));
KC_BUF_X5 T2384 ( .Y(T2384_Y), .A(T16023_Q));
KC_BUF_X5 T2441 ( .Y(T2441_Y), .A(T15381_Y));
KC_BUF_X5 T2443 ( .Y(T2443_Y), .A(T15381_Y));
KC_BUF_X5 T2488 ( .Y(T2488_Y), .A(T11278_Y));
KC_BUF_X5 T2495 ( .Y(T2495_Y), .A(T1964_Y));
KC_BUF_X5 T2529 ( .Y(T2529_Y), .A(T13012_Q));
KC_BUF_X5 T2589 ( .Y(T2589_Y), .A(T10194_Y));
KC_BUF_X5 T2667 ( .Y(T2667_Y), .A(T16446_Q));
KC_BUF_X5 T2736 ( .Y(T2736_Y), .A(T2157_Y));
KC_BUF_X5 T2744 ( .Y(T2744_Y), .A(T11463_Y));
KC_BUF_X5 T2753 ( .Y(T2753_Y), .A(T10640_Y));
KC_BUF_X5 T2789 ( .Y(T2789_Y), .A(T15991_Y));
KC_BUF_X5 T2790 ( .Y(T2790_Y), .A(T2736_Y));
KC_BUF_X5 T2791 ( .Y(T2791_Y), .A(T3876_Y));
KC_BUF_X5 T2811 ( .Y(T2811_Y), .A(T5570_Y));
KC_BUF_X5 T2813 ( .Y(T2813_Y), .A(T16134_Y));
KC_BUF_X5 T2871 ( .Y(T2871_Y), .A(T13142_Y));
KC_BUF_X5 T3026 ( .Y(T3026_Y), .A(T1964_Y));
KC_BUF_X5 T3061 ( .Y(T3061_Y), .A(T9739_Y));
KC_BUF_X5 T3075 ( .Y(T3075_Y), .A(T5715_Y));
KC_BUF_X5 T3122 ( .Y(T3122_Y), .A(T1964_Y));
KC_BUF_X5 T3153 ( .Y(T3153_Y), .A(T2623_Y));
KC_BUF_X5 T3158 ( .Y(T3158_Y), .A(T16303_Y));
KC_BUF_X5 T3188 ( .Y(T3188_Y), .A(T15551_Y));
KC_BUF_X5 T3191 ( .Y(T3191_Y), .A(T15551_Y));
KC_BUF_X5 T3198 ( .Y(T3198_Y), .A(T14953_Q));
KC_BUF_X5 T3199 ( .Y(T3199_Y), .A(T14953_Q));
KC_BUF_X5 T3209 ( .Y(T3209_Y), .A(T3217_Y));
KC_BUF_X5 T3215 ( .Y(T3215_Y), .A(T3216_Y));
KC_BUF_X5 T3216 ( .Y(T3216_Y), .A(T4897_Y));
KC_BUF_X5 T3234 ( .Y(T3234_Y), .A(T15565_Y));
KC_BUF_X5 T3239 ( .Y(T3239_Y), .A(T15565_Y));
KC_BUF_X5 T3254 ( .Y(T3254_Y), .A(T11457_Y));
KC_BUF_X5 T3263 ( .Y(T3263_Y), .A(T3315_Y));
KC_BUF_X5 T3264 ( .Y(T3264_Y), .A(T14556_Q));
KC_BUF_X5 T3279 ( .Y(T3279_Y), .A(T15182_Q));
KC_BUF_X5 T3282 ( .Y(T3282_Y), .A(T2127_Y));
KC_BUF_X5 T3307 ( .Y(T3307_Y), .A(T2761_Y));
KC_BUF_X5 T3311 ( .Y(T3311_Y), .A(T3991_Y));
KC_BUF_X5 T3314 ( .Y(T3314_Y), .A(T10638_Y));
KC_BUF_X5 T3316 ( .Y(T3316_Y), .A(T11477_Y));
KC_BUF_X5 T3332 ( .Y(T3332_Y), .A(T11561_Y));
KC_BUF_X5 T3333 ( .Y(T3333_Y), .A(T16202_Y));
KC_BUF_X5 T3340 ( .Y(T3340_Y), .A(T3291_Y));
KC_BUF_X5 T3414 ( .Y(T3414_Y), .A(T3403_Y));
KC_BUF_X5 T3496 ( .Y(T3496_Y), .A(T14963_Q));
KC_BUF_X5 T3584 ( .Y(T3584_Y), .A(T2059_Y));
KC_BUF_X5 T3638 ( .Y(T3638_Y), .A(T3290_Y));
KC_BUF_X5 T3643 ( .Y(T3643_Y), .A(T3290_Y));
KC_BUF_X5 T3681 ( .Y(T3681_Y), .A(T3658_Y));
KC_BUF_X5 T3879 ( .Y(T3879_Y), .A(T5351_Y));
KC_BUF_X5 T3934 ( .Y(T3934_Y), .A(T3933_Y));
KC_BUF_X5 T3938 ( .Y(T3938_Y), .A(T15594_Y));
KC_BUF_X5 T3939 ( .Y(T3939_Y), .A(T4174_Y));
KC_BUF_X5 T3957 ( .Y(T3957_Y), .A(T15594_Y));
KC_BUF_X5 T3993 ( .Y(T3993_Y), .A(T14556_Q));
KC_BUF_X5 T3994 ( .Y(T3994_Y), .A(T5501_Q));
KC_BUF_X5 T3995 ( .Y(T3995_Y), .A(T4056_Q));
KC_BUF_X5 T3999 ( .Y(T3999_Y), .A(T2809_Q));
KC_BUF_X5 T4000 ( .Y(T4000_Y), .A(T5499_Q));
KC_BUF_X5 T4001 ( .Y(T4001_Y), .A(T4714_Q));
KC_BUF_X5 T4002 ( .Y(T4002_Y), .A(T5502_Q));
KC_BUF_X5 T4003 ( .Y(T4003_Y), .A(T4663_Q));
KC_BUF_X5 T4004 ( .Y(T4004_Y), .A(T4675_Q));
KC_BUF_X5 T4005 ( .Y(T4005_Y), .A(T4043_Q));
KC_BUF_X5 T4012 ( .Y(T4012_Y), .A(T5496_Q));
KC_BUF_X5 T4013 ( .Y(T4013_Y), .A(T5498_Q));
KC_BUF_X5 T4014 ( .Y(T4014_Y), .A(T14959_Q));
KC_BUF_X5 T4039 ( .Y(T4039_Y), .A(T4352_Y));
KC_BUF_X5 T4045 ( .Y(T4045_Y), .A(T14963_Q));
KC_BUF_X5 T4047 ( .Y(T4047_Y), .A(T2081_Y));
KC_BUF_X5 T4175 ( .Y(T4175_Y), .A(T11659_Y));
KC_BUF_X5 T4190 ( .Y(T4190_Y), .A(T15366_Y));
KC_BUF_X5 T4191 ( .Y(T4191_Y), .A(T5552_Y));
KC_BUF_X5 T4198 ( .Y(T4198_Y), .A(T15366_Y));
KC_BUF_X5 T4227 ( .Y(T4227_Y), .A(T6455_Y));
KC_BUF_X5 T4282 ( .Y(T4282_Y), .A(T4897_Y));
KC_BUF_X5 T4331 ( .Y(T4331_Y), .A(T2724_Y));
KC_BUF_X5 T4332 ( .Y(T4332_Y), .A(T2724_Y));
KC_BUF_X5 T4350 ( .Y(T4350_Y), .A(T16253_Y));
KC_BUF_X5 T4501 ( .Y(T4501_Y), .A(T15557_Y));
KC_BUF_X5 T4502 ( .Y(T4502_Y), .A(T11443_Y));
KC_BUF_X5 T4524 ( .Y(T4524_Y), .A(T12207_Y));
KC_BUF_X5 T4531 ( .Y(T4531_Y), .A(T16152_Y));
KC_BUF_X5 T4542 ( .Y(T4542_Y), .A(T3315_Y));
KC_BUF_X5 T4570 ( .Y(T4570_Y), .A(T3334_Y));
KC_BUF_X5 T4601 ( .Y(T4601_Y), .A(T4580_Y));
KC_BUF_X5 T4605 ( .Y(T4605_Y), .A(T2719_Y));
KC_BUF_X5 T4610 ( .Y(T4610_Y), .A(T4686_Q));
KC_BUF_X5 T4618 ( .Y(T4618_Y), .A(T4669_Q));
KC_BUF_X5 T4619 ( .Y(T4619_Y), .A(T4693_Q));
KC_BUF_X5 T4620 ( .Y(T4620_Y), .A(T4685_Q));
KC_BUF_X5 T4668 ( .Y(T4668_Y), .A(T11558_Y));
KC_BUF_X5 T4691 ( .Y(T4691_Y), .A(T13139_Y));
KC_BUF_X5 T4692 ( .Y(T4692_Y), .A(T16046_Y));
KC_BUF_X5 T4728 ( .Y(T4728_Y), .A(T14959_Q));
KC_BUF_X5 T4749 ( .Y(T4749_Y), .A(T4733_Y));
KC_BUF_X5 T4754 ( .Y(T4754_Y), .A(T286_Y));
KC_BUF_X5 T4782 ( .Y(T4782_Y), .A(T4186_Y));
KC_BUF_X5 T4798 ( .Y(T4798_Y), .A(T13068_Y));
KC_BUF_X5 T4812 ( .Y(T4812_Y), .A(T14097_Q));
KC_BUF_X5 T16190 ( .Y(T16190_Y), .A(T15540_Y));
KC_BUF_X5 T4826 ( .Y(T4826_Y), .A(T13288_Y));
KC_BUF_X5 T4828 ( .Y(T4828_Y), .A(T13288_Y));
KC_BUF_X5 T4849 ( .Y(T4849_Y), .A(T706_Y));
KC_BUF_X5 T4851 ( .Y(T4851_Y), .A(T14369_Q));
KC_BUF_X5 T4881 ( .Y(T4881_Y), .A(T1385_Y));
KC_BUF_X5 T4882 ( .Y(T4882_Y), .A(T13064_Q));
KC_BUF_X5 T4900 ( .Y(T4900_Y), .A(T1964_Y));
KC_BUF_X5 T4929 ( .Y(T4929_Y), .A(T16481_Q));
KC_BUF_X5 T4977 ( .Y(T4977_Y), .A(T1964_Y));
KC_BUF_X5 T4979 ( .Y(T4979_Y), .A(T5527_Q));
KC_BUF_X5 T5064 ( .Y(T5064_Y), .A(T16152_Y));
KC_BUF_X5 T5127 ( .Y(T5127_Y), .A(T4352_Y));
KC_BUF_X5 T5156 ( .Y(T5156_Y), .A(T4567_Y));
KC_BUF_X5 T5175 ( .Y(T5175_Y), .A(T6455_Y));
KC_BUF_X5 T5197 ( .Y(T5197_Y), .A(T13935_Q));
KC_BUF_X5 T5298 ( .Y(T5298_Y), .A(T911_Y));
KC_BUF_X5 T5315 ( .Y(T5315_Y), .A(T1964_Y));
KC_BUF_X5 T5361 ( .Y(T5361_Y), .A(T2059_Y));
KC_BUF_X5 T5371 ( .Y(T5371_Y), .A(T1722_Y));
KC_BUF_X5 T5413 ( .Y(T5413_Y), .A(T1376_Y));
KC_BUF_X5 T5422 ( .Y(T5422_Y), .A(T2089_Q));
KC_BUF_X5 T5482 ( .Y(T5482_Y), .A(T16049_Q));
KC_BUF_X5 T5485 ( .Y(T5485_Y), .A(T3997_Y));
KC_BUF_X5 T5531 ( .Y(T5531_Y), .A(T15639_Y));
KC_BUF_X5 T5542 ( .Y(T5542_Y), .A(T15639_Y));
KC_BUF_X5 T5557 ( .Y(T5557_Y), .A(T15673_Y));
KC_XNOR2_X1 T232 ( .B(T8824_Y), .A(T8878_Y), .Y(T232_Y));
KC_XNOR2_X1 T239 ( .B(T9026_Y), .A(T9134_Y), .Y(T239_Y));
KC_XNOR2_X1 T252 ( .B(T253_Y), .A(T8141_Y), .Y(T252_Y));
KC_XNOR2_X1 T554 ( .B(T11277_Y), .A(T1417_Y), .Y(T554_Y));
KC_XNOR2_X1 T612 ( .B(T15104_Y), .A(T15880_Q), .Y(T612_Y));
KC_XNOR2_X1 T613 ( .B(T15103_Y), .A(T15880_Q), .Y(T613_Y));
KC_XNOR2_X1 T777 ( .B(T9224_S), .A(T9467_Y), .Y(T777_Y));
KC_XNOR2_X1 T778 ( .B(T9239_S), .A(T9465_Y), .Y(T778_Y));
KC_XNOR2_X1 T854 ( .B(T383_Y), .A(T279_Y), .Y(T854_Y));
KC_XNOR2_X1 T1279 ( .B(T15161_Y), .A(T15860_Q), .Y(T1279_Y));
KC_XNOR2_X1 T1371 ( .B(T1738_Y), .A(T4819_Y), .Y(T1371_Y));
KC_XNOR2_X1 T1372 ( .B(T1371_Y), .A(T1357_Y), .Y(T1372_Y));
KC_XNOR2_X1 T1521 ( .B(T13494_Q), .A(T6894_Y), .Y(T1521_Y));
KC_XNOR2_X1 T2006 ( .B(T9941_Y), .A(T16465_Q), .Y(T2006_Y));
KC_XNOR2_X1 T2021 ( .B(T2003_Y), .A(T13029_Q), .Y(T2021_Y));
KC_XNOR2_X1 T2122 ( .B(T8199_Y), .A(T11458_Y), .Y(T2122_Y));
KC_XNOR2_X1 T2164 ( .B(T11463_Y), .A(T15915_Y), .Y(T2164_Y));
KC_XNOR2_X1 T2189 ( .B(T2172_Y), .A(T2184_Y), .Y(T2189_Y));
KC_XNOR2_X1 T2354 ( .B(T8418_Y), .A(T6569_Y), .Y(T2354_Y));
KC_XNOR2_X1 T2376 ( .B(T6491_Y), .A(T2933_Y), .Y(T2376_Y));
KC_XNOR2_X1 T2389 ( .B(T6540_Y), .A(T4962_Y), .Y(T2389_Y));
KC_XNOR2_X1 T2399 ( .B(T11033_Y), .A(T5546_Y), .Y(T2399_Y));
KC_XNOR2_X1 T2541 ( .B(T2538_Q), .A(T8358_Y), .Y(T2541_Y));
KC_XNOR2_X1 T2576 ( .B(T2547_Y), .A(T5869_S), .Y(T2576_Y));
KC_XNOR2_X1 T2741 ( .B(T8208_Y), .A(T11472_Y), .Y(T2741_Y));
KC_XNOR2_X1 T2747 ( .B(T5449_Q), .A(T10640_Y), .Y(T2747_Y));
KC_XNOR2_X1 T2760 ( .B(T11498_Y), .A(T2764_Y), .Y(T2760_Y));
KC_XNOR2_X1 T2764 ( .B(T8269_Y), .A(T3352_Y), .Y(T2764_Y));
KC_XNOR2_X1 T2766 ( .B(T11516_Y), .A(T15991_Y), .Y(T2766_Y));
KC_XNOR2_X1 T2767 ( .B(T11489_Y), .A(T2759_Q), .Y(T2767_Y));
KC_XNOR2_X1 T2785 ( .B(T11567_Y), .A(T15444_Y), .Y(T2785_Y));
KC_XNOR2_X1 T2786 ( .B(T2122_Y), .A(T2789_Y), .Y(T2786_Y));
KC_XNOR2_X1 T2787 ( .B(T11565_Y), .A(T11593_Y), .Y(T2787_Y));
KC_XNOR2_X1 T2808 ( .B(T11580_Y), .A(T8334_Y), .Y(T2808_Y));
KC_XNOR2_X1 T2941 ( .B(T2945_Q), .A(T8435_Y), .Y(T2941_Y));
KC_XNOR2_X1 T2948 ( .B(T4159_Y), .A(T2942_Q), .Y(T2948_Y));
KC_XNOR2_X1 T2959 ( .B(T12878_Y), .A(T2954_Q), .Y(T2959_Y));
KC_XNOR2_X1 T3219 ( .B(T6726_Y), .A(T3205_Y), .Y(T3219_Y));
KC_XNOR2_X1 T3268 ( .B(T11456_Y), .A(T3270_Y), .Y(T3268_Y));
KC_XNOR2_X1 T3274 ( .B(T3263_Y), .A(T3255_Y), .Y(T3274_Y));
KC_XNOR2_X1 T3305 ( .B(T11457_Y), .A(T6206_Y), .Y(T3305_Y));
KC_XNOR2_X1 T3310 ( .B(T15944_Y), .A(T11497_Y), .Y(T3310_Y));
KC_XNOR2_X1 T3329 ( .B(T12027_Y), .A(T3318_Y), .Y(T3329_Y));
KC_XNOR2_X1 T3330 ( .B(T11558_Y), .A(T13126_Q), .Y(T3330_Y));
KC_XNOR2_X1 T3334 ( .B(T11559_Y), .A(T11592_Y), .Y(T3334_Y));
KC_XNOR2_X1 T3335 ( .B(T15127_Y), .A(T11579_Y), .Y(T3335_Y));
KC_XNOR2_X1 T3360 ( .B(T16015_Y), .A(T3351_Y), .Y(T3360_Y));
KC_XNOR2_X1 T3680 ( .B(T16230_Y), .A(T3658_Y), .Y(T3680_Y));
KC_XNOR2_X1 T3822 ( .B(T10282_Y), .A(T3814_Y), .Y(T3822_Y));
KC_XNOR2_X1 T3897 ( .B(T2077_Y), .A(T5905_Y), .Y(T3897_Y));
KC_XNOR2_X1 T3951 ( .B(T4565_Y), .A(T11525_Y), .Y(T3951_Y));
KC_XNOR2_X1 T3963 ( .B(T4411_Y), .A(T15981_Y), .Y(T3963_Y));
KC_XNOR2_X1 T3992 ( .B(T8330_Y), .A(T11545_Y), .Y(T3992_Y));
KC_XNOR2_X1 T4042 ( .B(T16029_Y), .A(T6033_Y), .Y(T4042_Y));
KC_XNOR2_X1 T4046 ( .B(T4053_Y), .A(T4044_Q), .Y(T4046_Y));
KC_XNOR2_X1 T4148 ( .B(T3528_Q), .A(T5072_Y), .Y(T4148_Y));
KC_XNOR2_X1 T4167 ( .B(T4173_Y), .A(T4161_Y), .Y(T4167_Y));
KC_XNOR2_X1 T4275 ( .B(T4284_Y), .A(T4277_Y), .Y(T4275_Y));
KC_XNOR2_X1 T4317 ( .B(T14158_Q), .A(T4275_Y), .Y(T4317_Y));
KC_XNOR2_X1 T4457 ( .B(T5044_Y), .A(T4456_Q), .Y(T4457_Y));
KC_XNOR2_X1 T4463 ( .B(T4454_Q), .A(T15121_Y), .Y(T4463_Y));
KC_XNOR2_X1 T4489 ( .B(T15126_Y), .A(T4490_Q), .Y(T4489_Y));
KC_XNOR2_X1 T4497 ( .B(T4476_Y), .A(T4498_Q), .Y(T4497_Y));
KC_XNOR2_X1 T4500 ( .B(T5164_Q), .A(T16147_Y), .Y(T4500_Y));
KC_XNOR2_X1 T4530 ( .B(T4537_Q), .A(T3961_Y), .Y(T4530_Y));
KC_XNOR2_X1 T4535 ( .B(T4538_Q), .A(T15954_Y), .Y(T4535_Y));
KC_XNOR2_X1 T4541 ( .B(T3939_Y), .A(T4542_Y), .Y(T4541_Y));
KC_XNOR2_X1 T4565 ( .B(T6779_Y), .A(T4566_Y), .Y(T4565_Y));
KC_XNOR2_X1 T4617 ( .B(T16020_Y), .A(T16021_Y), .Y(T4617_Y));
KC_XNOR2_X1 T4622 ( .B(T8300_Y), .A(T16459_Q), .Y(T4622_Y));
KC_XNOR2_X1 T4623 ( .B(T16045_Y), .A(T4638_Y), .Y(T4623_Y));
KC_XNOR2_X1 T4665 ( .B(T8366_Y), .A(T4690_Y), .Y(T4665_Y));
KC_XNOR2_X1 T4690 ( .B(T4661_Y), .A(T6029_Y), .Y(T4690_Y));
KC_XNOR2_X1 T4711 ( .B(T4713_Q), .A(T4719_Q), .Y(T4711_Y));
KC_XNOR2_X1 T4712 ( .B(T4709_Y), .A(T4699_Y), .Y(T4712_Y));
KC_XNOR2_X1 T4807 ( .B(T9452_Y), .A(T9494_Y), .Y(T4807_Y));
KC_XNOR2_X1 T4808 ( .B(T1449_Y), .A(T9451_Y), .Y(T4808_Y));
KC_XNOR2_X1 T9482 ( .B(T9485_Y), .A(T9495_Y), .Y(T9482_Y));
KC_XNOR2_X1 T4921 ( .B(T5289_Y), .A(T1694_Q), .Y(T4921_Y));
KC_XNOR2_X1 T4974 ( .B(T15052_Y), .A(T15153_Y), .Y(T4974_Y));
KC_XNOR2_X1 T5011 ( .B(T2761_Y), .A(T2779_Y), .Y(T5011_Y));
KC_XNOR2_X1 T5012 ( .B(T15998_Y), .A(T11566_Y), .Y(T5012_Y));
KC_XNOR2_X1 T5067 ( .B(T11578_Y), .A(T8323_Y), .Y(T5067_Y));
KC_XNOR2_X1 T5135 ( .B(T5543_Q), .A(T8165_Y), .Y(T5135_Y));
KC_XNOR2_X1 T5319 ( .B(T5320_Q), .A(T12649_Y), .Y(T5319_Y));
KC_XNOR2_X1 T5349 ( .B(T15056_Y), .A(T5355_Q), .Y(T5349_Y));
KC_XNOR2_X1 T5478 ( .B(T11578_Y), .A(T3347_Y), .Y(T5478_Y));
KC_XNOR2_X1 T5510 ( .B(T8348_Y), .A(T5511_Q), .Y(T5510_Y));
KC_XNOR2_X1 T5540 ( .B(T5538_Q), .A(T8423_Y), .Y(T5540_Y));
KC_XNOR2_X1 T9462 ( .B(T9188_S), .A(T9468_Y), .Y(T9462_Y));
KC_XNOR2_X1 T5569 ( .B(T10630_Y), .A(T10639_Y), .Y(T5569_Y));
KC_NOR2B_X1 T46 ( .B(T5606_Y), .AN(T5640_S), .Y(T46_Y));
KC_NOR2B_X1 T47 ( .B(T5606_Y), .AN(T5641_S), .Y(T47_Y));
KC_NOR2B_X1 T50 ( .B(T5606_Y), .AN(T5644_S), .Y(T50_Y));
KC_NOR2B_X1 T5591 ( .B(T5606_Y), .AN(T5643_S), .Y(T5591_Y));
KC_NOR2B_X1 T5585 ( .B(T5606_Y), .AN(T2397_Y), .Y(T5585_Y));
KC_NOR2B_X1 T51 ( .B(T5606_Y), .AN(T5639_S), .Y(T51_Y));
KC_NOR2B_X1 T5590 ( .B(T5606_Y), .AN(T5642_S), .Y(T5590_Y));
KC_NOR2B_X1 T57 ( .B(T5606_Y), .AN(T6850_S), .Y(T57_Y));
KC_NOR2B_X1 T61 ( .B(T5606_Y), .AN(T59_S), .Y(T61_Y));
KC_NOR2B_X1 T62 ( .B(T5606_Y), .AN(T5625_S), .Y(T62_Y));
KC_NOR2B_X1 T71 ( .B(T5606_Y), .AN(T5609_S), .Y(T71_Y));
KC_NOR2B_X1 T80 ( .B(T85_Q), .AN(T5187_Q), .Y(T80_Y));
KC_NOR2B_X1 T112 ( .B(T5618_Y), .AN(T8536_Y), .Y(T112_Y));
KC_NOR2B_X1 T120 ( .B(T5598_Y), .AN(T116_Y), .Y(T120_Y));
KC_NOR2B_X1 T127 ( .B(T14972_Y), .AN(T5613_Y), .Y(T127_Y));
KC_NOR2B_X1 T227 ( .B(T16006_Y), .AN(T234_Q), .Y(T227_Y));
KC_NOR2B_X1 T238 ( .B(T16006_Y), .AN(T238_AN), .Y(T238_Y));
KC_NOR2B_X1 T256 ( .B(T16006_Y), .AN(T15178_Q), .Y(T256_Y));
KC_NOR2B_X1 T279 ( .B(T15377_Y), .AN(T11048_Y), .Y(T279_Y));
KC_NOR2B_X1 T338 ( .B(T9350_Q), .AN(T5303_Q), .Y(T338_Y));
KC_NOR2B_X1 T508 ( .B(T521_Q), .AN(T522_Q), .Y(T508_Y));
KC_NOR2B_X1 T509 ( .B(T5283_Q), .AN(T9339_Q), .Y(T509_Y));
KC_NOR2B_X1 T723 ( .B(T15842_Y), .AN(T9446_Y), .Y(T723_Y));
KC_NOR2B_X1 T756 ( .B(T908_Y), .AN(T752_Q), .Y(T756_Y));
KC_NOR2B_X1 T775 ( .B(T11268_Y), .AN(T15658_Y), .Y(T775_Y));
KC_NOR2B_X1 T779 ( .B(T11268_Y), .AN(T9239_S), .Y(T779_Y));
KC_NOR2B_X1 T782 ( .B(T11268_Y), .AN(T16508_Y), .Y(T782_Y));
KC_NOR2B_X1 T787 ( .B(T11268_Y), .AN(T9225_S), .Y(T787_Y));
KC_NOR2B_X1 T788 ( .B(T11268_Y), .AN(T9224_S), .Y(T788_Y));
KC_NOR2B_X1 T934 ( .B(T15792_Y), .AN(T5309_Q), .Y(T934_Y));
KC_NOR2B_X1 T956 ( .B(T5376_Q), .AN(T8938_Y), .Y(T956_Y));
KC_NOR2B_X1 T965 ( .B(T961_Y), .AN(T758_Y), .Y(T965_Y));
KC_NOR2B_X1 T988 ( .B(T16006_Y), .AN(T3358_Y), .Y(T988_Y));
KC_NOR2B_X1 T1098 ( .B(T16423_Y), .AN(T12095_Y), .Y(T1098_Y));
KC_NOR2B_X1 T1111 ( .B(T5030_Y), .AN(T12095_Y), .Y(T1111_Y));
KC_NOR2B_X1 T1134 ( .B(T16149_Y), .AN(T10000_Y), .Y(T1134_Y));
KC_NOR2B_X1 T1258 ( .B(T10143_Y), .AN(T1365_Y), .Y(T1258_Y));
KC_NOR2B_X1 T1259 ( .B(T10143_Y), .AN(T4868_Y), .Y(T1259_Y));
KC_NOR2B_X1 T1260 ( .B(T10143_Y), .AN(T1362_Y), .Y(T1260_Y));
KC_NOR2B_X1 T1261 ( .B(T10143_Y), .AN(T1366_Y), .Y(T1261_Y));
KC_NOR2B_X1 T1263 ( .B(T10143_Y), .AN(T4902_Y), .Y(T1263_Y));
KC_NOR2B_X1 T1289 ( .B(T15544_Y), .AN(T1361_Q), .Y(T1289_Y));
KC_NOR2B_X1 T1326 ( .B(T6767_Y), .AN(T13609_Q), .Y(T1326_Y));
KC_NOR2B_X1 T1331 ( .B(T6767_Y), .AN(T13575_Q), .Y(T1331_Y));
KC_NOR2B_X1 T1332 ( .B(T6767_Y), .AN(T13597_Q), .Y(T1332_Y));
KC_NOR2B_X1 T1333 ( .B(T6767_Y), .AN(T13586_Q), .Y(T1333_Y));
KC_NOR2B_X1 T1351 ( .B(T4901_Y), .AN(T13946_Q), .Y(T1351_Y));
KC_NOR2B_X1 T1355 ( .B(T4901_Y), .AN(T14615_Q), .Y(T1355_Y));
KC_NOR2B_X1 T1375 ( .B(T13198_Q), .AN(T16081_Q), .Y(T1375_Y));
KC_NOR2B_X1 T1411 ( .B(T6767_Y), .AN(T13583_Q), .Y(T1411_Y));
KC_NOR2B_X1 T1412 ( .B(T6767_Y), .AN(T13585_Q), .Y(T1412_Y));
KC_NOR2B_X1 T1413 ( .B(T6767_Y), .AN(T13606_Q), .Y(T1413_Y));
KC_NOR2B_X1 T1414 ( .B(T6767_Y), .AN(T13573_Q), .Y(T1414_Y));
KC_NOR2B_X1 T1424 ( .B(T6767_Y), .AN(T13584_Q), .Y(T1424_Y));
KC_NOR2B_X1 T1432 ( .B(T6767_Y), .AN(T14726_Q), .Y(T1432_Y));
KC_NOR2B_X1 T1433 ( .B(T6767_Y), .AN(T14720_Q), .Y(T1433_Y));
KC_NOR2B_X1 T1434 ( .B(T6767_Y), .AN(T14728_Q), .Y(T1434_Y));
KC_NOR2B_X1 T1435 ( .B(T6767_Y), .AN(T13603_Q), .Y(T1435_Y));
KC_NOR2B_X1 T1436 ( .B(T6767_Y), .AN(T14725_Q), .Y(T1436_Y));
KC_NOR2B_X1 T1437 ( .B(T6767_Y), .AN(T14727_Q), .Y(T1437_Y));
KC_NOR2B_X1 T1441 ( .B(T6767_Y), .AN(T13692_Q), .Y(T1441_Y));
KC_NOR2B_X1 T1443 ( .B(T6767_Y), .AN(T13691_Q), .Y(T1443_Y));
KC_NOR2B_X1 T1444 ( .B(T6767_Y), .AN(T13717_Q), .Y(T1444_Y));
KC_NOR2B_X1 T1447 ( .B(T6767_Y), .AN(T14662_Q), .Y(T1447_Y));
KC_NOR2B_X1 T1461 ( .B(T4901_Y), .AN(T13812_Q), .Y(T1461_Y));
KC_NOR2B_X1 T1470 ( .B(T4901_Y), .AN(T13959_Q), .Y(T1470_Y));
KC_NOR2B_X1 T1473 ( .B(T4901_Y), .AN(T14013_Q), .Y(T1473_Y));
KC_NOR2B_X1 T1474 ( .B(T4901_Y), .AN(T13978_Q), .Y(T1474_Y));
KC_NOR2B_X1 T1475 ( .B(T4901_Y), .AN(T13958_Q), .Y(T1475_Y));
KC_NOR2B_X1 T1478 ( .B(T4901_Y), .AN(T14616_Q), .Y(T1478_Y));
KC_NOR2B_X1 T1486 ( .B(T4901_Y), .AN(T14127_Q), .Y(T1486_Y));
KC_NOR2B_X1 T1488 ( .B(T4901_Y), .AN(T14129_Q), .Y(T1488_Y));
KC_NOR2B_X1 T1489 ( .B(T4901_Y), .AN(T14126_Q), .Y(T1489_Y));
KC_NOR2B_X1 T1490 ( .B(T4901_Y), .AN(T14128_Q), .Y(T1490_Y));
KC_NOR2B_X1 T1494 ( .B(T4901_Y), .AN(T14614_Q), .Y(T1494_Y));
KC_NOR2B_X1 T1580 ( .B(T4901_Y), .AN(T14608_Q), .Y(T1580_Y));
KC_NOR2B_X1 T1581 ( .B(T16395_Y), .AN(T14125_Q), .Y(T1581_Y));
KC_NOR2B_X1 T1582 ( .B(T16395_Y), .AN(T14609_Q), .Y(T1582_Y));
KC_NOR2B_X1 T1583 ( .B(T16395_Y), .AN(T14611_Q), .Y(T1583_Y));
KC_NOR2B_X1 T1637 ( .B(T6765_Y), .AN(T5661_Y), .Y(T1637_Y));
KC_NOR2B_X1 T1727 ( .B(T16306_Q), .AN(T1723_Q), .Y(T1727_Y));
KC_NOR2B_X1 T1752 ( .B(T15904_Y), .AN(T1803_Q), .Y(T1752_Y));
KC_NOR2B_X1 T2018 ( .B(T1117_Y), .AN(T1996_Y), .Y(T2018_Y));
KC_NOR2B_X1 T2026 ( .B(T1102_Y), .AN(T13028_Q), .Y(T2026_Y));
KC_NOR2B_X1 T2121 ( .B(T5820_Y), .AN(T6097_S), .Y(T2121_Y));
KC_NOR2B_X1 T2163 ( .B(T11970_Y), .AN(T4943_Y), .Y(T2163_Y));
KC_NOR2B_X1 T2248 ( .B(T13132_Q), .AN(T2152_Q), .Y(T2248_Y));
KC_NOR2B_X1 T2352 ( .B(T6566_Y), .AN(T2317_Y), .Y(T2352_Y));
KC_NOR2B_X1 T2356 ( .B(T2329_Y), .AN(T2324_Y), .Y(T2356_Y));
KC_NOR2B_X1 T2386 ( .B(T7836_Y), .AN(T6502_Y), .Y(T2386_Y));
KC_NOR2B_X1 T2395 ( .B(T8436_Y), .AN(T6495_Y), .Y(T2395_Y));
KC_NOR2B_X1 T2434 ( .B(T15682_Y), .AN(T13639_Q), .Y(T2434_Y));
KC_NOR2B_X1 T2435 ( .B(T15682_Y), .AN(T14765_Q), .Y(T2435_Y));
KC_NOR2B_X1 T2436 ( .B(T15682_Y), .AN(T13656_Q), .Y(T2436_Y));
KC_NOR2B_X1 T2440 ( .B(T15682_Y), .AN(T13657_Q), .Y(T2440_Y));
KC_NOR2B_X1 T2453 ( .B(T15682_Y), .AN(T13782_Q), .Y(T2453_Y));
KC_NOR2B_X1 T2489 ( .B(T15422_Y), .AN(T14836_Q), .Y(T2489_Y));
KC_NOR2B_X1 T2493 ( .B(T15422_Y), .AN(T14856_Q), .Y(T2493_Y));
KC_NOR2B_X1 T2533 ( .B(T5026_Y), .AN(T14857_Q), .Y(T2533_Y));
KC_NOR2B_X1 T2536 ( .B(T5026_Y), .AN(T14083_Q), .Y(T2536_Y));
KC_NOR2B_X1 T2537 ( .B(T5026_Y), .AN(T14069_Q), .Y(T2537_Y));
KC_NOR2B_X1 T2585 ( .B(T2013_Y), .AN(T5869_Co), .Y(T2585_Y));
KC_NOR2B_X1 T2586 ( .B(T2573_Y), .AN(T2547_Y), .Y(T2586_Y));
KC_NOR2B_X1 T2587 ( .B(T2013_Y), .AN(T5869_Co), .Y(T2587_Y));
KC_NOR2B_X1 T2619 ( .B(T15533_Y), .AN(T14366_Q), .Y(T2619_Y));
KC_NOR2B_X1 T2623 ( .B(T2597_Y), .AN(T2844_Q), .Y(T2623_Y));
KC_NOR2B_X1 T2644 ( .B(T15533_Y), .AN(T14425_Q), .Y(T2644_Y));
KC_NOR2B_X1 T2645 ( .B(T15533_Y), .AN(T14427_Q), .Y(T2645_Y));
KC_NOR2B_X1 T2646 ( .B(T15533_Y), .AN(T14403_Q), .Y(T2646_Y));
KC_NOR2B_X1 T2647 ( .B(T15533_Y), .AN(T14426_Q), .Y(T2647_Y));
KC_NOR2B_X1 T2649 ( .B(T15533_Y), .AN(T14345_Q), .Y(T2649_Y));
KC_NOR2B_X1 T2650 ( .B(T15533_Y), .AN(T14363_Q), .Y(T2650_Y));
KC_NOR2B_X1 T2670 ( .B(T2643_Y), .AN(T2512_Y), .Y(T2670_Y));
KC_NOR2B_X1 T2671 ( .B(T2643_Y), .AN(T2509_Y), .Y(T2671_Y));
KC_NOR2B_X1 T2672 ( .B(T11355_Y), .AN(T10252_Y), .Y(T2672_Y));
KC_NOR2B_X1 T2673 ( .B(T2643_Y), .AN(T2513_Y), .Y(T2673_Y));
KC_NOR2B_X1 T2693 ( .B(T2676_Y), .AN(T2656_Y), .Y(T2693_Y));
KC_NOR2B_X1 T2695 ( .B(T11960_Y), .AN(T2686_Y), .Y(T2695_Y));
KC_NOR2B_X1 T2707 ( .B(T15943_Y), .AN(T16033_Y), .Y(T2707_Y));
KC_NOR2B_X1 T2718 ( .B(T2107_Y), .AN(T2106_Y), .Y(T2718_Y));
KC_NOR2B_X1 T2739 ( .B(T13112_Q), .AN(T2735_Q), .Y(T2739_Y));
KC_NOR2B_X1 T2740 ( .B(T13111_Q), .AN(T2746_Q), .Y(T2740_Y));
KC_NOR2B_X1 T2763 ( .B(T11463_Y), .AN(T6186_Y), .Y(T2763_Y));
KC_NOR2B_X1 T2838 ( .B(T8394_Y), .AN(T16305_Y), .Y(T2838_Y));
KC_NOR2B_X1 T2846 ( .B(T5014_Y), .AN(T5999_Y), .Y(T2846_Y));
KC_NOR2B_X1 T2869 ( .B(T11724_Y), .AN(T3214_Y), .Y(T2869_Y));
KC_NOR2B_X1 T2870 ( .B(T2871_Y), .AN(T3425_Y), .Y(T2870_Y));
KC_NOR2B_X1 T2927 ( .B(T6225_Y), .AN(T11770_Y), .Y(T2927_Y));
KC_NOR2B_X1 T2929 ( .B(T2926_Y), .AN(T2890_Y), .Y(T2929_Y));
KC_NOR2B_X1 T2946 ( .B(T11846_Y), .AN(T2932_Y), .Y(T2946_Y));
KC_NOR2B_X1 T3021 ( .B(T15422_Y), .AN(T13755_Q), .Y(T3021_Y));
KC_NOR2B_X1 T3022 ( .B(T15422_Y), .AN(T14930_Q), .Y(T3022_Y));
KC_NOR2B_X1 T3023 ( .B(T15422_Y), .AN(T14761_Q), .Y(T3023_Y));
KC_NOR2B_X1 T3074 ( .B(T5026_Y), .AN(T14882_Q), .Y(T3074_Y));
KC_NOR2B_X1 T3077 ( .B(T5026_Y), .AN(T14081_Q), .Y(T3077_Y));
KC_NOR2B_X1 T3078 ( .B(T422_Y), .AN(T2648_Y), .Y(T3078_Y));
KC_NOR2B_X1 T3116 ( .B(T5026_Y), .AN(T14152_Q), .Y(T3116_Y));
KC_NOR2B_X1 T3118 ( .B(T5026_Y), .AN(T14172_Q), .Y(T3118_Y));
KC_NOR2B_X1 T3119 ( .B(T5026_Y), .AN(T14892_Q), .Y(T3119_Y));
KC_NOR2B_X1 T3120 ( .B(T5026_Y), .AN(T14151_Q), .Y(T3120_Y));
KC_NOR2B_X1 T3121 ( .B(T5026_Y), .AN(T14198_Q), .Y(T3121_Y));
KC_NOR2B_X1 T3123 ( .B(T5026_Y), .AN(T15072_Q), .Y(T3123_Y));
KC_NOR2B_X1 T3147 ( .B(T5026_Y), .AN(T14893_Q), .Y(T3147_Y));
KC_NOR2B_X1 T3148 ( .B(T5026_Y), .AN(T14404_Q), .Y(T3148_Y));
KC_NOR2B_X1 T3157 ( .B(T5026_Y), .AN(T14303_Q), .Y(T3157_Y));
KC_NOR2B_X1 T3241 ( .B(T5575_Q), .AN(T10256_Y), .Y(T3241_Y));
KC_NOR2B_X1 T3267 ( .B(T3269_Y), .AN(T3252_Y), .Y(T3267_Y));
KC_NOR2B_X1 T3272 ( .B(T5022_Y), .AN(T13316_Q), .Y(T3272_Y));
KC_NOR2B_X1 T3273 ( .B(T5022_Y), .AN(T13103_Q), .Y(T3273_Y));
KC_NOR2B_X1 T3276 ( .B(T5022_Y), .AN(T13297_Q), .Y(T3276_Y));
KC_NOR2B_X1 T3343 ( .B(T12215_Y), .AN(T8275_Y), .Y(T3343_Y));
KC_NOR2B_X1 T3362 ( .B(T4052_Q), .AN(T9056_Y), .Y(T3362_Y));
KC_NOR2B_X1 T3364 ( .B(T6555_Q), .AN(T12263_Y), .Y(T3364_Y));
KC_NOR2B_X1 T3404 ( .B(T5052_Y), .AN(T12042_Y), .Y(T3404_Y));
KC_NOR2B_X1 T3409 ( .B(T11643_Y), .AN(T11645_Y), .Y(T3409_Y));
KC_NOR2B_X1 T3413 ( .B(T4035_Y), .AN(T11630_Y), .Y(T3413_Y));
KC_NOR2B_X1 T3454 ( .B(T6158_Y), .AN(T11644_Y), .Y(T3454_Y));
KC_NOR2B_X1 T3527 ( .B(T11006_Y), .AN(T3522_Q), .Y(T3527_Y));
KC_NOR2B_X1 T3530 ( .B(T11007_Y), .AN(T11833_Y), .Y(T3530_Y));
KC_NOR2B_X1 T3823 ( .B(T13308_Y), .AN(T3815_Y), .Y(T3823_Y));
KC_NOR2B_X1 T3854 ( .B(T3242_Q), .AN(T3241_Y), .Y(T3854_Y));
KC_NOR2B_X1 T3874 ( .B(T5454_Y), .AN(T16501_Y), .Y(T3874_Y));
KC_NOR2B_X1 T3875 ( .B(T5454_Y), .AN(T6146_S), .Y(T3875_Y));
KC_NOR2B_X1 T3881 ( .B(T5454_Y), .AN(T6131_S), .Y(T3881_Y));
KC_NOR2B_X1 T3886 ( .B(T6797_S), .AN(T15939_Y), .Y(T3886_Y));
KC_NOR2B_X1 T3887 ( .B(T3871_Y), .AN(T12184_Y), .Y(T3887_Y));
KC_NOR2B_X1 T3891 ( .B(T5454_Y), .AN(T6142_S), .Y(T3891_Y));
KC_NOR2B_X1 T3892 ( .B(T5454_Y), .AN(T6132_S), .Y(T3892_Y));
KC_NOR2B_X1 T3893 ( .B(T5454_Y), .AN(T6130_S), .Y(T3893_Y));
KC_NOR2B_X1 T3894 ( .B(T5454_Y), .AN(T6143_S), .Y(T3894_Y));
KC_NOR2B_X1 T3896 ( .B(T12804_Y), .AN(T15919_Y), .Y(T3896_Y));
KC_NOR2B_X1 T3925 ( .B(T8264_Y), .AN(T3904_Y), .Y(T3925_Y));
KC_NOR2B_X1 T3952 ( .B(T5022_Y), .AN(T13312_Q), .Y(T3952_Y));
KC_NOR2B_X1 T3961 ( .B(T15985_Y), .AN(T3962_Y), .Y(T3961_Y));
KC_NOR2B_X1 T3962 ( .B(T6277_Y), .AN(T3972_Y), .Y(T3962_Y));
KC_NOR2B_X1 T3969 ( .B(T5022_Y), .AN(T3971_Q), .Y(T3969_Y));
KC_NOR2B_X1 T3988 ( .B(T4596_Y), .AN(T11607_Y), .Y(T3988_Y));
KC_NOR2B_X1 T3989 ( .B(T5022_Y), .AN(T13155_Q), .Y(T3989_Y));
KC_NOR2B_X1 T3997 ( .B(T5022_Y), .AN(T16416_Y), .Y(T3997_Y));
KC_NOR2B_X1 T4053 ( .B(T16028_Y), .AN(T12346_Y), .Y(T4053_Y));
KC_NOR2B_X1 T4095 ( .B(T12851_Y), .AN(T4061_Y), .Y(T4095_Y));
KC_NOR2B_X1 T4102 ( .B(T4084_Y), .AN(T10586_Y), .Y(T4102_Y));
KC_NOR2B_X1 T4106 ( .B(T15760_Q), .AN(T4023_Y), .Y(T4106_Y));
KC_NOR2B_X1 T4165 ( .B(T9163_Y), .AN(T4173_Y), .Y(T4165_Y));
KC_NOR2B_X1 T4166 ( .B(T4156_Y), .AN(T4151_Y), .Y(T4166_Y));
KC_NOR2B_X1 T4355 ( .B(T10257_Y), .AN(T5170_Q), .Y(T4355_Y));
KC_NOR2B_X1 T4356 ( .B(T10257_Y), .AN(T4361_Q), .Y(T4356_Y));
KC_NOR2B_X1 T4357 ( .B(T10257_Y), .AN(T4359_Q), .Y(T4357_Y));
KC_NOR2B_X1 T4358 ( .B(T10257_Y), .AN(T4362_Q), .Y(T4358_Y));
KC_NOR2B_X1 T4364 ( .B(T10257_Y), .AN(T4370_Q), .Y(T4364_Y));
KC_NOR2B_X1 T4365 ( .B(T10257_Y), .AN(T4375_Q), .Y(T4365_Y));
KC_NOR2B_X1 T4366 ( .B(T10257_Y), .AN(T4367_Q), .Y(T4366_Y));
KC_NOR2B_X1 T4371 ( .B(T10257_Y), .AN(T4369_Q), .Y(T4371_Y));
KC_NOR2B_X1 T4372 ( .B(T10257_Y), .AN(T4368_Q), .Y(T4372_Y));
KC_NOR2B_X1 T4373 ( .B(T10257_Y), .AN(T4376_Q), .Y(T4373_Y));
KC_NOR2B_X1 T4377 ( .B(T10257_Y), .AN(T4374_Q), .Y(T4377_Y));
KC_NOR2B_X1 T4378 ( .B(T10257_Y), .AN(T4380_Q), .Y(T4378_Y));
KC_NOR2B_X1 T4379 ( .B(T10257_Y), .AN(T4360_Q), .Y(T4379_Y));
KC_NOR2B_X1 T4418 ( .B(T15837_Y), .AN(T420_Y), .Y(T4418_Y));
KC_NOR2B_X1 T4459 ( .B(T4462_Y), .AN(T8195_Y), .Y(T4459_Y));
KC_NOR2B_X1 T4482 ( .B(T4497_Y), .AN(T11454_Y), .Y(T4482_Y));
KC_NOR2B_X1 T4488 ( .B(T4470_Y), .AN(T5142_Y), .Y(T4488_Y));
KC_NOR2B_X1 T4495 ( .B(T4488_Y), .AN(T11466_Y), .Y(T4495_Y));
KC_NOR2B_X1 T4496 ( .B(T5454_Y), .AN(T6168_S), .Y(T4496_Y));
KC_NOR2B_X1 T4523 ( .B(T10925_Y), .AN(T10629_Y), .Y(T4523_Y));
KC_NOR2B_X1 T4529 ( .B(T5154_Y), .AN(T4531_Y), .Y(T4529_Y));
KC_NOR2B_X1 T4534 ( .B(T10939_Y), .AN(T4482_Y), .Y(T4534_Y));
KC_NOR2B_X1 T4539 ( .B(T9487_Y), .AN(T15963_Y), .Y(T4539_Y));
KC_NOR2B_X1 T4574 ( .B(T2757_Y), .AN(T4555_Y), .Y(T4574_Y));
KC_NOR2B_X1 T4577 ( .B(T4556_Y), .AN(T11542_Y), .Y(T4577_Y));
KC_NOR2B_X1 T4600 ( .B(T4621_Y), .AN(T4613_Y), .Y(T4600_Y));
KC_NOR2B_X1 T4603 ( .B(T2757_Y), .AN(T12018_Y), .Y(T4603_Y));
KC_NOR2B_X1 T4715 ( .B(T12281_Y), .AN(T6151_Y), .Y(T4715_Y));
KC_NOR2B_X1 T4724 ( .B(T8390_Y), .AN(T4697_Y), .Y(T4724_Y));
KC_NOR2B_X1 T4747 ( .B(T11758_Y), .AN(T6420_Co), .Y(T4747_Y));
KC_NOR2B_X1 T15725 ( .B(T524_Q), .AN(T363_Q), .Y(T15725_Y));
KC_NOR2B_X1 T4880 ( .B(T4901_Y), .AN(T14613_Q), .Y(T4880_Y));
KC_NOR2B_X1 T4887 ( .B(T16395_Y), .AN(T14661_Q), .Y(T4887_Y));
KC_NOR2B_X1 T4890 ( .B(T4901_Y), .AN(T13941_Q), .Y(T4890_Y));
KC_NOR2B_X1 T4891 ( .B(T4901_Y), .AN(T13942_Q), .Y(T4891_Y));
KC_NOR2B_X1 T4899 ( .B(T4901_Y), .AN(T14612_Q), .Y(T4899_Y));
KC_NOR2B_X1 T4903 ( .B(T16395_Y), .AN(T14607_Q), .Y(T4903_Y));
KC_NOR2B_X1 T4904 ( .B(T16395_Y), .AN(T14610_Q), .Y(T4904_Y));
KC_NOR2B_X1 T4920 ( .B(T4919_Y), .AN(T10757_Y), .Y(T4920_Y));
KC_NOR2B_X1 T16268 ( .B(T5508_Y), .AN(T16040_Y), .Y(T16268_Y));
KC_NOR2B_X1 T4973 ( .B(T4983_Y), .AN(T1665_Q), .Y(T4973_Y));
KC_NOR2B_X1 T4980 ( .B(T2374_Y), .AN(T2393_Y), .Y(T4980_Y));
KC_NOR2B_X1 T5020 ( .B(T13073_Y), .AN(T2654_Y), .Y(T5020_Y));
KC_NOR2B_X1 T5024 ( .B(T2583_Q), .AN(T10517_Y), .Y(T5024_Y));
KC_NOR2B_X1 T5062 ( .B(T16503_Y), .AN(T5064_Y), .Y(T5062_Y));
KC_NOR2B_X1 T5079 ( .B(T5026_Y), .AN(T14881_Q), .Y(T5079_Y));
KC_NOR2B_X1 T5081 ( .B(T15422_Y), .AN(T13653_Q), .Y(T5081_Y));
KC_NOR2B_X1 T5116 ( .B(T3383_Y), .AN(T11764_Y), .Y(T5116_Y));
KC_NOR2B_X1 T5163 ( .B(T13081_Y), .AN(T3800_Y), .Y(T5163_Y));
KC_NOR2B_X1 T5166 ( .B(T10257_Y), .AN(T4406_Q), .Y(T5166_Y));
KC_NOR2B_X1 T5167 ( .B(T10257_Y), .AN(T4427_Q), .Y(T5167_Y));
KC_NOR2B_X1 T5168 ( .B(T16157_Y), .AN(T12950_Y), .Y(T5168_Y));
KC_NOR2B_X1 T5171 ( .B(T10257_Y), .AN(T4363_Q), .Y(T5171_Y));
KC_NOR2B_X1 T5172 ( .B(T10257_Y), .AN(T4351_Q), .Y(T5172_Y));
KC_NOR2B_X1 T5236 ( .B(T6767_Y), .AN(T13607_Q), .Y(T5236_Y));
KC_NOR2B_X1 T5256 ( .B(T7254_Y), .AN(T4810_Q), .Y(T5256_Y));
KC_NOR2B_X1 T5295 ( .B(T4901_Y), .AN(T13943_Q), .Y(T5295_Y));
KC_NOR2B_X1 T5302 ( .B(T16091_Y), .AN(T5301_Q), .Y(T5302_Y));
KC_NOR2B_X1 T5316 ( .B(T5026_Y), .AN(T13894_Q), .Y(T5316_Y));
KC_NOR2B_X1 T5317 ( .B(T5026_Y), .AN(T14051_Q), .Y(T5317_Y));
KC_NOR2B_X1 T5338 ( .B(T4901_Y), .AN(T14124_Q), .Y(T5338_Y));
KC_NOR2B_X1 T5358 ( .B(T903_Y), .AN(T1249_Q), .Y(T5358_Y));
KC_NOR2B_X1 T5409 ( .B(T2717_Y), .AN(T5731_Y), .Y(T5409_Y));
KC_NOR2B_X1 T5419 ( .B(T11268_Y), .AN(T9188_S), .Y(T5419_Y));
KC_NOR2B_X1 T5453 ( .B(T5454_Y), .AN(T6167_S), .Y(T5453_Y));
KC_NOR2B_X1 T5454 ( .B(T5457_Y), .AN(T11451_Y), .Y(T5454_Y));
KC_NOR2B_X1 T5546 ( .B(T2395_Y), .AN(T2394_Y), .Y(T5546_Y));
KC_NOR2B_X1 T5570 ( .B(T6549_Q), .AN(T3364_Y), .Y(T5570_Y));
KC_OR2_X2 T23 ( .Y(T23_Y), .A(T24_Y), .B(T13068_Y));
KC_OR2_X2 T25 ( .Y(T25_Y), .A(T30_Y), .B(T13068_Y));
KC_OR2_X2 T38 ( .Y(T38_Y), .A(T37_Y), .B(T13075_Y));
KC_OR2_X2 T64 ( .Y(T64_Y), .A(T63_Y), .B(T70_Y));
KC_OR2_X2 T76 ( .Y(T76_Y), .A(T74_Y), .B(T70_Y));
KC_OR2_X2 T113 ( .Y(T113_Y), .A(T111_Y), .B(T15321_Y));
KC_OR2_X2 T194 ( .Y(T194_Y), .A(T193_Y), .B(T15407_Y));
KC_OR2_X2 T195 ( .Y(T195_Y), .A(T7608_Y), .B(T14972_Y));
KC_OR2_X2 T463 ( .Y(T463_Y), .A(T462_Y), .B(T15369_Y));
KC_OR2_X2 T471 ( .Y(T471_Y), .A(T470_Y), .B(T15369_Y));
KC_OR2_X2 T574 ( .Y(T574_Y), .A(T580_Y), .B(T15484_Y));
KC_OR2_X2 T581 ( .Y(T581_Y), .A(T537_Y), .B(T15484_Y));
KC_OR2_X2 T805 ( .Y(T805_Y), .A(T795_Y), .B(T15335_Y));
KC_OR2_X2 T806 ( .Y(T806_Y), .A(T804_Y), .B(T15335_Y));
KC_OR2_X2 T873 ( .Y(T873_Y), .A(T897_Y), .B(T15411_Y));
KC_OR2_X2 T888 ( .Y(T888_Y), .A(T887_Y), .B(T15411_Y));
KC_OR2_X2 T1180 ( .Y(T1180_Y), .A(T1179_Y), .B(T15673_Y));
KC_OR2_X2 T1227 ( .Y(T1227_Y), .A(T1226_Y), .B(T15496_Y));
KC_OR2_X2 T1236 ( .Y(T1236_Y), .A(T1235_Y), .B(T15496_Y));
KC_OR2_X2 T1380 ( .Y(T1380_Y), .A(T15181_Q), .B(T15189_Q));
KC_OR2_X2 T1389 ( .Y(T1389_Y), .A(T1388_Y), .B(T15342_Y));
KC_OR2_X2 T1396 ( .Y(T1396_Y), .A(T1392_Y), .B(T15342_Y));
KC_OR2_X2 T1455 ( .Y(T1455_Y), .A(T1454_Y), .B(T15415_Y));
KC_OR2_X2 T1462 ( .Y(T1462_Y), .A(T1460_Y), .B(T15415_Y));
KC_OR2_X2 T1537 ( .Y(T1537_Y), .A(T1529_Y), .B(T8671_Y));
KC_OR2_X2 T1539 ( .Y(T1539_Y), .A(T1543_Y), .B(T8671_Y));
KC_OR2_X2 T1564 ( .Y(T1564_Y), .A(T1595_Y), .B(T984_Y));
KC_OR2_X2 T1596 ( .Y(T1596_Y), .A(T1577_Y), .B(T984_Y));
KC_OR2_X2 T1869 ( .Y(T1869_Y), .A(T1868_Y), .B(T15347_Y));
KC_OR2_X2 T1960 ( .Y(T1960_Y), .A(T1959_Y), .B(T6848_Y));
KC_OR2_X2 T2408 ( .Y(T2408_Y), .A(T2409_Y), .B(T15347_Y));
KC_OR2_X2 T2439 ( .Y(T2439_Y), .A(T5246_Y), .B(T15381_Y));
KC_OR2_X2 T2498 ( .Y(T2498_Y), .A(T2497_Y), .B(T6848_Y));
KC_OR2_X2 T3010 ( .Y(T3010_Y), .A(T3009_Y), .B(T15381_Y));
KC_OR2_X2 T3150 ( .Y(T3150_Y), .A(T3156_Y), .B(T16303_Y));
KC_OR2_X2 T3151 ( .Y(T3151_Y), .A(T3149_Y), .B(T16303_Y));
KC_OR2_X2 T3187 ( .Y(T3187_Y), .A(T3197_Y), .B(T15551_Y));
KC_OR2_X2 T3231 ( .Y(T3231_Y), .A(T3229_Y), .B(T15565_Y));
KC_OR2_X2 T3238 ( .Y(T3238_Y), .A(T3243_Y), .B(T15565_Y));
KC_OR2_X2 T16026 ( .Y(T16026_Y), .A(T3366_Y), .B(T4352_Y));
KC_OR2_X2 T3503 ( .Y(T3503_Y), .A(T3532_Y), .B(T15639_Y));
KC_OR2_X2 T3531 ( .Y(T3531_Y), .A(T3529_Y), .B(T15639_Y));
KC_OR2_X2 T3647 ( .Y(T3647_Y), .A(T3646_Y), .B(T3290_Y));
KC_OR2_X2 T3956 ( .Y(T3956_Y), .A(T3955_Y), .B(T15594_Y));
KC_OR2_X2 T4188 ( .Y(T4188_Y), .A(T4193_Y), .B(T15366_Y));
KC_OR2_X2 T4195 ( .Y(T4195_Y), .A(T4194_Y), .B(T15366_Y));
KC_OR2_X2 T4207 ( .Y(T4207_Y), .A(T4206_Y), .B(T6455_Y));
KC_OR2_X2 T4225 ( .Y(T4225_Y), .A(T4224_Y), .B(T6455_Y));
KC_OR2_X2 T4328 ( .Y(T4328_Y), .A(T4327_Y), .B(T2724_Y));
KC_OR2_X2 T4329 ( .Y(T4329_Y), .A(T4336_Y), .B(T2724_Y));
KC_OR2_X2 T4866 ( .Y(T4866_Y), .A(T1181_Y), .B(T15673_Y));
KC_OR2_X2 T5078 ( .Y(T5078_Y), .A(T3190_Y), .B(T15551_Y));
KC_OR2_X2 T5118 ( .Y(T5118_Y), .A(T5117_Y), .B(T15594_Y));
KC_OR2_X2 T5132 ( .Y(T5132_Y), .A(T3642_Y), .B(T3290_Y));
KC_OR2_X2 T5188 ( .Y(T5188_Y), .A(T95_Y), .B(T15321_Y));
KC_OR2_X2 T5191 ( .Y(T5191_Y), .A(T49_Y), .B(T13075_Y));
KC_OR2_X2 T5572 ( .Y(T5572_Y), .A(T3407_Y), .B(T4352_Y));
KC_DFFRNHQ_X2 T44 ( .Q(T44_Q), .D(T46_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T45 ( .Q(T45_Q), .D(T50_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T48 ( .Q(T48_Q), .D(T47_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T5586 ( .Q(T5586_Q), .D(T5585_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T54 ( .Q(T54_Q), .D(T57_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T5589 ( .Q(T5589_Q), .D(T5590_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T81 ( .Q(T81_Q), .D(T12370_Y), .RN(T15024_Y),     .CK(T16477_Y));
KC_DFFRNHQ_X2 T83 ( .Q(T83_Q), .D(T9251_Y), .RN(T15024_Y),     .CK(T16477_Y));
KC_DFFRNHQ_X2 T84 ( .Q(T84_Q), .D(T15166_Y), .RN(T15024_Y),     .CK(T16477_Y));
KC_DFFRNHQ_X2 T85 ( .Q(T85_Q), .D(T61_Y), .RN(T15024_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T98 ( .Q(T98_Q), .D(T9252_Y), .RN(T15024_Y),     .CK(T16477_Y));
KC_DFFRNHQ_X2 T101 ( .Q(T101_Q), .D(T12377_Y), .RN(T15024_Y),     .CK(T16477_Y));
KC_DFFRNHQ_X2 T103 ( .Q(T103_Q), .D(T60_Y), .RN(T15024_Y),     .CK(T13330_Q));
KC_DFFRNHQ_X2 T105 ( .Q(T105_Q), .D(T8547_Y), .RN(T7074_Y),     .CK(T138_Y));
KC_DFFRNHQ_X2 T107 ( .Q(T107_Q), .D(T121_Y), .RN(T15024_Y),     .CK(T13330_Q));
KC_DFFRNHQ_X2 T114 ( .Q(T114_Q), .D(T122_Y), .RN(T15024_Y),     .CK(T13330_Q));
KC_DFFRNHQ_X2 T131 ( .Q(T131_Q), .D(T6910_Y), .RN(T7073_Y),     .CK(T130_Y));
KC_DFFRNHQ_X2 T132 ( .Q(T132_Q), .D(T100_Y), .RN(T7073_Y),     .CK(T138_Y));
KC_DFFRNHQ_X2 T133 ( .Q(T133_Q), .D(T9297_Y), .RN(T7073_Y),     .CK(T130_Y));
KC_DFFRNHQ_X2 T134 ( .Q(T134_Q), .D(T8552_Y), .RN(T7074_Y),     .CK(T13330_Q));
KC_DFFRNHQ_X2 T135 ( .Q(T135_Q), .D(T12376_Y), .RN(T7073_Y),     .CK(T138_Y));
KC_DFFRNHQ_X2 T136 ( .Q(T136_Q), .D(T9296_Y), .RN(T7073_Y),     .CK(T130_Y));
KC_DFFRNHQ_X2 T150 ( .Q(T150_Q), .D(T8567_Y), .RN(T7074_Y),     .CK(T130_Y));
KC_DFFRNHQ_X2 T151 ( .Q(T151_Q), .D(T186_Y), .RN(T14975_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T153 ( .Q(T153_Q), .D(T186_Y), .RN(T14975_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T154 ( .Q(T154_Q), .D(T186_Y), .RN(T14975_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T155 ( .Q(T155_Q), .D(T176_Y), .RN(T869_Y), .CK(T178_Y));
KC_DFFRNHQ_X2 T157 ( .Q(T157_Q), .D(T186_Y), .RN(T14975_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T158 ( .Q(T158_Q), .D(T11082_Y), .RN(T14975_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T160 ( .Q(T160_Q), .D(T7108_Y), .RN(T14975_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T161 ( .Q(T161_Q), .D(T322_Y), .RN(T7074_Y),     .CK(T352_Y));
KC_DFFRNHQ_X2 T162 ( .Q(T162_Q), .D(T198_Y), .RN(T7074_Y),     .CK(T138_Y));
KC_DFFRNHQ_X2 T163 ( .Q(T163_Q), .D(T214_Y), .RN(T15721_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T164 ( .Q(T164_Q), .D(T214_Y), .RN(T15721_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T165 ( .Q(T165_Q), .D(T214_Y), .RN(T15721_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T166 ( .Q(T166_Q), .D(T16429_Y), .RN(T15721_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T167 ( .Q(T167_Q), .D(T11870_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T169 ( .Q(T169_Q), .D(T16376_Y), .RN(T14978_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T170 ( .Q(T170_Q), .D(T7812_Y), .RN(T14978_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T171 ( .Q(T171_Q), .D(T16376_Y), .RN(T14978_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T172 ( .Q(T172_Q), .D(T16376_Y), .RN(T14978_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T173 ( .Q(T173_Q), .D(T214_Y), .RN(T15721_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T174 ( .Q(T174_Q), .D(T11100_Y), .RN(T14978_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T177 ( .Q(T177_Q), .D(T16376_Y), .RN(T15721_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T179 ( .Q(T179_Q), .D(T176_Y), .RN(T14978_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T180 ( .Q(T180_Q), .D(T176_Y), .RN(T14978_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T181 ( .Q(T181_Q), .D(T10264_Y), .RN(T15721_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T182 ( .Q(T182_Q), .D(T11871_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T183 ( .Q(T183_Q), .D(T16429_Y), .RN(T15721_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T184 ( .Q(T184_Q), .D(T15425_Y), .RN(T15721_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T189 ( .Q(T189_Q), .D(T16429_Y), .RN(T15029_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T190 ( .Q(T190_Q), .D(T10264_Y), .RN(T15029_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T191 ( .Q(T191_Q), .D(T16429_Y), .RN(T15721_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T204 ( .Q(T204_Q), .D(T8808_Y), .RN(T15029_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T207 ( .Q(T207_Q), .D(T206_Y), .RN(T14976_Y),     .CK(T14589_Q));
KC_DFFRNHQ_X2 T208 ( .Q(T208_Q), .D(T8755_Y), .RN(T14976_Y),     .CK(T14589_Q));
KC_DFFRNHQ_X2 T211 ( .Q(T211_Q), .D(T210_Y), .RN(T14976_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X2 T212 ( .Q(T212_Q), .D(T648_Y), .RN(T14976_Y),     .CK(T14589_Q));
KC_DFFRNHQ_X2 T215 ( .Q(T215_Q), .D(T9356_Y), .RN(T14976_Y),     .CK(T4826_Y));
KC_DFFRNHQ_X2 T223 ( .Q(T223_Q), .D(T8744_Y), .RN(T14976_Y),     .CK(T14589_Q));
KC_DFFRNHQ_X2 T224 ( .Q(T224_Q), .D(T222_Y), .RN(T14976_Y),     .CK(T14589_Q));
KC_DFFRNHQ_X2 T234 ( .Q(T234_Q), .D(T238_Y), .RN(T7675_Y),     .CK(T4828_Y));
KC_DFFRNHQ_X2 T235 ( .Q(T235_Q), .D(T8786_Y), .RN(T14976_Y),     .CK(T4828_Y));
KC_DFFRNHQ_X2 T272 ( .Q(T272_Q), .D(T16162_Y), .RN(T14974_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T273 ( .Q(T273_Q), .D(T16162_Y), .RN(T14974_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T274 ( .Q(T274_Q), .D(T16162_Y), .RN(T14974_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T275 ( .Q(T275_Q), .D(T11062_Y), .RN(T14974_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T276 ( .Q(T276_Q), .D(T6809_Y), .RN(T14974_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T277 ( .Q(T277_Q), .D(T7606_Y), .RN(T14974_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T278 ( .Q(T278_Q), .D(T16162_Y), .RN(T14974_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T281 ( .Q(T281_Q), .D(T7108_Y), .RN(T14975_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T282 ( .Q(T282_Q), .D(T156_Y), .RN(T14975_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T283 ( .Q(T283_Q), .D(T7606_Y), .RN(T14974_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T284 ( .Q(T284_Q), .D(T7606_Y), .RN(T14976_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T288 ( .Q(T288_Q), .D(T11058_Y), .RN(T14976_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T289 ( .Q(T289_Q), .D(T7108_Y), .RN(T14975_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T293 ( .Q(T293_Q), .D(T12387_Y), .RN(T14974_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T294 ( .Q(T294_Q), .D(T7606_Y), .RN(T14974_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T296 ( .Q(T296_Q), .D(T11071_Y), .RN(T14974_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T306 ( .Q(T306_Q), .D(T11083_Y), .RN(T14978_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T313 ( .Q(T313_Q), .D(T11074_Y), .RN(T14975_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T316 ( .Q(T316_Q), .D(T7812_Y), .RN(T14978_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T319 ( .Q(T319_Q), .D(T11868_Y), .RN(T14978_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T320 ( .Q(T320_Q), .D(T11867_Y), .RN(T14979_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T323 ( .Q(T323_Q), .D(T11107_Y), .RN(T14978_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T326 ( .Q(T326_Q), .D(T11097_Y), .RN(T14978_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T329 ( .Q(T329_Q), .D(T11098_Y), .RN(T14978_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T330 ( .Q(T330_Q), .D(T7812_Y), .RN(T14978_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T9354 ( .Q(T9354_Q), .D(T15425_Y), .RN(T15029_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T9352 ( .Q(T9352_Q), .D(T11148_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T335 ( .Q(T335_Q), .D(T11159_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T337 ( .Q(T337_Q), .D(T11151_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T341 ( .Q(T341_Q), .D(T10264_Y), .RN(T15029_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T343 ( .Q(T343_Q), .D(T11161_Y), .RN(T15030_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T344 ( .Q(T344_Q), .D(T11160_Y), .RN(T15030_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T359 ( .Q(T359_Q), .D(T357_Y), .RN(T15030_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T360 ( .Q(T360_Q), .D(T357_Y), .RN(T15029_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T362 ( .Q(T362_Q), .D(T11168_Y), .RN(T15030_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T363 ( .Q(T363_Q), .D(T8808_Y), .RN(T15030_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T432 ( .Q(T432_Q), .D(T11051_Y), .RN(T15027_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T434 ( .Q(T434_Q), .D(T472_Y), .RN(T14974_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T435 ( .Q(T435_Q), .D(T6809_Y), .RN(T15027_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T436 ( .Q(T436_Q), .D(T11052_Y), .RN(T15027_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T438 ( .Q(T438_Q), .D(T7318_Y), .RN(T14974_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T439 ( .Q(T439_Q), .D(T472_Y), .RN(T14974_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T440 ( .Q(T440_Q), .D(T7318_Y), .RN(T14974_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T441 ( .Q(T441_Q), .D(T7318_Y), .RN(T15027_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T442 ( .Q(T442_Q), .D(T472_Y), .RN(T15027_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T443 ( .Q(T443_Q), .D(T6809_Y), .RN(T14974_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T445 ( .Q(T445_Q), .D(T11855_Y), .RN(T7242_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T446 ( .Q(T446_Q), .D(T455_Y), .RN(T7242_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T449 ( .Q(T449_Q), .D(T447_Y), .RN(T15027_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T450 ( .Q(T450_Q), .D(T11061_Y), .RN(T7242_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T452 ( .Q(T452_Q), .D(T11858_Y), .RN(T7242_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T453 ( .Q(T453_Q), .D(T11057_Y), .RN(T15027_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T456 ( .Q(T456_Q), .D(T11054_Y), .RN(T7242_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T459 ( .Q(T459_Q), .D(T11079_Y), .RN(T7242_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T460 ( .Q(T460_Q), .D(T11086_Y), .RN(T7242_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T489 ( .Q(T489_Q), .D(T11096_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T9338 ( .Q(T9338_Q), .D(T357_Y), .RN(T14985_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T500 ( .Q(T500_Q), .D(T11144_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T501 ( .Q(T501_Q), .D(T11145_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T512 ( .Q(T512_Q), .D(T11890_Y), .RN(T15030_Y),     .CK(T13936_Q));
KC_DFFRNHQ_X2 T517 ( .Q(T517_Q), .D(T11892_Y), .RN(T15030_Y),     .CK(T13936_Q));
KC_DFFRNHQ_X2 T519 ( .Q(T519_Q), .D(T11882_Y), .RN(T15030_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T521 ( .Q(T521_Q), .D(T11884_Y), .RN(T15030_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T522 ( .Q(T522_Q), .D(T7813_Y), .RN(T15030_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T523 ( .Q(T523_Q), .D(T357_Y), .RN(T14985_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T524 ( .Q(T524_Q), .D(T11885_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T525 ( .Q(T525_Q), .D(T11196_Y), .RN(T15030_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T526 ( .Q(T526_Q), .D(T10264_Y), .RN(T15030_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T528 ( .Q(T528_Q), .D(T11891_Y), .RN(T15030_Y),     .CK(T13936_Q));
KC_DFFRNHQ_X2 T529 ( .Q(T529_Q), .D(T11220_Y), .RN(T15030_Y),     .CK(T14094_Q));
KC_DFFRNHQ_X2 T530 ( .Q(T530_Q), .D(T11224_Y), .RN(T15030_Y),     .CK(T14094_Q));
KC_DFFRNHQ_X2 T541 ( .Q(T541_Q), .D(T11240_Y), .RN(T14973_Y),     .CK(T14200_Q));
KC_DFFRNHQ_X2 T543 ( .Q(T543_Q), .D(T11231_Y), .RN(T14997_Y),     .CK(T14096_Q));
KC_DFFRNHQ_X2 T544 ( .Q(T544_Q), .D(T11229_Y), .RN(T14997_Y),     .CK(T14096_Q));
KC_DFFRNHQ_X2 T550 ( .Q(T550_Q), .D(T11219_Y), .RN(T15030_Y),     .CK(T14094_Q));
KC_DFFRNHQ_X2 T551 ( .Q(T551_Q), .D(T11241_Y), .RN(T14973_Y),     .CK(T14200_Q));
KC_DFFRNHQ_X2 T556 ( .Q(T556_Q), .D(T8069_Y), .RN(T14997_Y),     .CK(T14201_Q));
KC_DFFRNHQ_X2 T561 ( .Q(T561_Q), .D(T8124_Y), .RN(T14997_Y),     .CK(T352_Y));
KC_DFFRNHQ_X2 T566 ( .Q(T566_Q), .D(T1256_Y), .RN(T14997_Y),     .CK(T14201_Q));
KC_DFFRNHQ_X2 T567 ( .Q(T567_Q), .D(T16123_Y), .RN(T14997_Y),     .CK(T352_Y));
KC_DFFRNHQ_X2 T572 ( .Q(T572_Q), .D(T8044_Y), .RN(T14997_Y),     .CK(T14201_Q));
KC_DFFRNHQ_X2 T9469 ( .Q(T9469_Q), .D(T11298_Y), .RN(T10535_Y),     .CK(T594_Y));
KC_DFFRNHQ_X2 T604 ( .Q(T604_Q), .D(T11899_Y), .RN(T10535_Y),     .CK(T594_Y));
KC_DFFRNHQ_X2 T605 ( .Q(T605_Q), .D(T9055_Y), .RN(T10535_Y),     .CK(T594_Y));
KC_DFFRNHQ_X2 T606 ( .Q(T606_Q), .D(T11297_Y), .RN(T10535_Y),     .CK(T594_Y));
KC_DFFRNHQ_X2 T621 ( .Q(T621_Q), .D(T11049_Y), .RN(T14973_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T624 ( .Q(T624_Q), .D(T6350_Y), .RN(T15027_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T625 ( .Q(T625_Q), .D(T7607_Y), .RN(T15027_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T626 ( .Q(T626_Q), .D(T7810_Y), .RN(T15027_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T627 ( .Q(T627_Q), .D(T6350_Y), .RN(T15027_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T628 ( .Q(T628_Q), .D(T7810_Y), .RN(T15027_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T630 ( .Q(T630_Q), .D(T7603_Y), .RN(T15027_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T649 ( .Q(T649_Q), .D(T11063_Y), .RN(T14973_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T653 ( .Q(T653_Q), .D(T11848_Y), .RN(T7243_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T657 ( .Q(T657_Q), .D(T11850_Y), .RN(T7243_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T663 ( .Q(T663_Q), .D(T7623_Y), .RN(T7243_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T664 ( .Q(T664_Q), .D(T15028_Y), .RN(T14979_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T665 ( .Q(T665_Q), .D(T7623_Y), .RN(T14979_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T666 ( .Q(T666_Q), .D(T15031_Y), .RN(T14979_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T668 ( .Q(T668_Q), .D(T15031_Y), .RN(T7243_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T669 ( .Q(T669_Q), .D(T7623_Y), .RN(T7243_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T670 ( .Q(T670_Q), .D(T736_Y), .RN(T7243_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T671 ( .Q(T671_Q), .D(T736_Y), .RN(T7243_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T672 ( .Q(T672_Q), .D(T11106_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T674 ( .Q(T674_Q), .D(T736_Y), .RN(T7243_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T676 ( .Q(T676_Q), .D(T16382_Y), .RN(T7243_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T677 ( .Q(T677_Q), .D(T16382_Y), .RN(T7243_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T679 ( .Q(T679_Q), .D(T736_Y), .RN(T7243_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T9340 ( .Q(T9340_Q), .D(T15840_Y), .RN(T14973_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T7367 ( .Q(T7367_Q), .D(T7385_Y), .RN(T14985_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T680 ( .Q(T680_Q), .D(T7623_Y), .RN(T14979_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T681 ( .Q(T681_Q), .D(T11152_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T683 ( .Q(T683_Q), .D(T15722_Y), .RN(T14985_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T687 ( .Q(T687_Q), .D(T15839_Y), .RN(T14985_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T688 ( .Q(T688_Q), .D(T7385_Y), .RN(T14985_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T689 ( .Q(T689_Q), .D(T15722_Y), .RN(T14985_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T690 ( .Q(T690_Q), .D(T7385_Y), .RN(T14973_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T694 ( .Q(T694_Q), .D(T15031_Y), .RN(T14979_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T695 ( .Q(T695_Q), .D(T15839_Y), .RN(T14973_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T696 ( .Q(T696_Q), .D(T11156_Y), .RN(T14973_Y),     .CK(T923_Y));
KC_DFFRNHQ_X2 T697 ( .Q(T697_Q), .D(T15722_Y), .RN(T14985_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T698 ( .Q(T698_Q), .D(T15722_Y), .RN(T14985_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T699 ( .Q(T699_Q), .D(T11166_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T701 ( .Q(T701_Q), .D(T11182_Y), .RN(T14986_Y),     .CK(T13936_Q));
KC_DFFRNHQ_X2 T705 ( .Q(T705_Q), .D(T15839_Y), .RN(T14973_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T709 ( .Q(T709_Q), .D(T11201_Y), .RN(T15732_Y),     .CK(T923_Y));
KC_DFFRNHQ_X2 T710 ( .Q(T710_Q), .D(T15840_Y), .RN(T14986_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T711 ( .Q(T711_Q), .D(T15839_Y), .RN(T14986_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T712 ( .Q(T712_Q), .D(T15840_Y), .RN(T14973_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T713 ( .Q(T713_Q), .D(T12439_Y), .RN(T14986_Y),     .CK(T13936_Q));
KC_DFFRNHQ_X2 T714 ( .Q(T714_Q), .D(T11212_Y), .RN(T14986_Y),     .CK(T13936_Q));
KC_DFFRNHQ_X2 T716 ( .Q(T716_Q), .D(T11221_Y), .RN(T14986_Y),     .CK(T14094_Q));
KC_DFFRNHQ_X2 T717 ( .Q(T717_Q), .D(T11211_Y), .RN(T14986_Y),     .CK(T14094_Q));
KC_DFFRNHQ_X2 T722 ( .Q(T722_Q), .D(T11216_Y), .RN(T14997_Y),     .CK(T14096_Q));
KC_DFFRNHQ_X2 T724 ( .Q(T724_Q), .D(T11215_Y), .RN(T14986_Y),     .CK(T14096_Q));
KC_DFFRNHQ_X2 T725 ( .Q(T725_Q), .D(T11239_Y), .RN(T14986_Y),     .CK(T14096_Q));
KC_DFFRNHQ_X2 T729 ( .Q(T729_Q), .D(T11228_Y), .RN(T14986_Y),     .CK(T14200_Q));
KC_DFFRNHQ_X2 T741 ( .Q(T741_Q), .D(T11222_Y), .RN(T14986_Y),     .CK(T14094_Q));
KC_DFFRNHQ_X2 T747 ( .Q(T747_Q), .D(T8856_Y), .RN(T14997_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T750 ( .Q(T750_Q), .D(T8857_Y), .RN(T14996_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T751 ( .Q(T751_Q), .D(T8896_Y), .RN(T14997_Y),     .CK(T14201_Q));
KC_DFFRNHQ_X2 T752 ( .Q(T752_Q), .D(T8806_Y), .RN(T14997_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T754 ( .Q(T754_Q), .D(T8806_Y), .RN(T8030_Y),     .CK(T14369_Q));
KC_DFFRNHQ_X2 T760 ( .Q(T760_Q), .D(T8806_Y), .RN(T8030_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T761 ( .Q(T761_Q), .D(T8857_Y), .RN(T14996_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T762 ( .Q(T762_Q), .D(T8856_Y), .RN(T8030_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T765 ( .Q(T765_Q), .D(T8806_Y), .RN(T8030_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T767 ( .Q(T767_Q), .D(T8857_Y), .RN(T14996_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T768 ( .Q(T768_Q), .D(T8856_Y), .RN(T14996_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T9471 ( .Q(T9471_Q), .D(T9985_Y), .RN(T15001_Y),     .CK(T14370_Q));
KC_DFFRNHQ_X2 T9460 ( .Q(T9460_Q), .D(T9985_Y), .RN(T15001_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T769 ( .Q(T769_Q), .D(T10167_Y), .RN(T15001_Y),     .CK(T14370_Q));
KC_DFFRNHQ_X2 T770 ( .Q(T770_Q), .D(T10165_Y), .RN(T15001_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T771 ( .Q(T771_Q), .D(T10165_Y), .RN(T15001_Y),     .CK(T14370_Q));
KC_DFFRNHQ_X2 T772 ( .Q(T772_Q), .D(T10166_Y), .RN(T14997_Y),     .CK(T14370_Q));
KC_DFFRNHQ_X2 T780 ( .Q(T780_Q), .D(T10168_Y), .RN(T15001_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T781 ( .Q(T781_Q), .D(T775_Y), .RN(T10535_Y),     .CK(T14451_Q));
KC_DFFRNHQ_X2 T784 ( .Q(T784_Q), .D(T779_Y), .RN(T10535_Y),     .CK(T14451_Q));
KC_DFFRNHQ_X2 T789 ( .Q(T789_Q), .D(T788_Y), .RN(T10535_Y),     .CK(T14451_Q));
KC_DFFRNHQ_X2 T790 ( .Q(T790_Q), .D(T7603_Y), .RN(T14973_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T793 ( .Q(T793_Q), .D(T15731_Y), .RN(T15026_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T811 ( .Q(T811_Q), .D(T15731_Y), .RN(T15026_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T812 ( .Q(T812_Q), .D(T11854_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T813 ( .Q(T813_Q), .D(T7607_Y), .RN(T15026_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T814 ( .Q(T814_Q), .D(T7603_Y), .RN(T15026_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T815 ( .Q(T815_Q), .D(T11065_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T816 ( .Q(T816_Q), .D(T7607_Y), .RN(T15026_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T817 ( .Q(T817_Q), .D(T11066_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T820 ( .Q(T820_Q), .D(T11059_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T822 ( .Q(T822_Q), .D(T7607_Y), .RN(T15026_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T823 ( .Q(T823_Q), .D(T11056_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T824 ( .Q(T824_Q), .D(T11857_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T825 ( .Q(T825_Q), .D(T15731_Y), .RN(T15026_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T826 ( .Q(T826_Q), .D(T11050_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T828 ( .Q(T828_Q), .D(T11847_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T829 ( .Q(T829_Q), .D(T16382_Y), .RN(T14977_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T831 ( .Q(T831_Q), .D(T7603_Y), .RN(T15026_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T834 ( .Q(T834_Q), .D(T11076_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T838 ( .Q(T838_Q), .D(T11078_Y), .RN(T14977_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T843 ( .Q(T843_Q), .D(T11077_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T847 ( .Q(T847_Q), .D(T11073_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T848 ( .Q(T848_Q), .D(T11072_Y), .RN(T15026_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T860 ( .Q(T860_Q), .D(T11103_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T861 ( .Q(T861_Q), .D(T11093_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T862 ( .Q(T862_Q), .D(T11902_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T863 ( .Q(T863_Q), .D(T11901_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T865 ( .Q(T865_Q), .D(T11859_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T910 ( .Q(T910_Q), .D(T13280_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T935 ( .Q(T935_Q), .D(T11177_Y), .RN(T7798_Y),     .CK(T923_Y));
KC_DFFRNHQ_X2 T938 ( .Q(T938_Q), .D(T8889_Y), .RN(T8030_Y),     .CK(T14202_Q));
KC_DFFRNHQ_X2 T939 ( .Q(T939_Q), .D(T8844_Y), .RN(T8030_Y),     .CK(T14202_Q));
KC_DFFRNHQ_X2 T940 ( .Q(T940_Q), .D(T945_Y), .RN(T8030_Y),     .CK(T14202_Q));
KC_DFFRNHQ_X2 T949 ( .Q(T949_Q), .D(T7875_Y), .RN(T8030_Y),     .CK(T14202_Q));
KC_DFFRNHQ_X2 T963 ( .Q(T963_Q), .D(T8937_Y), .RN(T14996_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T974 ( .Q(T974_Q), .D(T8937_Y), .RN(T8030_Y),     .CK(T4851_Y));
KC_DFFRNHQ_X2 T976 ( .Q(T976_Q), .D(T13257_Y), .RN(T14996_Y),     .CK(T971_Y));
KC_DFFRNHQ_X2 T977 ( .Q(T977_Q), .D(T9413_Y), .RN(T14996_Y),     .CK(T4851_Y));
KC_DFFRNHQ_X2 T978 ( .Q(T978_Q), .D(T9413_Y), .RN(T14996_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T980 ( .Q(T980_Q), .D(T8932_Y), .RN(T8030_Y),     .CK(T16445_Q));
KC_DFFRNHQ_X2 T981 ( .Q(T981_Q), .D(T8887_Y), .RN(T8030_Y),     .CK(T14202_Q));
KC_DFFRNHQ_X2 T982 ( .Q(T982_Q), .D(T12453_Y), .RN(T14996_Y),     .CK(T971_Y));
KC_DFFRNHQ_X2 T983 ( .Q(T983_Q), .D(T9413_Y), .RN(T14996_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T992 ( .Q(T992_Q), .D(T8888_Y), .RN(T8030_Y),     .CK(T14202_Q));
KC_DFFRNHQ_X2 T9459 ( .Q(T9459_Q), .D(T9985_Y), .RN(T15001_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T9458 ( .Q(T9458_Q), .D(T10164_Y), .RN(T15002_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T9457 ( .Q(T9457_Q), .D(T9417_Y), .RN(T15001_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T995 ( .Q(T995_Q), .D(T8858_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T996 ( .Q(T996_Q), .D(T10167_Y), .RN(T15002_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T997 ( .Q(T997_Q), .D(T9417_Y), .RN(T15001_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T998 ( .Q(T998_Q), .D(T10166_Y), .RN(T15001_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T999 ( .Q(T999_Q), .D(T10166_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1000 ( .Q(T1000_Q), .D(T8858_Y), .RN(T15002_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T1001 ( .Q(T1001_Q), .D(T8858_Y), .RN(T14996_Y),     .CK(T4851_Y));
KC_DFFRNHQ_X2 T1002 ( .Q(T1002_Q), .D(T8858_Y), .RN(T14996_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T1003 ( .Q(T1003_Q), .D(T15520_Y), .RN(T15002_Y),     .CK(T14370_Q));
KC_DFFRNHQ_X2 T1004 ( .Q(T1004_Q), .D(T7889_Y), .RN(T14996_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T1005 ( .Q(T1005_Q), .D(T10166_Y), .RN(T15002_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T1012 ( .Q(T1012_Q), .D(T11275_Y), .RN(T15002_Y),     .CK(T971_Y));
KC_DFFRNHQ_X2 T1013 ( .Q(T1013_Q), .D(T7889_Y), .RN(T14996_Y),     .CK(T14369_Q));
KC_DFFRNHQ_X2 T1022 ( .Q(T1022_Q), .D(T5419_Y), .RN(T10535_Y),     .CK(T14451_Q));
KC_DFFRNHQ_X2 T6487 ( .Q(T6487_Q), .D(T11903_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T6486 ( .Q(T6486_Q), .D(T11906_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T1037 ( .Q(T1037_Q), .D(T10343_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1040 ( .Q(T1040_Q), .D(T11141_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1041 ( .Q(T1041_Q), .D(T11164_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1044 ( .Q(T1044_Q), .D(T7359_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1045 ( .Q(T1045_Q), .D(T11162_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1046 ( .Q(T1046_Q), .D(T11163_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1048 ( .Q(T1048_Q), .D(T7550_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T8714 ( .Q(T8714_Q), .D(T11191_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1061 ( .Q(T1061_Q), .D(T8686_Y), .RN(T14993_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1064 ( .Q(T1064_Q), .D(T9818_Y), .RN(T7797_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1065 ( .Q(T1065_Q), .D(T15440_Y), .RN(T7797_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T1066 ( .Q(T1066_Q), .D(T7589_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1067 ( .Q(T1067_Q), .D(T10330_Y), .RN(T7797_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T1068 ( .Q(T1068_Q), .D(T11190_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T1069 ( .Q(T1069_Q), .D(T10330_Y), .RN(T7797_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T1070 ( .Q(T1070_Q), .D(T9816_Y), .RN(T7797_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T1071 ( .Q(T1071_Q), .D(T9819_Y), .RN(T7797_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1072 ( .Q(T1072_Q), .D(T9816_Y), .RN(T7797_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T1073 ( .Q(T1073_Q), .D(T9815_Y), .RN(T7797_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1076 ( .Q(T1076_Q), .D(T9816_Y), .RN(T14993_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T1077 ( .Q(T1077_Q), .D(T16401_Y), .RN(T7797_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T1078 ( .Q(T1078_Q), .D(T8685_Y), .RN(T14993_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1084 ( .Q(T1084_Q), .D(T13279_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T8834 ( .Q(T8834_Q), .D(T8830_Y), .RN(T14993_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T16422 ( .Q(T16422_Q), .D(T1111_Y), .RN(T14993_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T1088 ( .Q(T1088_Q), .D(T10330_Y), .RN(T14993_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T1091 ( .Q(T1091_Q), .D(T10330_Y), .RN(T14993_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T1092 ( .Q(T1092_Q), .D(T15440_Y), .RN(T14993_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T1094 ( .Q(T1094_Q), .D(T13201_Y), .RN(T14993_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1095 ( .Q(T1095_Q), .D(T1093_Y), .RN(T14993_Y),     .CK(T971_Y));
KC_DFFRNHQ_X2 T1100 ( .Q(T1100_Q), .D(T1098_Y), .RN(T14993_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T1113 ( .Q(T1113_Q), .D(T13022_Y), .RN(T14993_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T1121 ( .Q(T1121_Q), .D(T9364_Y), .RN(T14993_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1122 ( .Q(T1122_Q), .D(T9368_Y), .RN(T14993_Y),     .CK(T1074_Y));
KC_DFFRNHQ_X2 T1127 ( .Q(T1127_Q), .D(T9890_Y), .RN(T10697_Y),     .CK(T1140_Y));
KC_DFFRNHQ_X2 T1128 ( .Q(T1128_Q), .D(T13023_Y), .RN(T10697_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T1129 ( .Q(T1129_Q), .D(T13037_Y), .RN(T10697_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T1130 ( .Q(T1130_Q), .D(T8973_Y), .RN(T10697_Y),     .CK(T16445_Q));
KC_DFFRNHQ_X2 T1131 ( .Q(T1131_Q), .D(T8933_Y), .RN(T10697_Y),     .CK(T16445_Q));
KC_DFFRNHQ_X2 T1133 ( .Q(T1133_Q), .D(T9988_Y), .RN(T10697_Y),     .CK(T16445_Q));
KC_DFFRNHQ_X2 T1135 ( .Q(T1135_Q), .D(T13038_Y), .RN(T10697_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T16232 ( .Q(T16232_Q), .D(T10168_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1151 ( .Q(T1151_Q), .D(T16277_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1152 ( .Q(T1152_Q), .D(T10168_Y), .RN(T15002_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T1153 ( .Q(T1153_Q), .D(T10165_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1154 ( .Q(T1154_Q), .D(T10165_Y), .RN(T15002_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T1156 ( .Q(T1156_Q), .D(T10167_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1157 ( .Q(T1157_Q), .D(T15520_Y), .RN(T10727_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T1158 ( .Q(T1158_Q), .D(T15520_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1159 ( .Q(T1159_Q), .D(T10164_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1160 ( .Q(T1160_Q), .D(T9985_Y), .RN(T15002_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T1183 ( .Q(T1183_Q), .D(T12641_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1184 ( .Q(T1184_Q), .D(T12619_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1185 ( .Q(T1185_Q), .D(T12642_Y), .RN(T7797_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1186 ( .Q(T1186_Q), .D(T12620_Y), .RN(T7797_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1187 ( .Q(T1187_Q), .D(T12905_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1188 ( .Q(T1188_Q), .D(T12903_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1189 ( .Q(T1189_Q), .D(T12705_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1190 ( .Q(T1190_Q), .D(T12900_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1191 ( .Q(T1191_Q), .D(T13203_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1195 ( .Q(T1195_Q), .D(T15464_Y), .RN(T15000_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T1202 ( .Q(T1202_Q), .D(T12902_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1203 ( .Q(T1203_Q), .D(T12704_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1204 ( .Q(T1204_Q), .D(T13202_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1207 ( .Q(T1207_Q), .D(T15464_Y), .RN(T14992_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T1208 ( .Q(T1208_Q), .D(T1086_Y), .RN(T14992_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T1209 ( .Q(T1209_Q), .D(T13025_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1210 ( .Q(T1210_Q), .D(T986_Y), .RN(T10697_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T1211 ( .Q(T1211_Q), .D(T1086_Y), .RN(T14992_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T1212 ( .Q(T1212_Q), .D(T15464_Y), .RN(T14992_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T1215 ( .Q(T1215_Q), .D(T12703_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1216 ( .Q(T1216_Q), .D(T16432_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T1220 ( .Q(T1220_Q), .D(T16393_Y), .RN(T15000_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T1221 ( .Q(T1221_Q), .D(T15464_Y), .RN(T14992_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T1222 ( .Q(T1222_Q), .D(T16393_Y), .RN(T15000_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T1223 ( .Q(T1223_Q), .D(T16393_Y), .RN(T15000_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T1224 ( .Q(T1224_Q), .D(T1086_Y), .RN(T14992_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T1231 ( .Q(T1231_Q), .D(T1086_Y), .RN(T15000_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T1232 ( .Q(T1232_Q), .D(T16393_Y), .RN(T15000_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T1247 ( .Q(T1247_Q), .D(T10295_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T1249 ( .Q(T1249_Q), .D(T10296_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T1250 ( .Q(T1250_Q), .D(T10294_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T1264 ( .Q(T1264_Q), .D(T1260_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T1265 ( .Q(T1265_Q), .D(T1258_Y), .RN(T10727_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T1270 ( .Q(T1270_Q), .D(T1263_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T1271 ( .Q(T1271_Q), .D(T1261_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T1283 ( .Q(T1283_Q), .D(T15545_Y), .RN(T1283_RN),     .CK(T5725_Y));
KC_DFFRNHQ_X2 T1361 ( .Q(T1361_Q), .D(T5558_Q), .RN(T13053_SN),     .CK(T16078_Y));
KC_DFFRNHQ_X2 T1660 ( .Q(T1660_Q), .D(T9785_Y), .RN(T1658_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1661 ( .Q(T1661_Q), .D(T809_Y), .RN(T1671_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1662 ( .Q(T1662_Q), .D(T13010_Q), .RN(T2000_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1665 ( .Q(T1665_Q), .D(T4702_Y), .RN(T1664_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1675 ( .Q(T1675_Q), .D(T15048_Y), .RN(T1679_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1678 ( .Q(T1678_Q), .D(T1662_Q), .RN(T2000_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1681 ( .Q(T1681_Q), .D(T4932_Q), .RN(T2000_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1682 ( .Q(T1682_Q), .D(T13009_Q), .RN(T2000_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1690 ( .Q(T1690_Q), .D(T16468_Q), .RN(T14988_Y),     .CK(T16392_Y));
KC_DFFRNHQ_X2 T16435 ( .Q(T16435_Q), .D(T15480_Y), .RN(T1692_Y),     .CK(T16392_Y));
KC_DFFRNHQ_X2 T16434 ( .Q(T16434_Q), .D(T1713_Y), .RN(T14988_Y),     .CK(T14998_Y));
KC_DFFRNHQ_X2 T16433 ( .Q(T16433_Q), .D(T11254_Y), .RN(T15000_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T8880 ( .Q(T8880_Q), .D(T11249_Y), .RN(T15003_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T8877 ( .Q(T8877_Q), .D(T11253_Y), .RN(T15003_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T16413 ( .Q(T16413_Q), .D(T11248_Y), .RN(T15003_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T1691 ( .Q(T1691_Q), .D(T11916_Y), .RN(T15000_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T1694 ( .Q(T1694_Q), .D(T1711_Y), .RN(T4923_Y),     .CK(T16392_Y));
KC_DFFRNHQ_X2 T1707 ( .Q(T1707_Q), .D(T11251_Y), .RN(T15000_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T1714 ( .Q(T1714_Q), .D(T2004_Y), .RN(T2000_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T1717 ( .Q(T1717_Q), .D(T11250_Y), .RN(T15003_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T1719 ( .Q(T1719_Q), .D(T5324_Y), .RN(T1112_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T16306 ( .Q(T16306_Q), .D(T1723_Q), .RN(T14999_Y),     .CK(T16392_Y));
KC_DFFRNHQ_X2 T16297 ( .Q(T16297_Q), .D(T16290_Q), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T16296 ( .Q(T16296_Q), .D(T16297_Q), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T16290 ( .Q(T16290_Q), .D(T1850_Y), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T1723 ( .Q(T1723_Q), .D(T16065_Y), .RN(T14999_Y),     .CK(T16392_Y));
KC_DFFRNHQ_X2 T1725 ( .Q(T1725_Q), .D(T5374_Q), .RN(T14999_Y),     .CK(T16392_Y));
KC_DFFRNHQ_X2 T1726 ( .Q(T1726_Q), .D(T1730_Q), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T1728 ( .Q(T1728_Q), .D(T16475_Y), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T1729 ( .Q(T1729_Q), .D(T16066_Y), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T1730 ( .Q(T1730_Q), .D(T1731_Q), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T1731 ( .Q(T1731_Q), .D(T1835_Y), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T1734 ( .Q(T1734_Q), .D(T16067_Y), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T1735 ( .Q(T1735_Q), .D(T1569_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T1736 ( .Q(T1736_Q), .D(T2488_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T1751 ( .Q(T1751_Q), .D(T2110_Y), .RN(T15011_Y),     .CK(T14554_Q));
KC_DFFRNHQ_X2 T1753 ( .Q(T1753_Q), .D(T2110_Y), .RN(T15011_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X2 T1759 ( .Q(T1759_Q), .D(T2158_Y), .RN(T15011_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X2 T1760 ( .Q(T1760_Q), .D(T5876_Y), .RN(T2169_Y),     .CK(T14565_Q));
KC_DFFRNHQ_X2 T1761 ( .Q(T1761_Q), .D(T20_Y), .RN(T15011_Y),     .CK(T14560_Q));
KC_DFFRNHQ_X2 T1774 ( .Q(T1774_Q), .D(T5063_Y), .RN(T15018_Y),     .CK(T14538_Q));
KC_DFFRNHQ_X2 T1775 ( .Q(T1775_Q), .D(T2213_Y), .RN(T15018_Y),     .CK(T14559_Q));
KC_DFFRNHQ_X2 T1777 ( .Q(T1777_Q), .D(T11596_Y), .RN(T15018_Y),     .CK(T14538_Q));
KC_DFFRNHQ_X2 T1778 ( .Q(T1778_Q), .D(T1776_Y), .RN(T15018_Y),     .CK(T14538_Q));
KC_DFFRNHQ_X2 T1779 ( .Q(T1779_Q), .D(T2214_Y), .RN(T15018_Y),     .CK(T14559_Q));
KC_DFFRNHQ_X2 T1785 ( .Q(T1785_Q), .D(T11601_Y), .RN(T15018_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1787 ( .Q(T1787_Q), .D(T12011_Y), .RN(T15018_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1789 ( .Q(T1789_Q), .D(T11600_Y), .RN(T15018_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1790 ( .Q(T1790_Q), .D(T1783_Y), .RN(T15018_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1803 ( .Q(T1803_Q), .D(T11654_Y), .RN(T15021_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1806 ( .Q(T1806_Q), .D(T11669_Y), .RN(T15018_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1807 ( .Q(T1807_Q), .D(T11653_Y), .RN(T15018_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1820 ( .Q(T1820_Q), .D(T11701_Y), .RN(T15021_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1821 ( .Q(T1821_Q), .D(T11700_Y), .RN(T15021_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1822 ( .Q(T1822_Q), .D(T11691_Y), .RN(T15037_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1823 ( .Q(T1823_Q), .D(T1792_Y), .RN(T15021_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1826 ( .Q(T1826_Q), .D(T1815_Y), .RN(T15037_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1829 ( .Q(T1829_Q), .D(T11690_Y), .RN(T15037_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T1830 ( .Q(T1830_Q), .D(T11753_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T1832 ( .Q(T1832_Q), .D(T6553_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T1833 ( .Q(T1833_Q), .D(T13189_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T1856 ( .Q(T1856_Q), .D(T13195_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T1857 ( .Q(T1857_Q), .D(T13196_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T1970 ( .Q(T1970_Q), .D(T1971_Q), .RN(T14988_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1971 ( .Q(T1971_Q), .D(T4974_Y), .RN(T14988_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1978 ( .Q(T1978_Q), .D(T13012_Q), .RN(T14988_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1981 ( .Q(T1981_Q), .D(T13006_Q), .RN(T14988_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1982 ( .Q(T1982_Q), .D(T13007_Q), .RN(T14988_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T1983 ( .Q(T1983_Q), .D(T1977_Y), .RN(T14988_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T2001 ( .Q(T2001_Q), .D(T2054_Q), .RN(T15003_Y),     .CK(T5725_Y));
KC_DFFRNHQ_X2 T2002 ( .Q(T2002_Q), .D(T11287_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T2005 ( .Q(T2005_Q), .D(T11255_Y), .RN(T1112_Y),     .CK(T14184_Q));
KC_DFFRNHQ_X2 T2008 ( .Q(T2008_Q), .D(T2017_Y), .RN(T1112_Y),     .CK(T14184_Q));
KC_DFFRNHQ_X2 T2012 ( .Q(T2012_Q), .D(T1589_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T2015 ( .Q(T2015_Q), .D(T11256_Y), .RN(T1112_Y),     .CK(T14184_Q));
KC_DFFRNHQ_X2 T2016 ( .Q(T2016_Q), .D(T12713_Y), .RN(T1112_Y),     .CK(T14184_Q));
KC_DFFRNHQ_X2 T2023 ( .Q(T2023_Q), .D(T13030_Y), .RN(T1112_Y),     .CK(T14184_Q));
KC_DFFRNHQ_X2 T2028 ( .Q(T2028_Q), .D(T12709_Y), .RN(T1112_Y),     .CK(T14184_Q));
KC_DFFRNHQ_X2 T2051 ( .Q(T2051_Q), .D(T10084_Y), .RN(T10083_Y),     .CK(T14967_Y));
KC_DFFRNHQ_X2 T2053 ( .Q(T2053_Q), .D(T11288_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T2054 ( .Q(T2054_Q), .D(T5394_Y), .RN(T15003_Y),     .CK(T5725_Y));
KC_DFFRNHQ_X2 T2080 ( .Q(T2080_Q), .D(T2079_Y), .RN(T15806_Q),     .CK(T5725_Y));
KC_DFFRNHQ_X2 T2082 ( .Q(T2082_Q), .D(T10258_Y), .RN(T2063_Y),     .CK(T2078_Y));
KC_DFFRNHQ_X2 T2095 ( .Q(T2095_Q), .D(T2123_Y), .RN(T15008_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T6071 ( .Q(T6071_Q), .D(T15913_Y), .RN(T15011_Y),     .CK(T14570_Q));
KC_DFFRNHQ_X2 T2112 ( .Q(T2112_Q), .D(T15893_Y), .RN(T15011_Y),     .CK(T14570_Q));
KC_DFFRNHQ_X2 T2113 ( .Q(T2113_Q), .D(T2117_Y), .RN(T15011_Y),     .CK(T14559_Q));
KC_DFFRNHQ_X2 T2114 ( .Q(T2114_Q), .D(T16151_Y), .RN(T15013_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X2 T2115 ( .Q(T2115_Q), .D(T15122_Y), .RN(T15013_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T2118 ( .Q(T2118_Q), .D(T15885_Y), .RN(T15011_Y),     .CK(T14570_Q));
KC_DFFRNHQ_X2 T2119 ( .Q(T2119_Q), .D(T15884_Y), .RN(T15011_Y),     .CK(T14570_Q));
KC_DFFRNHQ_X2 T2128 ( .Q(T2128_Q), .D(T13101_Y), .RN(T15008_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X2 T2129 ( .Q(T2129_Q), .D(T2111_Y), .RN(T15011_Y),     .CK(T14559_Q));
KC_DFFRNHQ_X2 T2150 ( .Q(T2150_Q), .D(T15926_Y), .RN(T15015_Y),     .CK(T14565_Q));
KC_DFFRNHQ_X2 T2151 ( .Q(T2151_Q), .D(T11474_Y), .RN(T2169_Y),     .CK(T14558_Q));
KC_DFFRNHQ_X2 T2152 ( .Q(T2152_Q), .D(T2149_Y), .RN(T15015_Y),     .CK(T14570_Q));
KC_DFFRNHQ_X2 T2153 ( .Q(T2153_Q), .D(T13114_Y), .RN(T15015_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X2 T2160 ( .Q(T2160_Q), .D(T11437_Y), .RN(T15011_Y),     .CK(T14558_Q));
KC_DFFRNHQ_X2 T2161 ( .Q(T2161_Q), .D(T13099_Y), .RN(T15013_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T2162 ( .Q(T2162_Q), .D(T11473_Y), .RN(T2169_Y),     .CK(T14558_Q));
KC_DFFRNHQ_X2 T2181 ( .Q(T2181_Q), .D(T2177_Y), .RN(T2169_Y),     .CK(T14559_Q));
KC_DFFRNHQ_X2 T2182 ( .Q(T2182_Q), .D(T2180_Y), .RN(T15015_Y),     .CK(T14559_Q));
KC_DFFRNHQ_X2 T2186 ( .Q(T2186_Q), .D(T5900_Y), .RN(T15015_Y),     .CK(T14565_Q));
KC_DFFRNHQ_X2 T2236 ( .Q(T2236_Q), .D(T12022_Y), .RN(T15018_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X2 T2237 ( .Q(T2237_Q), .D(T11612_Y), .RN(T15018_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X2 T2249 ( .Q(T2249_Q), .D(T5487_Y), .RN(T4047_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X2 T6419 ( .Q(T6419_Q), .D(T12050_Y), .RN(T15021_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2275 ( .Q(T2275_Q), .D(T12010_Y), .RN(T4047_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X2 T2276 ( .Q(T2276_Q), .D(T2821_Y), .RN(T15021_Y),     .CK(T14565_Q));
KC_DFFRNHQ_X2 T2278 ( .Q(T2278_Q), .D(T2262_Y), .RN(T15021_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2281 ( .Q(T2281_Q), .D(T11634_Y), .RN(T4047_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X2 T2311 ( .Q(T2311_Q), .D(T11732_Y), .RN(T15021_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2313 ( .Q(T2313_Q), .D(T2294_Y), .RN(T15037_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2314 ( .Q(T2314_Q), .D(T4948_Y), .RN(T15037_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2315 ( .Q(T2315_Q), .D(T12051_Y), .RN(T15037_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2316 ( .Q(T2316_Q), .D(T2304_Y), .RN(T15037_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2345 ( .Q(T2345_Q), .D(T4950_Y), .RN(T15037_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T2353 ( .Q(T2353_Q), .D(T11754_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T2355 ( .Q(T2355_Q), .D(T11748_Y), .RN(T2322_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T2359 ( .Q(T2359_Q), .D(T15628_Y), .RN(T2322_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T2364 ( .Q(T2364_Q), .D(T6544_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T2381 ( .Q(T2381_Q), .D(T2378_Y), .RN(T2709_Y),     .CK(T14560_Q));
KC_DFFRNHQ_X2 T2385 ( .Q(T2385_Q), .D(T4782_Y), .RN(T2709_Y),     .CK(T14560_Q));
KC_DFFRNHQ_X2 T2388 ( .Q(T2388_Q), .D(T13194_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T2525 ( .Q(T2525_Q), .D(T1983_Q), .RN(T2522_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T2526 ( .Q(T2526_Q), .D(T2525_Q), .RN(T2522_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T2538 ( .Q(T2538_Q), .D(T5319_Y), .RN(T2542_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T2570 ( .Q(T2570_Q), .D(T6692_Y), .RN(T1112_Y),     .CK(T14185_Q));
KC_DFFRNHQ_X2 T2571 ( .Q(T2571_Q), .D(T3153_Y), .RN(T1112_Y),     .CK(T14185_Q));
KC_DFFRNHQ_X2 T2572 ( .Q(T2572_Q), .D(T2588_Y), .RN(T2582_Y),     .CK(T14326_Q));
KC_DFFRNHQ_X2 T2575 ( .Q(T2575_Q), .D(T16362_Y), .RN(T1112_Y),     .CK(T14185_Q));
KC_DFFRNHQ_X2 T2583 ( .Q(T2583_Q), .D(T11282_Y), .RN(T1112_Y),     .CK(T14185_Q));
KC_DFFRNHQ_X2 T2584 ( .Q(T2584_Q), .D(T13289_Y), .RN(T1112_Y),     .CK(T14185_Q));
KC_DFFRNHQ_X2 T2591 ( .Q(T2591_Q), .D(T1141_Y), .RN(T2582_Y),     .CK(T14326_Q));
KC_DFFRNHQ_X2 T2592 ( .Q(T2592_Q), .D(T9948_Y), .RN(T2582_Y),     .CK(T14326_Q));
KC_DFFRNHQ_X2 T2625 ( .Q(T2625_Q), .D(T10089_Y), .RN(T2063_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T2626 ( .Q(T2626_Q), .D(T12740_Y), .RN(T1112_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T2627 ( .Q(T2627_Q), .D(T12943_Y), .RN(T1112_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T2628 ( .Q(T2628_Q), .D(T10077_Y), .RN(T1112_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T2631 ( .Q(T2631_Q), .D(T12733_Y), .RN(T1112_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T2639 ( .Q(T2639_Q), .D(T5731_Y), .RN(T2062_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T2669 ( .Q(T2669_Q), .D(T6707_Y), .RN(T2062_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T2689 ( .Q(T2689_Q), .D(T11017_Y), .RN(T15008_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X2 T2692 ( .Q(T2692_Q), .D(T15850_Y), .RN(T15008_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T2710 ( .Q(T2710_Q), .D(T12169_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T2711 ( .Q(T2711_Q), .D(T12175_Y), .RN(T15013_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T2713 ( .Q(T2713_Q), .D(T12170_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T2715 ( .Q(T2715_Q), .D(T12162_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T2716 ( .Q(T2716_Q), .D(T12161_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T2735 ( .Q(T2735_Q), .D(T10930_Y), .RN(T15013_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2737 ( .Q(T2737_Q), .D(T6153_Y), .RN(T15013_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2738 ( .Q(T2738_Q), .D(T6154_Y), .RN(T15013_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2746 ( .Q(T2746_Q), .D(T10929_Y), .RN(T15013_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2748 ( .Q(T2748_Q), .D(T6152_Y), .RN(T15013_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2749 ( .Q(T2749_Q), .D(T6736_Y), .RN(T15013_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2752 ( .Q(T2752_Q), .D(T8211_Y), .RN(T15013_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2759 ( .Q(T2759_Q), .D(T15960_Y), .RN(VDD),     .CK(T2790_Y));
KC_DFFRNHQ_X2 T2793 ( .Q(T2793_Q), .D(T2794_Q), .RN(T2808_Y),     .CK(T2790_Y));
KC_DFFRNHQ_X2 T2794 ( .Q(T2794_Q), .D(T11547_Y), .RN(T2808_Y),     .CK(T2790_Y));
KC_DFFRNHQ_X2 T2814 ( .Q(T2814_Q), .D(T5997_Y), .RN(T4047_Y),     .CK(T14570_Q));
KC_DFFRNHQ_X2 T2815 ( .Q(T2815_Q), .D(T8472_Y), .RN(T15020_Y),     .CK(T5725_Y));
KC_DFFRNHQ_X2 T2832 ( .Q(T2832_Q), .D(T2834_Y), .RN(T2081_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T2833 ( .Q(T2833_Q), .D(T11649_Y), .RN(T2081_Y),     .CK(T14570_Q));
KC_DFFRNHQ_X2 T2835 ( .Q(T2835_Q), .D(T2826_Y), .RN(T15021_Y),     .CK(T14961_Q));
KC_DFFRNHQ_X2 T2841 ( .Q(T2841_Q), .D(T12967_Y), .RN(T2081_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T2842 ( .Q(T2842_Q), .D(T2845_Y), .RN(T15020_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T2843 ( .Q(T2843_Q), .D(T11648_Y), .RN(T4047_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X2 T2874 ( .Q(T2874_Q), .D(T8387_Y), .RN(T15021_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T2878 ( .Q(T2878_Q), .D(T11718_Y), .RN(T15021_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T2942 ( .Q(T2942_Q), .D(T12068_Y), .RN(T15023_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T2943 ( .Q(T2943_Q), .D(T6488_Y), .RN(T15023_Y),     .CK(T14582_Q));
KC_DFFRNHQ_X2 T2944 ( .Q(T2944_Q), .D(T2946_Y), .RN(T15023_Y),     .CK(T14582_Q));
KC_DFFRNHQ_X2 T2945 ( .Q(T2945_Q), .D(T13193_Y), .RN(T15023_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T2949 ( .Q(T2949_Q), .D(T8153_Y), .RN(T15023_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T2952 ( .Q(T2952_Q), .D(T12296_Y), .RN(T2709_Y),     .CK(T3496_Y));
KC_DFFRNHQ_X2 T2953 ( .Q(T2953_Q), .D(T11819_Y), .RN(T15023_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T2954 ( .Q(T2954_Q), .D(T11820_Y), .RN(T2709_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T2955 ( .Q(T2955_Q), .D(T2940_Y), .RN(T2709_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T3213 ( .Q(T3213_Q), .D(T12146_Y), .RN(T3221_Y),     .CK(T3209_Y));
KC_DFFRNHQ_X2 T3218 ( .Q(T3218_Q), .D(T12793_Y), .RN(T3221_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T3226 ( .Q(T3226_Q), .D(T12179_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T3227 ( .Q(T3227_Q), .D(T12177_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T3228 ( .Q(T3228_Q), .D(T12171_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T3242 ( .Q(T3242_Q), .D(T10257_Y), .RN(T15009_Y),     .CK(T3209_Y));
KC_DFFRNHQ_X2 T3244 ( .Q(T3244_Q), .D(T12152_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T3245 ( .Q(T3245_Q), .D(T12154_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T3246 ( .Q(T3246_Q), .D(T12176_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T3256 ( .Q(T3256_Q), .D(T3273_Y), .RN(T15034_Y),     .CK(T3264_Y));
KC_DFFRNHQ_X2 T3257 ( .Q(T3257_Q), .D(T3276_Y), .RN(T15034_Y),     .CK(T3264_Y));
KC_DFFRNHQ_X2 T3258 ( .Q(T3258_Q), .D(T12339_Y), .RN(T869_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T3412 ( .Q(T3412_Q), .D(T13162_Y), .RN(T15020_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T3519 ( .Q(T3519_Q), .D(T11798_Y), .RN(T15023_Y),     .CK(T14579_Q));
KC_DFFRNHQ_X2 T3520 ( .Q(T3520_Q), .D(T13190_Y), .RN(T15023_Y),     .CK(T14579_Q));
KC_DFFRNHQ_X2 T3521 ( .Q(T3521_Q), .D(T11689_Y), .RN(T15023_Y),     .CK(T14579_Q));
KC_DFFRNHQ_X2 T3522 ( .Q(T3522_Q), .D(T3470_Y), .RN(T15023_Y),     .CK(T14579_Q));
KC_DFFRNHQ_X2 T3523 ( .Q(T3523_Q), .D(T11799_Y), .RN(T15023_Y),     .CK(T14579_Q));
KC_DFFRNHQ_X2 T3524 ( .Q(T3524_Q), .D(T8151_Y), .RN(T15023_Y),     .CK(T5725_Y));
KC_DFFRNHQ_X2 T3525 ( .Q(T3525_Q), .D(T12059_Y), .RN(T15023_Y),     .CK(T14579_Q));
KC_DFFRNHQ_X2 T3528 ( .Q(T3528_Q), .D(T3500_Y), .RN(T15023_Y),     .CK(T3496_Y));
KC_DFFRNHQ_X2 T3873 ( .Q(T3873_Q), .D(T10634_Y), .RN(T3888_Y),     .CK(T14562_Q));
KC_DFFRNHQ_X2 T3877 ( .Q(T3877_Q), .D(T3875_Y), .RN(T869_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T3878 ( .Q(T3878_Q), .D(T3891_Y), .RN(T869_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T3883 ( .Q(T3883_Q), .D(T3881_Y), .RN(T3888_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T3884 ( .Q(T3884_Q), .D(T8229_Y), .RN(T869_Y),     .CK(T14562_Q));
KC_DFFRNHQ_X2 T3885 ( .Q(T3885_Q), .D(T15932_Y), .RN(T3888_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T3889 ( .Q(T3889_Q), .D(T8222_Y), .RN(T869_Y),     .CK(T14562_Q));
KC_DFFRNHQ_X2 T3890 ( .Q(T3890_Q), .D(T15931_Y), .RN(T869_Y),     .CK(T14562_Q));
KC_DFFRNHQ_X2 T3895 ( .Q(T3895_Q), .D(T3894_Y), .RN(T869_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T3900 ( .Q(T3900_Q), .D(T3893_Y), .RN(T3888_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T3935 ( .Q(T3935_Q), .D(T8255_Y), .RN(T3888_Y),     .CK(T3879_Y));
KC_DFFRNHQ_X2 T3936 ( .Q(T3936_Q), .D(T8256_Y), .RN(T3888_Y),     .CK(T3879_Y));
KC_DFFRNHQ_X2 T3937 ( .Q(T3937_Q), .D(T15576_Y), .RN(T3888_Y),     .CK(T3879_Y));
KC_DFFRNHQ_X2 T3964 ( .Q(T3964_Q), .D(T3948_Y), .RN(T15016_Y),     .CK(T14567_Q));
KC_DFFRNHQ_X2 T3965 ( .Q(T3965_Q), .D(T12225_Y), .RN(T15016_Y),     .CK(T14567_Q));
KC_DFFRNHQ_X2 T3968 ( .Q(T3968_Q), .D(T12226_Y), .RN(T15016_Y),     .CK(T14567_Q));
KC_DFFRNHQ_X2 T3970 ( .Q(T3970_Q), .D(T3969_Y), .RN(T5023_Y),     .CK(T3993_Y));
KC_DFFRNHQ_X2 T3971 ( .Q(T3971_Q), .D(T12214_Y), .RN(T5023_Y),     .CK(T3993_Y));
KC_DFFRNHQ_X2 T3974 ( .Q(T3974_Q), .D(T11543_Y), .RN(T15016_Y),     .CK(T14567_Q));
KC_DFFRNHQ_X2 T3990 ( .Q(T3990_Q), .D(T3989_Y), .RN(T5023_Y),     .CK(T3993_Y));
KC_DFFRNHQ_X2 T4006 ( .Q(T4006_Q), .D(T3997_Y), .RN(T5023_Y),     .CK(T3993_Y));
KC_DFFRNHQ_X2 T4043 ( .Q(T4043_Q), .D(T4679_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4044 ( .Q(T4044_Q), .D(T12964_Y), .RN(T15035_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T4048 ( .Q(T4048_Q), .D(T16210_Y), .RN(T15035_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T4050 ( .Q(T4050_Q), .D(T4038_Y), .RN(T15035_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T4051 ( .Q(T4051_Q), .D(T11635_Y), .RN(T15035_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T4052 ( .Q(T4052_Q), .D(T12841_Y), .RN(T15035_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X2 T4056 ( .Q(T4056_Q), .D(T4680_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4147 ( .Q(T4147_Q), .D(T4108_Y), .RN(T4047_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X2 T4163 ( .Q(T4163_Q), .D(T11003_Y), .RN(T15023_Y),     .CK(T14580_Q));
KC_DFFRNHQ_X2 T4164 ( .Q(T4164_Q), .D(T11841_Y), .RN(T15023_Y),     .CK(T14580_Q));
KC_DFFRNHQ_X2 T4168 ( .Q(T4168_Q), .D(T3507_Y), .RN(T15023_Y),     .CK(T14580_Q));
KC_DFFRNHQ_X2 T4169 ( .Q(T4169_Q), .D(T4170_Y), .RN(T15023_Y),     .CK(T14580_Q));
KC_DFFRNHQ_X2 T4171 ( .Q(T4171_Q), .D(T6528_Y), .RN(T15023_Y),     .CK(T14580_Q));
KC_DFFRNHQ_X2 T4178 ( .Q(T4178_Q), .D(T8513_Y), .RN(T4047_Y),     .CK(T3496_Y));
KC_DFFRNHQ_X2 T4351 ( .Q(T4351_Q), .D(T5171_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4359 ( .Q(T4359_Q), .D(T4373_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4360 ( .Q(T4360_Q), .D(T4378_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4361 ( .Q(T4361_Q), .D(T4355_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4362 ( .Q(T4362_Q), .D(T4357_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4363 ( .Q(T4363_Q), .D(T4365_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4367 ( .Q(T4367_Q), .D(T5172_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4368 ( .Q(T4368_Q), .D(T4371_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4369 ( .Q(T4369_Q), .D(T12116_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4370 ( .Q(T4370_Q), .D(T4372_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4374 ( .Q(T4374_Q), .D(T4366_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4375 ( .Q(T4375_Q), .D(T4364_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4376 ( .Q(T4376_Q), .D(T4379_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4380 ( .Q(T4380_Q), .D(T4377_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4381 ( .Q(T4381_Q), .D(T4356_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4406 ( .Q(T4406_Q), .D(T4358_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4427 ( .Q(T4427_Q), .D(T5166_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T4454 ( .Q(T4454_Q), .D(T4442_Y), .RN(T4402_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T4455 ( .Q(T4455_Q), .D(T6099_Y), .RN(T4402_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T4456 ( .Q(T4456_Q), .D(T4433_Y), .RN(T4402_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T4465 ( .Q(T4465_Q), .D(T8200_Y), .RN(T4402_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T4484 ( .Q(T4484_Q), .D(T6218_Y), .RN(T3888_Y),     .CK(T14561_Q));
KC_DFFRNHQ_X2 T4487 ( .Q(T4487_Q), .D(T11418_Y), .RN(T4402_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T4490 ( .Q(T4490_Q), .D(T15937_Y), .RN(T3888_Y),     .CK(T14561_Q));
KC_DFFRNHQ_X2 T4491 ( .Q(T4491_Q), .D(T5453_Y), .RN(T3888_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T4492 ( .Q(T4492_Q), .D(T8220_Y), .RN(T3888_Y),     .CK(T14561_Q));
KC_DFFRNHQ_X2 T4493 ( .Q(T4493_Q), .D(T4496_Y), .RN(T3888_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T4498 ( .Q(T4498_Q), .D(T11452_Y), .RN(T3888_Y),     .CK(T14561_Q));
KC_DFFRNHQ_X2 T4526 ( .Q(T4526_Q), .D(T4512_Y), .RN(T3888_Y),     .CK(T14569_Q));
KC_DFFRNHQ_X2 T4527 ( .Q(T4527_Q), .D(T11508_Y), .RN(T3888_Y),     .CK(T14569_Q));
KC_DFFRNHQ_X2 T4528 ( .Q(T4528_Q), .D(T12193_Y), .RN(T3888_Y),     .CK(T14569_Q));
KC_DFFRNHQ_X2 T4537 ( .Q(T4537_Q), .D(T8243_Y), .RN(T3888_Y),     .CK(T14561_Q));
KC_DFFRNHQ_X2 T4568 ( .Q(T4568_Q), .D(T12351_Y), .RN(T15016_Y),     .CK(T14569_Q));
KC_DFFRNHQ_X2 T4572 ( .Q(T4572_Q), .D(T8284_Y), .RN(T15016_Y),     .CK(T14568_Q));
KC_DFFRNHQ_X2 T4573 ( .Q(T4573_Q), .D(T4574_Y), .RN(T15016_Y),     .CK(T14568_Q));
KC_DFFRNHQ_X2 T4575 ( .Q(T4575_Q), .D(T8291_Y), .RN(T15016_Y),     .CK(T14568_Q));
KC_DFFRNHQ_X2 T4576 ( .Q(T4576_Q), .D(T11589_Y), .RN(T15016_Y),     .CK(T14568_Q));
KC_DFFRNHQ_X2 T4578 ( .Q(T4578_Q), .D(T6261_Y), .RN(T15016_Y),     .CK(T14568_Q));
KC_DFFRNHQ_X2 T4579 ( .Q(T4579_Q), .D(T8288_Y), .RN(T15016_Y),     .CK(T14568_Q));
KC_DFFRNHQ_X2 T4602 ( .Q(T4602_Q), .D(T4603_Y), .RN(T15016_Y),     .CK(T14958_Q));
KC_DFFRNHQ_X2 T4606 ( .Q(T4606_Q), .D(T6242_Y), .RN(T15016_Y),     .CK(T14958_Q));
KC_DFFRNHQ_X2 T4607 ( .Q(T4607_Q), .D(T4604_Y), .RN(T15016_Y),     .CK(T14958_Q));
KC_DFFRNHQ_X2 T4608 ( .Q(T4608_Q), .D(T8475_Y), .RN(T15016_Y),     .CK(T14958_Q));
KC_DFFRNHQ_X2 T4626 ( .Q(T4626_Q), .D(T8304_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T4627 ( .Q(T4627_Q), .D(T8301_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T4628 ( .Q(T4628_Q), .D(T8303_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T4629 ( .Q(T4629_Q), .D(T8464_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T4630 ( .Q(T4630_Q), .D(T8302_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T4663 ( .Q(T4663_Q), .D(T12840_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4669 ( .Q(T4669_Q), .D(T6056_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4675 ( .Q(T4675_Q), .D(T16062_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4685 ( .Q(T4685_Q), .D(T4677_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4686 ( .Q(T4686_Q), .D(T4670_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4693 ( .Q(T4693_Q), .D(T12839_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4713 ( .Q(T4713_Q), .D(T10613_Y), .RN(T15022_Y),     .CK(T4728_Y));
KC_DFFRNHQ_X2 T4714 ( .Q(T4714_Q), .D(T16059_Y), .RN(T15022_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T4717 ( .Q(T4717_Q), .D(T12850_Y), .RN(T15022_Y),     .CK(T4728_Y));
KC_DFFRNHQ_X2 T4718 ( .Q(T4718_Q), .D(T6129_Y), .RN(T15022_Y),     .CK(T2667_Y));
KC_DFFRNHQ_X2 T4719 ( .Q(T4719_Q), .D(T10600_Y), .RN(T15022_Y),     .CK(T4728_Y));
KC_DFFRNHQ_X2 T4720 ( .Q(T4720_Q), .D(T12260_Y), .RN(T15022_Y),     .CK(T4728_Y));
KC_DFFRNHQ_X2 T4721 ( .Q(T4721_Q), .D(T8379_Y), .RN(T15022_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T4722 ( .Q(T4722_Q), .D(T12261_Y), .RN(T15022_Y),     .CK(T4728_Y));
KC_DFFRNHQ_X2 T4723 ( .Q(T4723_Q), .D(T11681_Y), .RN(T15022_Y),     .CK(T4728_Y));
KC_DFFRNHQ_X2 T4746 ( .Q(T4746_Q), .D(T11785_Y), .RN(T15022_Y),     .CK(T4728_Y));
KC_DFFRNHQ_X2 T4750 ( .Q(T4750_Q), .D(T4745_Y), .RN(T15022_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T4755 ( .Q(T4755_Q), .D(T13185_Y), .RN(T15022_Y),     .CK(T14578_Q));
KC_DFFRNHQ_X2 T4756 ( .Q(T4756_Q), .D(T11759_Y), .RN(T15020_Y),     .CK(T14578_Q));
KC_DFFRNHQ_X2 T4757 ( .Q(T4757_Q), .D(T4751_Y), .RN(T15022_Y),     .CK(T14578_Q));
KC_DFFRNHQ_X2 T4758 ( .Q(T4758_Q), .D(T6548_Y), .RN(T15020_Y),     .CK(T14578_Q));
KC_DFFRNHQ_X2 T4759 ( .Q(T4759_Q), .D(T11733_Y), .RN(T15020_Y),     .CK(T14578_Q));
KC_DFFRNHQ_X2 T4760 ( .Q(T4760_Q), .D(T4753_Y), .RN(T15020_Y),     .CK(T14578_Q));
KC_DFFRNHQ_X2 T4799 ( .Q(T4799_Q), .D(T15028_Y), .RN(T15029_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T4802 ( .Q(T4802_Q), .D(T227_Y), .RN(T7675_Y),     .CK(T4828_Y));
KC_DFFRNHQ_X2 T4803 ( .Q(T4803_Q), .D(T16315_Y), .RN(T14976_Y),     .CK(T14589_Q));
KC_DFFRNHQ_X2 T4810 ( .Q(T4810_Q), .D(T176_Y), .RN(T14978_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T9351 ( .Q(T9351_Q), .D(T7813_Y), .RN(T15029_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T9350 ( .Q(T9350_Q), .D(T11883_Y), .RN(T15030_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T9349 ( .Q(T9349_Q), .D(T11147_Y), .RN(T15030_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T4822 ( .Q(T4822_Q), .D(T11075_Y), .RN(T14975_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T4823 ( .Q(T4823_Q), .D(T11088_Y), .RN(T14978_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T9472 ( .Q(T9472_Q), .D(T12889_Y), .RN(T10535_Y),     .CK(T594_Y));
KC_DFFRNHQ_X2 T4827 ( .Q(T4827_Q), .D(T11889_Y), .RN(T15030_Y),     .CK(T13936_Q));
KC_DFFRNHQ_X2 T4835 ( .Q(T4835_Q), .D(T11852_Y), .RN(T7242_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T4836 ( .Q(T4836_Q), .D(T15031_Y), .RN(T14979_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T4837 ( .Q(T4837_Q), .D(T15028_Y), .RN(T14979_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T4840 ( .Q(T4840_Q), .D(T11223_Y), .RN(T14986_Y),     .CK(T14094_Q));
KC_DFFRNHQ_X2 T4843 ( .Q(T4843_Q), .D(T9417_Y), .RN(T14997_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T4845 ( .Q(T4845_Q), .D(T11851_Y), .RN(T7243_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T4846 ( .Q(T4846_Q), .D(T11849_Y), .RN(T7243_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T9456 ( .Q(T9456_Q), .D(T1015_Y), .RN(T15002_Y),     .CK(T971_Y));
KC_DFFRNHQ_X2 T4854 ( .Q(T4854_Q), .D(T11091_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T4855 ( .Q(T4855_Q), .D(T16382_Y), .RN(T14977_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T4858 ( .Q(T4858_Q), .D(T9327_Y), .RN(T7740_Y),     .CK(T1047_Y));
KC_DFFRNHQ_X2 T4860 ( .Q(T4860_Q), .D(T9816_Y), .RN(T14993_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T4861 ( .Q(T4861_Q), .D(T16401_Y), .RN(T14993_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T4862 ( .Q(T4862_Q), .D(T16277_Y), .RN(T15002_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T4869 ( .Q(T4869_Q), .D(T12901_Y), .RN(T14992_Y),     .CK(T1115_Y));
KC_DFFRNHQ_X2 T4925 ( .Q(T4925_Q), .D(T1816_Y), .RN(T15037_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T4930 ( .Q(T4930_Q), .D(T1757_Y), .RN(T15011_Y),     .CK(T14960_Q));
KC_DFFRNHQ_X2 T4932 ( .Q(T4932_Q), .D(T2021_Y), .RN(T2000_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T4964 ( .Q(T4964_Q), .D(T2301_Y), .RN(T15037_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T4967 ( .Q(T4967_Q), .D(T2187_Y), .RN(T15015_Y),     .CK(T14559_Q));
KC_DFFRNHQ_X2 T4969 ( .Q(T4969_Q), .D(T2126_Y), .RN(T15008_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T4970 ( .Q(T4970_Q), .D(T2159_Y), .RN(T2169_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T4971 ( .Q(T4971_Q), .D(T13100_Y), .RN(T15013_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T5015 ( .Q(T5015_Q), .D(T10895_Y), .RN(T2688_Y),     .CK(T3209_Y));
KC_DFFRNHQ_X2 T5016 ( .Q(T5016_Q), .D(T15231_Y), .RN(T2688_Y),     .CK(T3879_Y));
KC_DFFRNHQ_X2 T5018 ( .Q(T5018_Q), .D(T11008_Y), .RN(T2688_Y),     .CK(T14497_Q));
KC_DFFRNHQ_X2 T5025 ( .Q(T5025_Q), .D(T16094_Y), .RN(T2582_Y),     .CK(T14326_Q));
KC_DFFRNHQ_X2 T5027 ( .Q(T5027_Q), .D(T2526_Q), .RN(T2522_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T5074 ( .Q(T5074_Q), .D(T15862_Y), .RN(T15009_Y),     .CK(T3209_Y));
KC_DFFRNHQ_X2 T5075 ( .Q(T5075_Q), .D(T12153_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T5076 ( .Q(T5076_Q), .D(T12338_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T5129 ( .Q(T5129_Q), .D(T3874_Y), .RN(T869_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T5130 ( .Q(T5130_Q), .D(T3892_Y), .RN(T869_Y),     .CK(T14555_Q));
KC_DFFRNHQ_X2 T5158 ( .Q(T5158_Q), .D(T8474_Y), .RN(T15016_Y),     .CK(T14958_Q));
KC_DFFRNHQ_X2 T5159 ( .Q(T5159_Q), .D(T15993_Y), .RN(T15016_Y),     .CK(T14958_Q));
KC_DFFRNHQ_X2 T5162 ( .Q(T5162_Q), .D(T8463_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T5164 ( .Q(T5164_Q), .D(T15899_Y), .RN(T4402_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T5165 ( .Q(T5165_Q), .D(T8203_Y), .RN(T4402_Y),     .CK(T14542_Q));
KC_DFFRNHQ_X2 T5170 ( .Q(T5170_Q), .D(T5167_Y), .RN(T15033_Y),     .CK(T4350_Y));
KC_DFFRNHQ_X2 T5184 ( .Q(T5184_Q), .D(T71_Y), .RN(T15024_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T5185 ( .Q(T5185_Q), .D(T12372_Y), .RN(T15024_Y),     .CK(T16477_Y));
KC_DFFRNHQ_X2 T5187 ( .Q(T5187_Q), .D(T62_Y), .RN(T15024_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T5189 ( .Q(T5189_Q), .D(T5591_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T5190 ( .Q(T5190_Q), .D(T51_Y), .RN(T14970_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T5192 ( .Q(T5192_Q), .D(T8595_Y), .RN(T7074_Y),     .CK(T130_Y));
KC_DFFRNHQ_X2 T5193 ( .Q(T5193_Q), .D(T11055_Y), .RN(T14974_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T5194 ( .Q(T5194_Q), .D(T11053_Y), .RN(T15027_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T5195 ( .Q(T5195_Q), .D(T6350_Y), .RN(T14973_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T5196 ( .Q(T5196_Q), .D(T6809_Y), .RN(T14974_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T5198 ( .Q(T5198_Q), .D(T7810_Y), .RN(T15027_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T5199 ( .Q(T5199_Q), .D(T15731_Y), .RN(T14973_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T5200 ( .Q(T5200_Q), .D(T7318_Y), .RN(T15027_Y),     .CK(T644_Y));
KC_DFFRNHQ_X2 T5202 ( .Q(T5202_Q), .D(T8551_Y), .RN(T7074_Y),     .CK(T13330_Q));
KC_DFFRNHQ_X2 T5203 ( .Q(T5203_Q), .D(T5597_Y), .RN(T7074_Y),     .CK(T13330_Q));
KC_DFFRNHQ_X2 T5204 ( .Q(T5204_Q), .D(T472_Y), .RN(T14974_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T5205 ( .Q(T5205_Q), .D(T7810_Y), .RN(T15027_Y),     .CK(T5197_Y));
KC_DFFRNHQ_X2 T5206 ( .Q(T5206_Q), .D(T6350_Y), .RN(T15027_Y),     .CK(T846_Y));
KC_DFFRNHQ_X2 T5220 ( .Q(T5220_Q), .D(T9254_Y), .RN(T15024_Y),     .CK(T13331_Q));
KC_DFFRNHQ_X2 T5221 ( .Q(T5221_Q), .D(T11856_Y), .RN(T7242_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T5222 ( .Q(T5222_Q), .D(T6967_Y), .RN(T7073_Y),     .CK(T130_Y));
KC_DFFRNHQ_X2 T5223 ( .Q(T5223_Q), .D(T11067_Y), .RN(T15027_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T5225 ( .Q(T5225_Q), .D(T6909_Y), .RN(T7073_Y),     .CK(T130_Y));
KC_DFFRNHQ_X2 T5226 ( .Q(T5226_Q), .D(T11070_Y), .RN(T14974_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T5227 ( .Q(T5227_Q), .D(T11069_Y), .RN(T15027_Y),     .CK(T226_Y));
KC_DFFRNHQ_X2 T5229 ( .Q(T5229_Q), .D(T808_Y), .RN(T14973_Y),     .CK(T810_Y));
KC_DFFRNHQ_X2 T7085 ( .Q(T7085_Q), .D(T7108_Y), .RN(T14975_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T5237 ( .Q(T5237_Q), .D(T11089_Y), .RN(T869_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T5238 ( .Q(T5238_Q), .D(T11102_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T5239 ( .Q(T5239_Q), .D(T11084_Y), .RN(T14975_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T5240 ( .Q(T5240_Q), .D(T11080_Y), .RN(T7242_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T5241 ( .Q(T5241_Q), .D(T11081_Y), .RN(T7242_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T5242 ( .Q(T5242_Q), .D(T156_Y), .RN(T14975_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T5243 ( .Q(T5243_Q), .D(T156_Y), .RN(T14975_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T5251 ( .Q(T5251_Q), .D(T11911_Y), .RN(T14978_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T5252 ( .Q(T5252_Q), .D(T15028_Y), .RN(T14979_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T5253 ( .Q(T5253_Q), .D(T7812_Y), .RN(T14979_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T5254 ( .Q(T5254_Q), .D(T11910_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T5255 ( .Q(T5255_Q), .D(T11108_Y), .RN(T14978_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T5257 ( .Q(T5257_Q), .D(T11094_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T5258 ( .Q(T5258_Q), .D(T1036_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T5259 ( .Q(T5259_Q), .D(T11092_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T5260 ( .Q(T5260_Q), .D(T11095_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T5261 ( .Q(T5261_Q), .D(T11090_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T5262 ( .Q(T5262_Q), .D(T11905_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T5263 ( .Q(T5263_Q), .D(T11099_Y), .RN(T14978_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T5264 ( .Q(T5264_Q), .D(T11904_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T5265 ( .Q(T5265_Q), .D(T11105_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T9355 ( .Q(T9355_Q), .D(T15425_Y), .RN(T15721_Y),     .CK(T503_Y));
KC_DFFRNHQ_X2 T9339 ( .Q(T9339_Q), .D(T7813_Y), .RN(T14985_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T5275 ( .Q(T5275_Q), .D(T11153_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T5276 ( .Q(T5276_Q), .D(T11866_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T5277 ( .Q(T5277_Q), .D(T11150_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T5278 ( .Q(T5278_Q), .D(T15425_Y), .RN(T15029_Y),     .CK(T510_Y));
KC_DFFRNHQ_X2 T5279 ( .Q(T5279_Q), .D(T11158_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T5280 ( .Q(T5280_Q), .D(T7385_Y), .RN(T14985_Y),     .CK(T693_Y));
KC_DFFRNHQ_X2 T5281 ( .Q(T5281_Q), .D(T11149_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T5282 ( .Q(T5282_Q), .D(T11146_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T5283 ( .Q(T5283_Q), .D(T11167_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T5292 ( .Q(T5292_Q), .D(T15440_Y), .RN(T7797_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T5293 ( .Q(T5293_Q), .D(T16401_Y), .RN(T7797_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T5294 ( .Q(T5294_Q), .D(T16401_Y), .RN(T7797_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T5297 ( .Q(T5297_Q), .D(T13277_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T5300 ( .Q(T5300_Q), .D(T15840_Y), .RN(T14986_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T5301 ( .Q(T5301_Q), .D(T7597_Y), .RN(T14986_Y),     .CK(T923_Y));
KC_DFFRNHQ_X2 T5303 ( .Q(T5303_Q), .D(T8808_Y), .RN(T15029_Y),     .CK(T4812_Y));
KC_DFFRNHQ_X2 T5304 ( .Q(T5304_Q), .D(T11169_Y), .RN(T15030_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T5305 ( .Q(T5305_Q), .D(T11881_Y), .RN(T14985_Y),     .CK(T495_Y));
KC_DFFRNHQ_X2 T5306 ( .Q(T5306_Q), .D(T7813_Y), .RN(T14985_Y),     .CK(T686_Y));
KC_DFFRNHQ_X2 T5308 ( .Q(T5308_Q), .D(T7643_Y), .RN(T14986_Y),     .CK(T923_Y));
KC_DFFRNHQ_X2 T5309 ( .Q(T5309_Q), .D(T7562_Y), .RN(T14986_Y),     .CK(T923_Y));
KC_DFFRNHQ_X2 T5310 ( .Q(T5310_Q), .D(T13278_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T5311 ( .Q(T5311_Q), .D(T1681_Q), .RN(T14988_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T5313 ( .Q(T5313_Q), .D(T13015_Q), .RN(T14988_Y),     .CK(T16407_Y));
KC_DFFRNHQ_X2 T5320 ( .Q(T5320_Q), .D(T1976_Y), .RN(T2527_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T5333 ( .Q(T5333_Q), .D(T15440_Y), .RN(T14993_Y),     .CK(T14199_Q));
KC_DFFRNHQ_X2 T5334 ( .Q(T5334_Q), .D(T13200_Y), .RN(T15000_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T5337 ( .Q(T5337_Q), .D(T986_Y), .RN(T10697_Y),     .CK(T14137_Q));
KC_DFFRNHQ_X2 T5340 ( .Q(T5340_Q), .D(T986_Y), .RN(T10697_Y),     .CK(T14113_Q));
KC_DFFRNHQ_X2 T5341 ( .Q(T5341_Q), .D(T986_Y), .RN(T15000_Y),     .CK(T14138_Q));
KC_DFFRNHQ_X2 T5342 ( .Q(T5342_Q), .D(T11225_Y), .RN(T14973_Y),     .CK(T14200_Q));
KC_DFFRNHQ_X2 T5343 ( .Q(T5343_Q), .D(T16439_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T5346 ( .Q(T5346_Q), .D(T7893_Y), .RN(T14997_Y),     .CK(T14200_Q));
KC_DFFRNHQ_X2 T5348 ( .Q(T5348_Q), .D(T11243_Y), .RN(T14986_Y),     .CK(T14200_Q));
KC_DFFRNHQ_X2 T5350 ( .Q(T5350_Q), .D(T11232_Y), .RN(T14986_Y),     .CK(T14200_Q));
KC_DFFRNHQ_X2 T5353 ( .Q(T5353_Q), .D(T8793_Y), .RN(T14993_Y),     .CK(T971_Y));
KC_DFFRNHQ_X2 T5354 ( .Q(T5354_Q), .D(T13284_Y), .RN(T14976_Y),     .CK(T4828_Y));
KC_DFFRNHQ_X2 T5355 ( .Q(T5355_Q), .D(T8813_Y), .RN(T7675_Y),     .CK(T4828_Y));
KC_DFFRNHQ_X2 T5356 ( .Q(T5356_Q), .D(T11226_Y), .RN(T14986_Y),     .CK(T14096_Q));
KC_DFFRNHQ_X2 T5357 ( .Q(T5357_Q), .D(T11242_Y), .RN(T14986_Y),     .CK(T14096_Q));
KC_DFFRNHQ_X2 T5359 ( .Q(T5359_Q), .D(T1696_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T5360 ( .Q(T5360_Q), .D(T16438_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T5362 ( .Q(T5362_Q), .D(T1995_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T5363 ( .Q(T5363_Q), .D(T13039_Y), .RN(T1112_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T5364 ( .Q(T5364_Q), .D(T11261_Y), .RN(T1112_Y),     .CK(T14174_Q));
KC_DFFRNHQ_X2 T5365 ( .Q(T5365_Q), .D(T5906_Y), .RN(T1112_Y),     .CK(T5725_Y));
KC_DFFRNHQ_X2 T5366 ( .Q(T5366_Q), .D(T13031_Q), .RN(T14999_Y),     .CK(T15190_Y));
KC_DFFRNHQ_X2 T5373 ( .Q(T5373_Q), .D(T13035_Y), .RN(T10697_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T5374 ( .Q(T5374_Q), .D(T1728_Q), .RN(T14999_Y),     .CK(T1604_Y));
KC_DFFRNHQ_X2 T5375 ( .Q(T5375_Q), .D(T13036_Y), .RN(T10697_Y),     .CK(T1120_Y));
KC_DFFRNHQ_X2 T5376 ( .Q(T5376_Q), .D(T10300_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T5377 ( .Q(T5377_Q), .D(T8897_Y), .RN(T14997_Y),     .CK(T14201_Q));
KC_DFFRNHQ_X2 T5378 ( .Q(T5378_Q), .D(T8906_Y), .RN(T14997_Y),     .CK(T14201_Q));
KC_DFFRNHQ_X2 T5379 ( .Q(T5379_Q), .D(T8937_Y), .RN(T14996_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T5383 ( .Q(T5383_Q), .D(T9413_Y), .RN(T14996_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T5384 ( .Q(T5384_Q), .D(T8937_Y), .RN(T14996_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T5385 ( .Q(T5385_Q), .D(T7889_Y), .RN(T14996_Y),     .CK(T14216_Q));
KC_DFFRNHQ_X2 T5386 ( .Q(T5386_Q), .D(T8857_Y), .RN(T14996_Y),     .CK(T14369_Q));
KC_DFFRNHQ_X2 T5387 ( .Q(T5387_Q), .D(T7889_Y), .RN(T14996_Y),     .CK(T9048_Q));
KC_DFFRNHQ_X2 T5388 ( .Q(T5388_Q), .D(T15813_Y), .RN(T15003_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T5389 ( .Q(T5389_Q), .D(T11290_Y), .RN(T2063_Y),     .CK(T14304_Q));
KC_DFFRNHQ_X2 T5390 ( .Q(T5390_Q), .D(T11289_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T5391 ( .Q(T5391_Q), .D(T11286_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T5397 ( .Q(T5397_Q), .D(T11283_Y), .RN(T15003_Y),     .CK(T14173_Q));
KC_DFFRNHQ_X2 T9470 ( .Q(T9470_Q), .D(T10168_Y), .RN(T15001_Y),     .CK(T14370_Q));
KC_DFFRNHQ_X2 T9461 ( .Q(T9461_Q), .D(T10164_Y), .RN(T15001_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T5404 ( .Q(T5404_Q), .D(T1259_Y), .RN(T10661_Y),     .CK(T14227_Q));
KC_DFFRNHQ_X2 T5406 ( .Q(T5406_Q), .D(T11300_Y), .RN(T10535_Y),     .CK(T594_Y));
KC_DFFRNHQ_X2 T5407 ( .Q(T5407_Q), .D(T10167_Y), .RN(T15001_Y),     .CK(T14203_Q));
KC_DFFRNHQ_X2 T5408 ( .Q(T5408_Q), .D(T5409_Y), .RN(T2062_Y),     .CK(T2050_Y));
KC_DFFRNHQ_X2 T5416 ( .Q(T5416_Q), .D(T10164_Y), .RN(T15001_Y),     .CK(T14370_Q));
KC_DFFRNHQ_X2 T5417 ( .Q(T5417_Q), .D(T782_Y), .RN(T10535_Y),     .CK(T14451_Q));
KC_DFFRNHQ_X2 T5420 ( .Q(T5420_Q), .D(T787_Y), .RN(T10535_Y),     .CK(T14451_Q));
KC_DFFRNHQ_X2 T5421 ( .Q(T5421_Q), .D(T4996_Y), .RN(T2063_Y),     .CK(T14497_Q));
KC_DFFRNHQ_X2 T5424 ( .Q(T5424_Q), .D(T2679_Y), .RN(T2063_Y),     .CK(T14497_Q));
KC_DFFRNHQ_X2 T5425 ( .Q(T5425_Q), .D(T11326_Y), .RN(T2063_Y),     .CK(T14497_Q));
KC_DFFRNHQ_X2 T5428 ( .Q(T5428_Q), .D(T11991_Y), .RN(T3221_Y),     .CK(T3209_Y));
KC_DFFRNHQ_X2 T5429 ( .Q(T5429_Q), .D(T2093_Y), .RN(T15008_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T5432 ( .Q(T5432_Q), .D(T2096_Y), .RN(T15008_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T5434 ( .Q(T5434_Q), .D(T15123_Y), .RN(T15008_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T5438 ( .Q(T5438_Q), .D(T2116_Y), .RN(T15011_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T5439 ( .Q(T5439_Q), .D(T12178_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T5441 ( .Q(T5441_Q), .D(T12802_Y), .RN(T15009_Y),     .CK(T14552_Q));
KC_DFFRNHQ_X2 T5442 ( .Q(T5442_Q), .D(T15883_Y), .RN(T15008_Y),     .CK(T14955_Q));
KC_DFFRNHQ_X2 T5449 ( .Q(T5449_Q), .D(T2751_Y), .RN(VDD),     .CK(T2790_Y));
KC_DFFRNHQ_X2 T5451 ( .Q(T5451_Q), .D(T3272_Y), .RN(T15034_Y),     .CK(T3264_Y));
KC_DFFRNHQ_X2 T5452 ( .Q(T5452_Q), .D(T5872_Y), .RN(T15015_Y),     .CK(T14565_Q));
KC_DFFRNHQ_X2 T5455 ( .Q(T5455_Q), .D(T11438_Y), .RN(T15011_Y),     .CK(T14558_Q));
KC_DFFRNHQ_X2 T5461 ( .Q(T5461_Q), .D(T11528_Y), .RN(T15015_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T5462 ( .Q(T5462_Q), .D(T11526_Y), .RN(T2709_Y),     .CK(T3264_Y));
KC_DFFRNHQ_X2 T5463 ( .Q(T5463_Q), .D(T15958_Y), .RN(T15015_Y),     .CK(T14538_Q));
KC_DFFRNHQ_X2 T5465 ( .Q(T5465_Q), .D(T12812_Y), .RN(T15015_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T5473 ( .Q(T5473_Q), .D(T15972_Y), .RN(T2169_Y),     .CK(T14538_Q));
KC_DFFRNHQ_X2 T5474 ( .Q(T5474_Q), .D(T12828_Y), .RN(T2169_Y),     .CK(T14538_Q));
KC_DFFRNHQ_X2 T5479 ( .Q(T5479_Q), .D(T3952_Y), .RN(T15035_Y),     .CK(T3993_Y));
KC_DFFRNHQ_X2 T5481 ( .Q(T5481_Q), .D(T11621_Y), .RN(T4047_Y),     .CK(T14573_Q));
KC_DFFRNHQ_X2 T5486 ( .Q(T5486_Q), .D(T11602_Y), .RN(T15018_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T5488 ( .Q(T5488_Q), .D(T8305_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T16049 ( .Q(T16049_Q), .D(T4683_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T5494 ( .Q(T5494_Q), .D(T11668_Y), .RN(T15021_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T5495 ( .Q(T5495_Q), .D(T8504_Y), .RN(T15035_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T5496 ( .Q(T5496_Q), .D(T12837_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T5497 ( .Q(T5497_Q), .D(T11667_Y), .RN(T15021_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T5498 ( .Q(T5498_Q), .D(T11670_Y), .RN(T5023_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T5499 ( .Q(T5499_Q), .D(T11655_Y), .RN(T5023_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T5501 ( .Q(T5501_Q), .D(T4673_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T5502 ( .Q(T5502_Q), .D(T12836_Y), .RN(T15017_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T5511 ( .Q(T5511_Q), .D(T13171_Y), .RN(T4047_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T5512 ( .Q(T5512_Q), .D(T16127_Y), .RN(T4047_Y),     .CK(T2736_Y));
KC_DFFRNHQ_X2 T5513 ( .Q(T5513_Q), .D(T4727_Y), .RN(T15022_Y),     .CK(T4014_Y));
KC_DFFRNHQ_X2 T5524 ( .Q(T5524_Q), .D(T1828_Y), .RN(T15037_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T5526 ( .Q(T5526_Q), .D(T11755_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T5527 ( .Q(T5527_Q), .D(T13183_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T5528 ( .Q(T5528_Q), .D(T8421_Y), .RN(T4047_Y),     .CK(T3496_Y));
KC_DFFRNHQ_X2 T5529 ( .Q(T5529_Q), .D(T12983_Y), .RN(T2322_Y),     .CK(T14577_Q));
KC_DFFRNHQ_X2 T5530 ( .Q(T5530_Q), .D(T12292_Y), .RN(T4047_Y),     .CK(T14575_Q));
KC_DFFRNHQ_X2 T5532 ( .Q(T5532_Q), .D(T8405_Y), .RN(T4047_Y),     .CK(T3496_Y));
KC_DFFRNHQ_X2 T5536 ( .Q(T5536_Q), .D(T8152_Y), .RN(T15023_Y),     .CK(T14582_Q));
KC_DFFRNHQ_X2 T5538 ( .Q(T5538_Q), .D(T11821_Y), .RN(T2709_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T5541 ( .Q(T5541_Q), .D(T11039_Y), .RN(T15037_Y),     .CK(T14581_Q));
KC_DFFRNHQ_X2 T5543 ( .Q(T5543_Q), .D(T12037_Y), .RN(T4047_Y),     .CK(T3496_Y));
KC_DFFRNHQ_X2 T9353 ( .Q(T9353_Q), .D(T8808_Y), .RN(T15029_Y),     .CK(T178_Y));
KC_DFFRNHQ_X2 T5558 ( .Q(T5558_Q), .D(T1375_Y), .RN(T13053_SN),     .CK(T16078_Y));
KC_DFFRNHQ_X2 T5559 ( .Q(T5559_Q), .D(T11912_Y), .RN(T15029_Y),     .CK(T536_Y));
KC_DFFRNHQ_X2 T5560 ( .Q(T5560_Q), .D(T11865_Y), .RN(T14979_Y),     .CK(T398_Y));
KC_DFFRNHQ_X2 T5561 ( .Q(T5561_Q), .D(T13276_Y), .RN(T7798_Y),     .CK(T14095_Q));
KC_DFFRNHQ_X2 T5562 ( .Q(T5562_Q), .D(T156_Y), .RN(T14975_Y),     .CK(T640_Y));
KC_DFFRNHQ_X2 T5564 ( .Q(T5564_Q), .D(T11853_Y), .RN(T14978_Y),     .CK(T309_Y));
KC_DFFRNHQ_X2 T5565 ( .Q(T5565_Q), .D(T11101_Y), .RN(T14977_Y),     .CK(T855_Y));
KC_DFFRNHQ_X2 T5566 ( .Q(T5566_Q), .D(T11692_Y), .RN(T15037_Y),     .CK(T14576_Q));
KC_DFFRNHQ_X2 T5567 ( .Q(T5567_Q), .D(T15139_Y), .RN(T15021_Y),     .CK(T14557_Q));
KC_DFFRNHQ_X2 T5568 ( .Q(T5568_Q), .D(T8399_Y), .RN(T15035_Y),     .CK(T4045_Y));
KC_DFFRNHQ_X2 T5571 ( .Q(T5571_Q), .D(T12012_Y), .RN(T15018_Y),     .CK(T14574_Q));
KC_DFFRNHQ_X2 T5573 ( .Q(T5573_Q), .D(T4625_Y), .RN(T15017_Y),     .CK(T14962_Q));
KC_DFFRNHQ_X2 T5574 ( .Q(T5574_Q), .D(T10908_Y), .RN(T15008_Y),     .CK(T14553_Q));
KC_DFFRNHQ_X2 T5575 ( .Q(T5575_Q), .D(T10256_Y), .RN(T15009_Y),     .CK(T3209_Y));
KC_DFFRNHQ_X2 T5576 ( .Q(T5576_Q), .D(T12336_Y), .RN(T2063_Y),     .CK(T14497_Q));
KC_DFFRNHQ_X2 T5577 ( .Q(T5577_Q), .D(T2080_Q), .RN(T15806_Q),     .CK(T5725_Y));
KC_NOR2_X1 T21 ( .Y(T21_Y), .A(T22_Y), .B(T15330_Y));
KC_NOR2_X1 T32 ( .Y(T32_Y), .A(T31_Y), .B(T15330_Y));
KC_NOR2_X1 T5582 ( .Y(T5582_Y), .A(T43_Y), .B(T15326_Y));
KC_NOR2_X1 T41 ( .Y(T41_Y), .A(T42_Y), .B(T15326_Y));
KC_NOR2_X1 T66 ( .Y(T66_Y), .A(T67_Y), .B(T13317_Y));
KC_NOR2_X1 T77 ( .Y(T77_Y), .A(T78_Y), .B(T13317_Y));
KC_NOR2_X1 T36 ( .Y(T36_Y), .A(T99_Y), .B(T15322_Y));
KC_NOR2_X1 T96 ( .Y(T96_Y), .A(T91_Y), .B(T15322_Y));
KC_NOR2_X1 T6833 ( .Y(T6833_Y), .A(T200_Y), .B(T6832_Y));
KC_NOR2_X1 T196 ( .Y(T196_Y), .A(GND), .B(T6832_Y));
KC_NOR2_X1 T531 ( .Y(T531_Y), .A(T479_Y), .B(T15370_Y));
KC_NOR2_X1 T464 ( .Y(T464_Y), .A(T467_Y), .B(T15370_Y));
KC_NOR2_X1 T10071 ( .Y(T10071_Y), .A(T533_Y), .B(T15657_Y));
KC_NOR2_X1 T532 ( .Y(T532_Y), .A(T583_Y), .B(T15657_Y));
KC_NOR2_X1 T692 ( .Y(T692_Y), .A(T7685_Y), .B(T7646_Y));
KC_NOR2_X1 T796 ( .Y(T796_Y), .A(T799_Y), .B(T15333_Y));
KC_NOR2_X1 T807 ( .Y(T807_Y), .A(T15720_Y), .B(T15333_Y));
KC_NOR2_X1 T6827 ( .Y(T6827_Y), .A(T892_Y), .B(T15410_Y));
KC_NOR2_X1 T889 ( .Y(T889_Y), .A(T893_Y), .B(T15410_Y));
KC_NOR2_X1 T1029 ( .Y(T1029_Y), .A(T1031_Y), .B(T15672_Y));
KC_NOR2_X1 T1219 ( .Y(T1219_Y), .A(T1241_Y), .B(T15499_Y));
KC_NOR2_X1 T1228 ( .Y(T1228_Y), .A(T1194_Y), .B(T15499_Y));
KC_NOR2_X1 T6435 ( .Y(T6435_Y), .A(T1319_Y), .B(T15345_Y));
KC_NOR2_X1 T6450 ( .Y(T6450_Y), .A(T7351_Y), .B(T9631_Y));
KC_NOR2_X1 T1336 ( .Y(T1336_Y), .A(T7351_Y), .B(T9633_Y));
KC_NOR2_X1 T1343 ( .Y(T1343_Y), .A(T7339_Y), .B(T10424_Y));
KC_NOR2_X1 T1344 ( .Y(T1344_Y), .A(T6748_Y), .B(T10425_Y));
KC_NOR2_X1 T1393 ( .Y(T1393_Y), .A(T1397_Y), .B(T15345_Y));
KC_NOR2_X1 T10240 ( .Y(T10240_Y), .A(T1466_Y), .B(T15416_Y));
KC_NOR2_X1 T6463 ( .Y(T6463_Y), .A(T1528_Y), .B(T15376_Y));
KC_NOR2_X1 T6449 ( .Y(T6449_Y), .A(T1530_Y), .B(T15376_Y));
KC_NOR2_X1 T1547 ( .Y(T1547_Y), .A(T15392_Y), .B(T9610_Y));
KC_NOR2_X1 T16424 ( .Y(T16424_Y), .A(T1570_Y), .B(T15459_Y));
KC_NOR2_X1 T1584 ( .Y(T1584_Y), .A(T8004_Y), .B(T9920_Y));
KC_NOR2_X1 T1585 ( .Y(T1585_Y), .A(T8004_Y), .B(T10319_Y));
KC_NOR2_X1 T1588 ( .Y(T1588_Y), .A(T1590_Y), .B(T15459_Y));
KC_NOR2_X1 T1617 ( .Y(T1617_Y), .A(T15904_Y), .B(T2240_Y));
KC_NOR2_X1 T6452 ( .Y(T6452_Y), .A(T7334_Y), .B(T9611_Y));
KC_NOR2_X1 T1632 ( .Y(T1632_Y), .A(T7334_Y), .B(T9613_Y));
KC_NOR2_X1 T1742 ( .Y(T1742_Y), .A(T15904_Y), .B(T6565_Y));
KC_NOR2_X1 T6434 ( .Y(T6434_Y), .A(T1867_Y), .B(T15346_Y));
KC_NOR2_X1 T6433 ( .Y(T6433_Y), .A(T1864_Y), .B(T15346_Y));
KC_NOR2_X1 T1961 ( .Y(T1961_Y), .A(T1962_Y), .B(T15426_Y));
KC_NOR2_X1 T1980 ( .Y(T1980_Y), .A(T16240_Y), .B(T15426_Y));
KC_NOR2_X1 T6451 ( .Y(T6451_Y), .A(T2444_Y), .B(T15380_Y));
KC_NOR2_X1 T2437 ( .Y(T2437_Y), .A(T2438_Y), .B(T15380_Y));
KC_NOR2_X1 T2531 ( .Y(T2531_Y), .A(T883_Y), .B(T2504_Y));
KC_NOR2_X1 T2532 ( .Y(T2532_Y), .A(T2861_Y), .B(T2504_Y));
KC_NOR2_X1 T2535 ( .Y(T2535_Y), .A(T2501_Y), .B(T2500_Y));
KC_NOR2_X1 T2630 ( .Y(T2630_Y), .A(T2551_Y), .B(T1987_Y));
KC_NOR2_X1 T2761 ( .Y(T2761_Y), .A(T10949_Y), .B(T15853_Y));
KC_NOR2_X1 T2876 ( .Y(T2876_Y), .A(T2838_Y), .B(T6180_Y));
KC_NOR2_X1 T3024 ( .Y(T3024_Y), .A(T475_Y), .B(T9649_Y));
KC_NOR2_X1 T3027 ( .Y(T3027_Y), .A(T475_Y), .B(T9650_Y));
KC_NOR2_X1 T3117 ( .Y(T3117_Y), .A(T16403_Y), .B(T10506_Y));
KC_NOR2_X1 T16304 ( .Y(T16304_Y), .A(T3154_Y), .B(T15508_Y));
KC_NOR2_X1 T3152 ( .Y(T3152_Y), .A(T3159_Y), .B(T15508_Y));
KC_NOR2_X1 T16166 ( .Y(T16166_Y), .A(T3193_Y), .B(T5737_Y));
KC_NOR2_X1 T10255 ( .Y(T10255_Y), .A(T3192_Y), .B(T5737_Y));
KC_NOR2_X1 T3225 ( .Y(T3225_Y), .A(T16239_Y), .B(T15561_Y));
KC_NOR2_X1 T3233 ( .Y(T3233_Y), .A(T3235_Y), .B(T15561_Y));
KC_NOR2_X1 T3315 ( .Y(T3315_Y), .A(T2777_Y), .B(T15858_Y));
KC_NOR2_X1 T3336 ( .Y(T3336_Y), .A(T2778_Y), .B(T15895_Y));
KC_NOR2_X1 T3367 ( .Y(T3367_Y), .A(T16242_Y), .B(T15599_Y));
KC_NOR2_X1 T3411 ( .Y(T3411_Y), .A(T16039_Y), .B(T15623_Y));
KC_NOR2_X1 T6552 ( .Y(T6552_Y), .A(T3501_Y), .B(T6551_Y));
KC_NOR2_X1 T3533 ( .Y(T3533_Y), .A(T3534_Y), .B(T6551_Y));
KC_NOR2_X1 T3611 ( .Y(T3611_Y), .A(T15402_Y), .B(T10470_Y));
KC_NOR2_X1 T3645 ( .Y(T3645_Y), .A(T3648_Y), .B(T15423_Y));
KC_NOR2_X1 T3954 ( .Y(T3954_Y), .A(T5121_Y), .B(T15707_Y));
KC_NOR2_X1 T4196 ( .Y(T4196_Y), .A(T4184_Y), .B(T15362_Y));
KC_NOR2_X1 T4197 ( .Y(T4197_Y), .A(T4192_Y), .B(T15362_Y));
KC_NOR2_X1 T4226 ( .Y(T4226_Y), .A(T4228_Y), .B(T15678_Y));
KC_NOR2_X1 T4330 ( .Y(T4330_Y), .A(T5913_Y), .B(T15510_Y));
KC_NOR2_X1 T6470 ( .Y(T6470_Y), .A(T4856_Y), .B(T15672_Y));
KC_NOR2_X1 T5022 ( .Y(T5022_Y), .A(T4872_Y), .B(T2633_Y));
KC_NOR2_X1 T16443 ( .Y(T16443_Y), .A(T3069_Y), .B(T9832_Y));
KC_NOR2_X1 T5066 ( .Y(T5066_Y), .A(T3317_Y), .B(T15707_Y));
KC_NOR2_X1 T5071 ( .Y(T5071_Y), .A(T4040_Y), .B(T15599_Y));
KC_NOR2_X1 T5131 ( .Y(T5131_Y), .A(T3639_Y), .B(T15423_Y));
KC_NOR2_X1 T5174 ( .Y(T5174_Y), .A(T5176_Y), .B(T15678_Y));
KC_NOR2_X1 T5290 ( .Y(T5290_Y), .A(T1465_Y), .B(T15416_Y));
KC_NOR2_X1 T5393 ( .Y(T5393_Y), .A(T4333_Y), .B(T15510_Y));
KC_NOR2_X1 T5579 ( .Y(T5579_Y), .A(T16402_Y), .B(T9834_Y));
KC_BUF_X10 T26 ( .Y(T26_Y), .A(T21_Y));
KC_BUF_X10 T39 ( .Y(T39_Y), .A(T5582_Y));
KC_BUF_X10 T65 ( .Y(T65_Y), .A(T66_Y));
KC_BUF_X10 T75 ( .Y(T75_Y), .A(T77_Y));
KC_BUF_X10 T104 ( .Y(T104_Y), .A(T36_Y));
KC_BUF_X10 T188 ( .Y(T188_Y), .A(T196_Y));
KC_BUF_X10 T202 ( .Y(T202_Y), .A(T256_Y));
KC_BUF_X10 T469 ( .Y(T469_Y), .A(T464_Y));
KC_BUF_X10 T481 ( .Y(T481_Y), .A(T531_Y));
KC_BUF_X10 T534 ( .Y(T534_Y), .A(T532_Y));
KC_BUF_X10 T539 ( .Y(T539_Y), .A(T10071_Y));
KC_BUF_X10 T117 ( .Y(T117_Y), .A(T807_Y));
KC_BUF_X10 T898 ( .Y(T898_Y), .A(T6827_Y));
KC_BUF_X10 T901 ( .Y(T901_Y), .A(T889_Y));
KC_BUF_X10 T1182 ( .Y(T1182_Y), .A(T6470_Y));
KC_BUF_X10 T1233 ( .Y(T1233_Y), .A(T1219_Y));
KC_BUF_X10 T1234 ( .Y(T1234_Y), .A(T1228_Y));
KC_BUF_X10 T1322 ( .Y(T1322_Y), .A(T6435_Y));
KC_BUF_X10 T1387 ( .Y(T1387_Y), .A(T1393_Y));
KC_BUF_X10 T1531 ( .Y(T1531_Y), .A(T6449_Y));
KC_BUF_X10 T1573 ( .Y(T1573_Y), .A(T16424_Y));
KC_BUF_X10 T1592 ( .Y(T1592_Y), .A(T1588_Y));
KC_BUF_X10 T1871 ( .Y(T1871_Y), .A(T6434_Y));
KC_BUF_X10 T1865 ( .Y(T1865_Y), .A(T6433_Y));
KC_BUF_X10 T2024 ( .Y(T2024_Y), .A(T1970_Q));
KC_BUF_X10 T3008 ( .Y(T3008_Y), .A(T2437_Y));
KC_BUF_X10 T3195 ( .Y(T3195_Y), .A(T10255_Y));
KC_BUF_X10 T3196 ( .Y(T3196_Y), .A(T16166_Y));
KC_BUF_X10 T3232 ( .Y(T3232_Y), .A(T3225_Y));
KC_BUF_X10 T3240 ( .Y(T3240_Y), .A(T3233_Y));
KC_BUF_X10 T3365 ( .Y(T3365_Y), .A(T3367_Y));
KC_BUF_X10 T3502 ( .Y(T3502_Y), .A(T6552_Y));
KC_BUF_X10 T3535 ( .Y(T3535_Y), .A(T3533_Y));
KC_BUF_X10 T3649 ( .Y(T3649_Y), .A(T3645_Y));
KC_BUF_X10 T3959 ( .Y(T3959_Y), .A(T3954_Y));
KC_BUF_X10 T4173 ( .Y(T4173_Y), .A(T10602_Y));
KC_BUF_X10 T4185 ( .Y(T4185_Y), .A(T4196_Y));
KC_BUF_X10 T4201 ( .Y(T4201_Y), .A(T4197_Y));
KC_BUF_X10 T4209 ( .Y(T4209_Y), .A(T5174_Y));
KC_BUF_X10 T4223 ( .Y(T4223_Y), .A(T4226_Y));
KC_BUF_X10 T4337 ( .Y(T4337_Y), .A(T4330_Y));
KC_BUF_X10 T4621 ( .Y(T4621_Y), .A(T8265_Y));
KC_BUF_X10 T4888 ( .Y(T4888_Y), .A(T10240_Y));
KC_BUF_X10 T4894 ( .Y(T4894_Y), .A(T6463_Y));
KC_BUF_X10 T5073 ( .Y(T5073_Y), .A(T5071_Y));
KC_BUF_X10 T5133 ( .Y(T5133_Y), .A(T5131_Y));
KC_BUF_X10 T5186 ( .Y(T5186_Y), .A(T96_Y));
KC_BUF_X10 T5201 ( .Y(T5201_Y), .A(T796_Y));
KC_BUF_X10 T5584 ( .Y(T5584_Y), .A(T41_Y));
KC_BUF_X10 T5230 ( .Y(T5230_Y), .A(T32_Y));
KC_BUF_X10 T5235 ( .Y(T5235_Y), .A(T1029_Y));
KC_BUF_X10 T5245 ( .Y(T5245_Y), .A(T6451_Y));
KC_BUF_X10 T5285 ( .Y(T5285_Y), .A(T1961_Y));
KC_BUF_X10 T5291 ( .Y(T5291_Y), .A(T5290_Y));
KC_BUF_X10 T5314 ( .Y(T5314_Y), .A(T13013_Q));
KC_BUF_X10 T1497 ( .Y(T1497_Y), .A(T5393_Y));
KC_BUF_X10 T5392 ( .Y(T5392_Y), .A(T16304_Y));
KC_BUF_X10 T5398 ( .Y(T5398_Y), .A(T3152_Y));
KC_BUF_X10 T5475 ( .Y(T5475_Y), .A(T5066_Y));
KC_BUF_X10 T5580 ( .Y(T5580_Y), .A(T1980_Y));
KC_BUF_X2 T152 ( .Y(T152_Y), .A(T5349_Y));
KC_BUF_X2 T156 ( .Y(T156_Y), .A(T15786_Y));
KC_BUF_X2 T176 ( .Y(T176_Y), .A(T11205_Y));
KC_BUF_X2 T186 ( .Y(T186_Y), .A(T11234_Y));
KC_BUF_X2 T205 ( .Y(T205_Y), .A(T9394_Y));
KC_BUF_X2 T206 ( .Y(T206_Y), .A(T220_Y));
KC_BUF_X2 T214 ( .Y(T214_Y), .A(T11235_Y));
KC_BUF_X2 T221 ( .Y(T221_Y), .A(T8706_Y));
KC_BUF_X2 T222 ( .Y(T222_Y), .A(T221_Y));
KC_BUF_X2 T254 ( .Y(T254_Y), .A(T1430_Y));
KC_BUF_X2 T271 ( .Y(T271_Y), .A(T15718_Y));
KC_BUF_X2 T295 ( .Y(T295_Y), .A(T6961_Y));
KC_BUF_X2 T305 ( .Y(T305_Y), .A(T8722_Y));
KC_BUF_X2 T325 ( .Y(T325_Y), .A(T7290_Y));
KC_BUF_X2 T328 ( .Y(T328_Y), .A(T7288_Y));
KC_BUF_X2 T336 ( .Y(T336_Y), .A(T7431_Y));
KC_BUF_X2 T346 ( .Y(T346_Y), .A(T7424_Y));
KC_BUF_X2 T357 ( .Y(T357_Y), .A(T11198_Y));
KC_BUF_X2 T371 ( .Y(T371_Y), .A(T350_Y));
KC_BUF_X2 T382 ( .Y(T382_Y), .A(T350_Y));
KC_BUF_X2 T390 ( .Y(T390_Y), .A(T841_Y));
KC_BUF_X2 T393 ( .Y(T393_Y), .A(T15109_Y));
KC_BUF_X2 T395 ( .Y(T395_Y), .A(T11308_Y));
KC_BUF_X2 T427 ( .Y(T427_Y), .A(T2392_Y));
KC_BUF_X2 T430 ( .Y(T430_Y), .A(T15905_Y));
KC_BUF_X2 T447 ( .Y(T447_Y), .A(T11060_Y));
KC_BUF_X2 T454 ( .Y(T454_Y), .A(T6904_Y));
KC_BUF_X2 T455 ( .Y(T455_Y), .A(T11068_Y));
KC_BUF_X2 T472 ( .Y(T472_Y), .A(T8813_Y));
KC_BUF_X2 T492 ( .Y(T492_Y), .A(T7245_Y));
KC_BUF_X2 T565 ( .Y(T565_Y), .A(T8984_Y));
KC_BUF_X2 T586 ( .Y(T586_Y), .A(T604_Q));
KC_BUF_X2 T593 ( .Y(T593_Y), .A(T5406_Q));
KC_BUF_X2 T615 ( .Y(T615_Y), .A(T15914_Y));
KC_BUF_X2 T616 ( .Y(T616_Y), .A(T13088_Y));
KC_BUF_X2 T617 ( .Y(T617_Y), .A(T16150_Y));
KC_BUF_X2 T618 ( .Y(T618_Y), .A(T15922_Y));
KC_BUF_X2 T619 ( .Y(T619_Y), .A(T1752_Y));
KC_BUF_X2 T675 ( .Y(T675_Y), .A(T7370_Y));
KC_BUF_X2 T746 ( .Y(T746_Y), .A(T9008_Y));
KC_BUF_X2 T748 ( .Y(T748_Y), .A(T749_Y));
KC_BUF_X2 T749 ( .Y(T749_Y), .A(T8115_Y));
KC_BUF_X2 T753 ( .Y(T753_Y), .A(T8094_Y));
KC_BUF_X2 T757 ( .Y(T757_Y), .A(T754_Q));
KC_BUF_X2 T758 ( .Y(T758_Y), .A(T977_Q));
KC_BUF_X2 T759 ( .Y(T759_Y), .A(T5384_Q));
KC_BUF_X2 T766 ( .Y(T766_Y), .A(T1157_Q));
KC_BUF_X2 T773 ( .Y(T773_Y), .A(T1154_Q));
KC_BUF_X2 T808 ( .Y(T808_Y), .A(T11064_Y));
KC_BUF_X2 T819 ( .Y(T819_Y), .A(T6948_Y));
KC_BUF_X2 T839 ( .Y(T839_Y), .A(T7078_Y));
KC_BUF_X2 T842 ( .Y(T842_Y), .A(T7075_Y));
KC_BUF_X2 T867 ( .Y(T867_Y), .A(T7298_Y));
KC_BUF_X2 T962 ( .Y(T962_Y), .A(T8095_Y));
KC_BUF_X2 T972 ( .Y(T972_Y), .A(T15485_Y));
KC_BUF_X2 T973 ( .Y(T973_Y), .A(T9038_Y));
KC_BUF_X2 T985 ( .Y(T985_Y), .A(T4862_Q));
KC_BUF_X2 T10534 ( .Y(T10534_Y), .A(T760_Q));
KC_BUF_X2 T993 ( .Y(T993_Y), .A(T1244_Y));
KC_BUF_X2 T994 ( .Y(T994_Y), .A(T995_Q));
KC_BUF_X2 T1014 ( .Y(T1014_Y), .A(T978_Q));
KC_BUF_X2 T1015 ( .Y(T1015_Y), .A(T10259_Y));
KC_BUF_X2 T1017 ( .Y(T1017_Y), .A(T1000_Q));
KC_BUF_X2 T1018 ( .Y(T1018_Y), .A(T983_Q));
KC_BUF_X2 T1019 ( .Y(T1019_Y), .A(T761_Q));
KC_BUF_X2 T1020 ( .Y(T1020_Y), .A(T997_Q));
KC_BUF_X2 T1021 ( .Y(T1021_Y), .A(T765_Q));
KC_BUF_X2 T1025 ( .Y(T1025_Y), .A(T9457_Q));
KC_BUF_X2 T1036 ( .Y(T1036_Y), .A(T11104_Y));
KC_BUF_X2 T1093 ( .Y(T1093_Y), .A(T8789_Y));
KC_BUF_X2 T1146 ( .Y(T1146_Y), .A(T996_Q));
KC_BUF_X2 T1155 ( .Y(T1155_Y), .A(T1152_Q));
KC_BUF_X2 T1161 ( .Y(T1161_Y), .A(T767_Q));
KC_BUF_X2 T1171 ( .Y(T1171_Y), .A(T9459_Q));
KC_BUF_X2 T1172 ( .Y(T1172_Y), .A(T9458_Q));
KC_BUF_X2 T1173 ( .Y(T1173_Y), .A(T5385_Q));
KC_BUF_X2 T1174 ( .Y(T1174_Y), .A(T999_Q));
KC_BUF_X2 T1175 ( .Y(T1175_Y), .A(T1159_Q));
KC_BUF_X2 T1176 ( .Y(T1176_Y), .A(T1160_Q));
KC_BUF_X2 T1177 ( .Y(T1177_Y), .A(T1158_Q));
KC_BUF_X2 T1178 ( .Y(T1178_Y), .A(T963_Q));
KC_BUF_X2 T1251 ( .Y(T1251_Y), .A(T1156_Q));
KC_BUF_X2 T1253 ( .Y(T1253_Y), .A(T1254_Y));
KC_BUF_X2 T1254 ( .Y(T1254_Y), .A(T1309_Y));
KC_BUF_X2 T1267 ( .Y(T1267_Y), .A(T1151_Q));
KC_BUF_X2 T1268 ( .Y(T1268_Y), .A(T16232_Q));
KC_BUF_X2 T1269 ( .Y(T1269_Y), .A(T1153_Q));
KC_BUF_X2 T1280 ( .Y(T1280_Y), .A(T1300_Y));
KC_BUF_X2 T1281 ( .Y(T1281_Y), .A(T15920_Y));
KC_BUF_X2 T1282 ( .Y(T1282_Y), .A(T1292_Y));
KC_BUF_X2 T1291 ( .Y(T1291_Y), .A(T1315_Y));
KC_BUF_X2 T1292 ( .Y(T1292_Y), .A(T1280_Y));
KC_BUF_X2 T1293 ( .Y(T1293_Y), .A(T1301_Y));
KC_BUF_X2 T1294 ( .Y(T1294_Y), .A(T1312_Y));
KC_BUF_X2 T1295 ( .Y(T1295_Y), .A(T1294_Y));
KC_BUF_X2 T1296 ( .Y(T1296_Y), .A(T1307_Y));
KC_BUF_X2 T1297 ( .Y(T1297_Y), .A(T1314_Y));
KC_BUF_X2 T1298 ( .Y(T1298_Y), .A(T1299_Y));
KC_BUF_X2 T1299 ( .Y(T1299_Y), .A(T1282_Y));
KC_BUF_X2 T1300 ( .Y(T1300_Y), .A(T1293_Y));
KC_BUF_X2 T1301 ( .Y(T1301_Y), .A(T1274_Y));
KC_BUF_X2 T1302 ( .Y(T1302_Y), .A(T4875_Y));
KC_BUF_X2 T1303 ( .Y(T1303_Y), .A(T1253_Y));
KC_BUF_X2 T1304 ( .Y(T1304_Y), .A(T4877_Y));
KC_BUF_X2 T1305 ( .Y(T1305_Y), .A(T1311_Y));
KC_BUF_X2 T1306 ( .Y(T1306_Y), .A(T1296_Y));
KC_BUF_X2 T1307 ( .Y(T1307_Y), .A(T1313_Y));
KC_BUF_X2 T1308 ( .Y(T1308_Y), .A(T1303_Y));
KC_BUF_X2 T1309 ( .Y(T1309_Y), .A(T4874_Y));
KC_BUF_X2 T1310 ( .Y(T1310_Y), .A(T1305_Y));
KC_BUF_X2 T1311 ( .Y(T1311_Y), .A(T1295_Y));
KC_BUF_X2 T1312 ( .Y(T1312_Y), .A(T1306_Y));
KC_BUF_X2 T1313 ( .Y(T1313_Y), .A(T1297_Y));
KC_BUF_X2 T1314 ( .Y(T1314_Y), .A(T1316_Y));
KC_BUF_X2 T1315 ( .Y(T1315_Y), .A(T1310_Y));
KC_BUF_X2 T1316 ( .Y(T1316_Y), .A(T1317_Y));
KC_BUF_X2 T1317 ( .Y(T1317_Y), .A(T10218_Y));
KC_BUF_X2 T1337 ( .Y(T1337_Y), .A(T7338_Y));
KC_BUF_X2 T1338 ( .Y(T1338_Y), .A(T2027_Y));
KC_BUF_X2 T1377 ( .Y(T1377_Y), .A(T5414_Y));
KC_BUF_X2 T1418 ( .Y(T1418_Y), .A(T9059_Y));
KC_BUF_X2 T1419 ( .Y(T1419_Y), .A(T9059_Y));
KC_BUF_X2 T1431 ( .Y(T1431_Y), .A(T9059_Y));
KC_BUF_X2 T1453 ( .Y(T1453_Y), .A(T4885_Y));
KC_BUF_X2 T1476 ( .Y(T1476_Y), .A(T16449_Y));
KC_BUF_X2 T1483 ( .Y(T1483_Y), .A(T16245_Y));
KC_BUF_X2 T1484 ( .Y(T1484_Y), .A(T9957_Y));
KC_BUF_X2 T1491 ( .Y(T1491_Y), .A(T9059_Y));
KC_BUF_X2 T1492 ( .Y(T1492_Y), .A(T9059_Y));
KC_BUF_X2 T1493 ( .Y(T1493_Y), .A(T9059_Y));
KC_BUF_X2 T1535 ( .Y(T1535_Y), .A(T7017_Y));
KC_BUF_X2 T1545 ( .Y(T1545_Y), .A(T2027_Y));
KC_BUF_X2 T1571 ( .Y(T1571_Y), .A(T10195_Y));
KC_BUF_X2 T1586 ( .Y(T1586_Y), .A(T16164_Y));
KC_BUF_X2 T1654 ( .Y(T1654_Y), .A(T1656_Y));
KC_BUF_X2 T1655 ( .Y(T1655_Y), .A(T1672_Y));
KC_BUF_X2 T1656 ( .Y(T1656_Y), .A(T1669_Y));
KC_BUF_X2 T1657 ( .Y(T1657_Y), .A(T1655_Y));
KC_BUF_X2 T1658 ( .Y(T1658_Y), .A(T1657_Y));
KC_BUF_X2 T1659 ( .Y(T1659_Y), .A(T844_Y));
KC_BUF_X2 T1663 ( .Y(T1663_Y), .A(T1673_Y));
KC_BUF_X2 T1664 ( .Y(T1664_Y), .A(T4918_Y));
KC_BUF_X2 T1667 ( .Y(T1667_Y), .A(T844_Y));
KC_BUF_X2 T1668 ( .Y(T1668_Y), .A(T844_Y));
KC_BUF_X2 T1669 ( .Y(T1669_Y), .A(T1670_Y));
KC_BUF_X2 T1670 ( .Y(T1670_Y), .A(T1674_Y));
KC_BUF_X2 T1671 ( .Y(T1671_Y), .A(T1654_Y));
KC_BUF_X2 T1672 ( .Y(T1672_Y), .A(T1677_Y));
KC_BUF_X2 T1673 ( .Y(T1673_Y), .A(T1667_Y));
KC_BUF_X2 T1674 ( .Y(T1674_Y), .A(T844_Y));
KC_BUF_X2 T1677 ( .Y(T1677_Y), .A(T1659_Y));
KC_BUF_X2 T1679 ( .Y(T1679_Y), .A(T1684_Y));
KC_BUF_X2 T1680 ( .Y(T1680_Y), .A(T5366_Q));
KC_BUF_X2 T1683 ( .Y(T1683_Y), .A(T1685_Y));
KC_BUF_X2 T1684 ( .Y(T1684_Y), .A(T1683_Y));
KC_BUF_X2 T1685 ( .Y(T1685_Y), .A(T1668_Y));
KC_BUF_X2 T1688 ( .Y(T1688_Y), .A(T1700_Y));
KC_BUF_X2 T1689 ( .Y(T1689_Y), .A(T1712_Y));
KC_BUF_X2 T1692 ( .Y(T1692_Y), .A(T1715_Y));
KC_BUF_X2 T1693 ( .Y(T1693_Y), .A(T1699_Y));
KC_BUF_X2 T1698 ( .Y(T1698_Y), .A(T1704_Y));
KC_BUF_X2 T1699 ( .Y(T1699_Y), .A(T1688_Y));
KC_BUF_X2 T1700 ( .Y(T1700_Y), .A(T1701_Y));
KC_BUF_X2 T1701 ( .Y(T1701_Y), .A(T16192_Y));
KC_BUF_X2 T1702 ( .Y(T1702_Y), .A(T16192_Y));
KC_BUF_X2 T1703 ( .Y(T1703_Y), .A(T1698_Y));
KC_BUF_X2 T1704 ( .Y(T1704_Y), .A(T1705_Y));
KC_BUF_X2 T1705 ( .Y(T1705_Y), .A(T1706_Y));
KC_BUF_X2 T1706 ( .Y(T1706_Y), .A(T1702_Y));
KC_BUF_X2 T1710 ( .Y(T1710_Y), .A(T1689_Y));
KC_BUF_X2 T1711 ( .Y(T1711_Y), .A(T1716_Y));
KC_BUF_X2 T1712 ( .Y(T1712_Y), .A(T16435_Q));
KC_BUF_X2 T1713 ( .Y(T1713_Y), .A(T1718_Y));
KC_BUF_X2 T1715 ( .Y(T1715_Y), .A(T1693_Y));
KC_BUF_X2 T1716 ( .Y(T1716_Y), .A(T1710_Y));
KC_BUF_X2 T1718 ( .Y(T1718_Y), .A(T16470_Q));
KC_BUF_X2 T1733 ( .Y(T1733_Y), .A(T2021_Y));
KC_BUF_X2 T1737 ( .Y(T1737_Y), .A(T1723_Q));
KC_BUF_X2 T1827 ( .Y(T1827_Y), .A(T2351_Y));
KC_BUF_X2 T1828 ( .Y(T1828_Y), .A(T1827_Y));
KC_BUF_X2 T1831 ( .Y(T1831_Y), .A(T6216_Y));
KC_BUF_X2 T1845 ( .Y(T1845_Y), .A(T1845_A));
KC_BUF_X2 T1846 ( .Y(T1846_Y), .A(T1845_Y));
KC_BUF_X2 T1847 ( .Y(T1847_Y), .A(T11838_Y));
KC_BUF_X2 T1930 ( .Y(T1930_Y), .A(T9059_Y));
KC_BUF_X2 T1972 ( .Y(T1972_Y), .A(T1675_Q));
KC_BUF_X2 T1973 ( .Y(T1973_Y), .A(T1972_Y));
KC_BUF_X2 T1974 ( .Y(T1974_Y), .A(T1975_Y));
KC_BUF_X2 T1975 ( .Y(T1975_Y), .A(T1675_Q));
KC_BUF_X2 T1976 ( .Y(T1976_Y), .A(T1979_Y));
KC_BUF_X2 T1977 ( .Y(T1977_Y), .A(T4976_Y));
KC_BUF_X2 T1979 ( .Y(T1979_Y), .A(T1973_Y));
KC_BUF_X2 T2004 ( .Y(T2004_Y), .A(T2022_Y));
KC_BUF_X2 T2011 ( .Y(T2011_Y), .A(T5549_Y));
KC_BUF_X2 T2019 ( .Y(T2019_Y), .A(T2582_Y));
KC_BUF_X2 T2022 ( .Y(T2022_Y), .A(T4975_Y));
KC_BUF_X2 T2044 ( .Y(T2044_Y), .A(T1734_Q));
KC_BUF_X2 T2045 ( .Y(T2045_Y), .A(T2046_Y));
KC_BUF_X2 T2046 ( .Y(T2046_Y), .A(T2044_Y));
KC_BUF_X2 T2052 ( .Y(T2052_Y), .A(T1737_Y));
KC_BUF_X2 T2076 ( .Y(T2076_Y), .A(T2113_Q));
KC_BUF_X2 T2077 ( .Y(T2077_Y), .A(T13060_Y));
KC_BUF_X2 T2079 ( .Y(T2079_Y), .A(T14966_Y));
KC_BUF_X2 T2111 ( .Y(T2111_Y), .A(T15990_Q));
KC_BUF_X2 T2117 ( .Y(T2117_Y), .A(T5987_Q));
KC_BUF_X2 T2177 ( .Y(T2177_Y), .A(T2178_Y));
KC_BUF_X2 T2178 ( .Y(T2178_Y), .A(T16007_Q));
KC_BUF_X2 T2179 ( .Y(T2179_Y), .A(T16018_Q));
KC_BUF_X2 T2180 ( .Y(T2180_Y), .A(T2179_Y));
KC_BUF_X2 T2184 ( .Y(T2184_Y), .A(T2761_Y));
KC_BUF_X2 T2187 ( .Y(T2187_Y), .A(T4966_Y));
KC_BUF_X2 T2213 ( .Y(T2213_Y), .A(T5480_Q));
KC_BUF_X2 T2214 ( .Y(T2214_Y), .A(T2809_Q));
KC_BUF_X2 T2351 ( .Y(T2351_Y), .A(T4927_Y));
KC_BUF_X2 T2358 ( .Y(T2358_Y), .A(T11042_Y));
KC_BUF_X2 T2365 ( .Y(T2365_Y), .A(T16151_Y));
KC_BUF_X2 T2400 ( .Y(T2400_Y), .A(T2362_Y));
KC_BUF_X2 T2449 ( .Y(T2449_Y), .A(T10239_Y));
KC_BUF_X2 T2450 ( .Y(T2450_Y), .A(T10195_Y));
KC_BUF_X2 T2452 ( .Y(T2452_Y), .A(T9059_Y));
KC_BUF_X2 T2491 ( .Y(T2491_Y), .A(T10195_Y));
KC_BUF_X2 T2494 ( .Y(T2494_Y), .A(T4252_Y));
KC_BUF_X2 T2524 ( .Y(T2524_Y), .A(T8453_Y));
KC_BUF_X2 T2527 ( .Y(T2527_Y), .A(T2524_Y));
KC_BUF_X2 T2528 ( .Y(T2528_Y), .A(T8453_Y));
KC_BUF_X2 T2542 ( .Y(T2542_Y), .A(T2528_Y));
KC_BUF_X2 T2543 ( .Y(T2543_Y), .A(T16169_Y));
KC_BUF_X2 T2544 ( .Y(T2544_Y), .A(T12670_Y));
KC_BUF_X2 T2578 ( .Y(T2578_Y), .A(T2581_Y));
KC_BUF_X2 T2579 ( .Y(T2579_Y), .A(T1103_Y));
KC_BUF_X2 T2580 ( .Y(T2580_Y), .A(T2579_Y));
KC_BUF_X2 T2581 ( .Y(T2581_Y), .A(T2580_Y));
KC_BUF_X2 T2582 ( .Y(T2582_Y), .A(T2578_Y));
KC_BUF_X2 T2590 ( .Y(T2590_Y), .A(T10195_Y));
KC_BUF_X2 T2651 ( .Y(T2651_Y), .A(T9059_Y));
KC_BUF_X2 T2688 ( .Y(T2688_Y), .A(T2709_Y));
KC_BUF_X2 T2762 ( .Y(T2762_Y), .A(T11546_Y));
KC_BUF_X2 T2840 ( .Y(T2840_Y), .A(T2825_Y));
KC_BUF_X2 T2845 ( .Y(T2845_Y), .A(T16052_Y));
KC_BUF_X2 T2951 ( .Y(T2951_Y), .A(T2912_Y));
KC_BUF_X2 T2956 ( .Y(T2956_Y), .A(T4142_Y));
KC_BUF_X2 T3025 ( .Y(T3025_Y), .A(T9059_Y));
KC_BUF_X2 T3080 ( .Y(T3080_Y), .A(T3781_Y));
KC_BUF_X2 T3081 ( .Y(T3081_Y), .A(T3780_Y));
KC_BUF_X2 T3210 ( .Y(T3210_Y), .A(T11986_Y));
KC_BUF_X2 T3221 ( .Y(T3221_Y), .A(T2709_Y));
KC_BUF_X2 T3255 ( .Y(T3255_Y), .A(T10637_Y));
KC_BUF_X2 T3265 ( .Y(T3265_Y), .A(T5874_Y));
KC_BUF_X2 T3266 ( .Y(T3266_Y), .A(T3268_Y));
KC_BUF_X2 T3269 ( .Y(T3269_Y), .A(T2747_Y));
KC_BUF_X2 T3280 ( .Y(T3280_Y), .A(T3248_Y));
KC_BUF_X2 T3283 ( .Y(T3283_Y), .A(T11456_Y));
KC_BUF_X2 T3303 ( .Y(T3303_Y), .A(T10639_Y));
KC_BUF_X2 T3308 ( .Y(T3308_Y), .A(T9227_Y));
KC_BUF_X2 T3585 ( .Y(T3585_Y), .A(T9059_Y));
KC_BUF_X2 T3640 ( .Y(T3640_Y), .A(T2027_Y));
KC_BUF_X2 T3676 ( .Y(T3676_Y), .A(T3775_Y));
KC_BUF_X2 T3677 ( .Y(T3677_Y), .A(T3774_Y));
KC_BUF_X2 T3678 ( .Y(T3678_Y), .A(T9059_Y));
KC_BUF_X2 T3679 ( .Y(T3679_Y), .A(T16449_Y));
KC_BUF_X2 T3682 ( .Y(T3682_Y), .A(T9059_Y));
KC_BUF_X2 T3684 ( .Y(T3684_Y), .A(T2027_Y));
KC_BUF_X2 T3719 ( .Y(T3719_Y), .A(T16063_Y));
KC_BUF_X2 T3735 ( .Y(T3735_Y), .A(T9059_Y));
KC_BUF_X2 T3973 ( .Y(T3973_Y), .A(T3301_Y));
KC_BUF_X2 T3984 ( .Y(T3984_Y), .A(T15892_Y));
KC_BUF_X2 T3996 ( .Y(T3996_Y), .A(T11429_Y));
KC_BUF_X2 T4008 ( .Y(T4008_Y), .A(T3373_Y));
KC_BUF_X2 T4097 ( .Y(T4097_Y), .A(T4715_Y));
KC_BUF_X2 T4283 ( .Y(T4283_Y), .A(T9059_Y));
KC_BUF_X2 T4426 ( .Y(T4426_Y), .A(T5148_Y));
KC_BUF_X2 T4462 ( .Y(T4462_Y), .A(T11370_Y));
KC_BUF_X2 T4505 ( .Y(T4505_Y), .A(T11455_Y));
KC_BUF_X2 T4571 ( .Y(T4571_Y), .A(T11558_Y));
KC_BUF_X2 T4611 ( .Y(T4611_Y), .A(T3969_Y));
KC_BUF_X2 T4612 ( .Y(T4612_Y), .A(T6326_Y));
KC_BUF_X2 T4613 ( .Y(T4613_Y), .A(T4598_Y));
KC_BUF_X2 T4624 ( .Y(T4624_Y), .A(T5160_Y));
KC_BUF_X2 T4625 ( .Y(T4625_Y), .A(T4624_Y));
KC_BUF_X2 T4745 ( .Y(T4745_Y), .A(T4718_Q));
KC_BUF_X2 T15425 ( .Y(T15425_Y), .A(T11238_Y));
KC_BUF_X2 T15732 ( .Y(T15732_Y), .A(T7668_Y));
KC_BUF_X2 T4842 ( .Y(T4842_Y), .A(T15795_Q));
KC_BUF_X2 T4844 ( .Y(T4844_Y), .A(T1005_Q));
KC_BUF_X2 T15327 ( .Y(T15327_Y), .A(T5387_Q));
KC_BUF_X2 T10262 ( .Y(T10262_Y), .A(T762_Q));
KC_BUF_X2 T10260 ( .Y(T10260_Y), .A(T768_Q));
KC_BUF_X2 T10259 ( .Y(T10259_Y), .A(T9005_Y));
KC_BUF_X2 T4853 ( .Y(T4853_Y), .A(T6245_Y));
KC_BUF_X2 T4873 ( .Y(T4873_Y), .A(T4951_Y));
KC_BUF_X2 T4874 ( .Y(T4874_Y), .A(T4876_Y));
KC_BUF_X2 T4875 ( .Y(T4875_Y), .A(T1308_Y));
KC_BUF_X2 T4876 ( .Y(T4876_Y), .A(T1304_Y));
KC_BUF_X2 T4877 ( .Y(T4877_Y), .A(T4878_Y));
KC_BUF_X2 T4878 ( .Y(T4878_Y), .A(T4873_Y));
KC_BUF_X2 T4884 ( .Y(T4884_Y), .A(T16449_Y));
KC_BUF_X2 T4885 ( .Y(T4885_Y), .A(T9059_Y));
KC_BUF_X2 T4889 ( .Y(T4889_Y), .A(T16063_Y));
KC_BUF_X2 T4918 ( .Y(T4918_Y), .A(T1663_Y));
KC_BUF_X2 T4923 ( .Y(T4923_Y), .A(T1703_Y));
KC_BUF_X2 T4927 ( .Y(T4927_Y), .A(T8350_Y));
KC_BUF_X2 T4965 ( .Y(T4965_Y), .A(T11728_Y));
KC_BUF_X2 T4966 ( .Y(T4966_Y), .A(T16010_Q));
KC_BUF_X2 T4975 ( .Y(T4975_Y), .A(T5578_Y));
KC_BUF_X2 T4976 ( .Y(T4976_Y), .A(T1974_Y));
KC_BUF_X2 T5028 ( .Y(T5028_Y), .A(T10239_Y));
KC_BUF_X2 T5068 ( .Y(T5068_Y), .A(T11578_Y));
KC_BUF_X2 T5134 ( .Y(T5134_Y), .A(T16063_Y));
KC_BUF_X2 T5154 ( .Y(T5154_Y), .A(T15981_Y));
KC_BUF_X2 T5160 ( .Y(T5160_Y), .A(T5161_Y));
KC_BUF_X2 T5161 ( .Y(T5161_Y), .A(T8465_Y));
KC_BUF_X2 T5169 ( .Y(T5169_Y), .A(T5168_Y));
KC_BUF_X2 T5173 ( .Y(T5173_Y), .A(T13873_Q));
KC_BUF_X2 T5318 ( .Y(T5318_Y), .A(T809_Y));
KC_BUF_X2 T5394 ( .Y(T5394_Y), .A(T2052_Y));
KC_BUF_X2 T5418 ( .Y(T5418_Y), .A(T15921_Y));
KC_BUF_X2 T5578 ( .Y(T5578_Y), .A(T13008_Q));
KC_BUF_X2 T1 ( .Y(T1_Y), .A(T11567_Y));

endmodule
